//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 0 1 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n829, new_n830, new_n831, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT86), .Z(new_n203));
  XNOR2_X1  g002(.A(G141gat), .B(G148gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n204), .A2(KEYINPUT2), .ZN(new_n205));
  XNOR2_X1  g004(.A(G155gat), .B(G162gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n204), .A2(KEYINPUT80), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n204), .A2(KEYINPUT80), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(new_n206), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT81), .B(G155gat), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n212), .B1(new_n213), .B2(G162gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n208), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G211gat), .B(G218gat), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT22), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT75), .B(G211gat), .ZN(new_n220));
  INV_X1    g019(.A(G218gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT76), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n222), .B(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT77), .ZN(new_n225));
  XNOR2_X1  g024(.A(G197gat), .B(G204gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n225), .B1(new_n224), .B2(new_n226), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n218), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n224), .A2(new_n226), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT77), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n232), .A2(new_n217), .A3(new_n227), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT29), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n230), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  XOR2_X1   g034(.A(KEYINPUT83), .B(KEYINPUT3), .Z(new_n236));
  AOI21_X1  g035(.A(new_n216), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n230), .A2(new_n233), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n216), .A2(new_n236), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(new_n234), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n203), .B1(new_n237), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n235), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n215), .B(KEYINPUT82), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n202), .B1(new_n238), .B2(new_n240), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n242), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT87), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G22gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n250), .A2(new_n251), .ZN(new_n255));
  XNOR2_X1  g054(.A(G78gat), .B(G106gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(KEYINPUT31), .ZN(new_n257));
  INV_X1    g056(.A(G50gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n254), .B1(new_n255), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT87), .B1(new_n242), .B2(new_n249), .ZN(new_n261));
  INV_X1    g060(.A(new_n259), .ZN(new_n262));
  NOR3_X1   g061(.A1(new_n261), .A2(G22gat), .A3(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n253), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n255), .A2(new_n254), .A3(new_n259), .ZN(new_n265));
  OAI21_X1  g064(.A(G22gat), .B1(new_n261), .B2(new_n262), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(new_n252), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G15gat), .B(G43gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(G71gat), .B(G99gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT25), .ZN(new_n273));
  XOR2_X1   g072(.A(KEYINPUT67), .B(G190gat), .Z(new_n274));
  INV_X1    g073(.A(G183gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n279));
  AND2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n273), .B1(new_n276), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G169gat), .ZN(new_n282));
  INV_X1    g081(.A(G176gat), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT66), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT23), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n282), .A2(new_n283), .ZN(new_n287));
  NOR2_X1   g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288));
  NOR3_X1   g087(.A1(new_n288), .A2(KEYINPUT66), .A3(KEYINPUT23), .ZN(new_n289));
  NOR3_X1   g088(.A1(new_n286), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  AND2_X1   g089(.A1(new_n281), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(G190gat), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n277), .B1(new_n275), .B2(new_n292), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n279), .A2(KEYINPUT65), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT65), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT25), .B1(new_n290), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(KEYINPUT68), .B1(new_n291), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n297), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT68), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n281), .A2(new_n290), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT27), .B(G183gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n274), .A2(new_n303), .ZN(new_n304));
  AOI22_X1  g103(.A1(new_n304), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT26), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n287), .B1(new_n306), .B2(new_n288), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n307), .B1(new_n306), .B2(new_n288), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n305), .B(new_n308), .C1(KEYINPUT28), .C2(new_n304), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n298), .A2(new_n302), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G113gat), .ZN(new_n311));
  INV_X1    g110(.A(G120gat), .ZN(new_n312));
  AOI21_X1  g111(.A(KEYINPUT1), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n313), .B1(new_n311), .B2(new_n312), .ZN(new_n314));
  XNOR2_X1  g113(.A(KEYINPUT69), .B(G134gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n315), .A2(KEYINPUT70), .A3(G127gat), .ZN(new_n316));
  INV_X1    g115(.A(G127gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G134gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT70), .B1(new_n315), .B2(G127gat), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n314), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  XOR2_X1   g120(.A(G127gat), .B(G134gat), .Z(new_n322));
  OR2_X1    g121(.A1(new_n314), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT71), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT71), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n321), .A2(new_n326), .A3(new_n323), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n310), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT72), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n310), .A2(new_n328), .A3(KEYINPUT72), .ZN(new_n332));
  OR2_X1    g131(.A1(new_n310), .A2(new_n328), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G227gat), .A2(G233gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n335), .B(KEYINPUT64), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT33), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n272), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT73), .B1(new_n337), .B2(KEYINPUT32), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT73), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT32), .ZN(new_n342));
  AOI211_X1 g141(.A(new_n341), .B(new_n342), .C1(new_n334), .C2(new_n336), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n339), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n337), .B(KEYINPUT32), .C1(new_n338), .C2(new_n272), .ZN(new_n345));
  INV_X1    g144(.A(new_n336), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n331), .A2(new_n333), .A3(new_n346), .A4(new_n332), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT74), .ZN(new_n348));
  AND3_X1   g147(.A1(new_n347), .A2(new_n348), .A3(KEYINPUT34), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n348), .B1(new_n347), .B2(KEYINPUT34), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n347), .A2(KEYINPUT34), .ZN(new_n351));
  NOR3_X1   g150(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n344), .A2(new_n345), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n352), .B1(new_n344), .B2(new_n345), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT35), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n328), .A2(new_n215), .ZN(new_n358));
  OR2_X1    g157(.A1(new_n358), .A2(KEYINPUT4), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n216), .A2(new_n236), .B1(new_n321), .B2(new_n323), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n360), .B1(new_n245), .B2(new_n243), .ZN(new_n361));
  OR3_X1    g160(.A1(new_n324), .A2(new_n215), .A3(KEYINPUT84), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT84), .B1(new_n324), .B2(new_n215), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n362), .A2(KEYINPUT4), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(G225gat), .A2(G233gat), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n366), .A2(KEYINPUT5), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n359), .A2(new_n361), .A3(new_n364), .A4(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n358), .A2(KEYINPUT4), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(new_n361), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n362), .A2(new_n363), .B1(KEYINPUT4), .B2(new_n365), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI22_X1  g171(.A1(new_n246), .A2(new_n324), .B1(new_n362), .B2(new_n363), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT5), .B1(new_n373), .B2(new_n365), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n368), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(KEYINPUT85), .B(KEYINPUT0), .Z(new_n376));
  XNOR2_X1  g175(.A(G1gat), .B(G29gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G57gat), .B(G85gat), .ZN(new_n379));
  XOR2_X1   g178(.A(new_n378), .B(new_n379), .Z(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT6), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n380), .B(new_n368), .C1(new_n372), .C2(new_n374), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n375), .A2(KEYINPUT6), .A3(new_n381), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AND2_X1   g186(.A1(new_n230), .A2(new_n233), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n309), .B1(new_n291), .B2(new_n297), .ZN(new_n389));
  NAND2_X1  g188(.A1(G226gat), .A2(G233gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(new_n234), .A3(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n391), .B1(new_n310), .B2(new_n390), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT79), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n393), .B(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n390), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n396), .B1(new_n310), .B2(new_n234), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT78), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n389), .A2(new_n396), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n400), .B1(new_n397), .B2(KEYINPUT78), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n238), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G8gat), .B(G36gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(G64gat), .ZN(new_n404));
  INV_X1    g203(.A(G92gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n404), .B(new_n405), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n395), .A2(new_n402), .A3(KEYINPUT30), .A4(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n406), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n393), .B(KEYINPUT79), .ZN(new_n409));
  INV_X1    g208(.A(new_n401), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n388), .B1(new_n410), .B2(new_n398), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n408), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n395), .A2(new_n402), .A3(new_n406), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT30), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n387), .A2(new_n407), .A3(new_n412), .A4(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n269), .A2(new_n356), .A3(new_n357), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n344), .A2(new_n345), .ZN(new_n419));
  INV_X1    g218(.A(new_n352), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n264), .A2(new_n421), .A3(new_n353), .A4(new_n267), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT35), .B1(new_n422), .B2(new_n416), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n418), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT91), .B(KEYINPUT38), .ZN(new_n425));
  AND2_X1   g224(.A1(new_n408), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT37), .B1(new_n395), .B2(new_n402), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT37), .B1(new_n388), .B2(new_n392), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n399), .A2(new_n401), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n428), .B1(new_n429), .B2(new_n388), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n426), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n431), .A2(new_n386), .A3(new_n385), .A4(new_n413), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT37), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n433), .B1(new_n409), .B2(new_n411), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n395), .A2(new_n402), .A3(KEYINPUT37), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n425), .B1(new_n436), .B2(new_n408), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n264), .B(new_n267), .C1(new_n432), .C2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT39), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n361), .B(new_n364), .C1(KEYINPUT4), .C2(new_n358), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n440), .A2(KEYINPUT88), .A3(new_n366), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT88), .B1(new_n440), .B2(new_n366), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n440), .A2(new_n366), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT88), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n440), .A2(KEYINPUT88), .A3(new_n366), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n439), .B1(new_n373), .B2(new_n365), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n443), .A2(new_n449), .A3(KEYINPUT40), .A4(new_n380), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n450), .B(KEYINPUT89), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n443), .A2(new_n449), .A3(new_n380), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT40), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n452), .A2(new_n453), .B1(new_n381), .B2(new_n375), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n415), .A2(new_n407), .A3(new_n412), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT90), .B1(new_n451), .B2(new_n456), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n449), .A2(new_n380), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n458), .A2(KEYINPUT89), .A3(KEYINPUT40), .A4(new_n443), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT89), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n450), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT90), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n462), .A2(new_n463), .A3(new_n455), .A4(new_n454), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n438), .B1(new_n457), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n268), .A2(new_n416), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT36), .B1(new_n354), .B2(new_n355), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT36), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n421), .A2(new_n468), .A3(new_n353), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n466), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n424), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT95), .ZN(new_n472));
  NAND2_X1  g271(.A1(G229gat), .A2(G233gat), .ZN(new_n473));
  XOR2_X1   g272(.A(new_n473), .B(KEYINPUT13), .Z(new_n474));
  AND2_X1   g273(.A1(G43gat), .A2(G50gat), .ZN(new_n475));
  NOR2_X1   g274(.A1(G43gat), .A2(G50gat), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT15), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(G43gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n258), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT15), .ZN(new_n480));
  NAND2_X1  g279(.A1(G43gat), .A2(G50gat), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(G29gat), .ZN(new_n484));
  INV_X1    g283(.A(G36gat), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(new_n485), .A3(KEYINPUT14), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT14), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n487), .B1(G29gat), .B2(G36gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(G29gat), .A2(G36gat), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n486), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT94), .B1(new_n483), .B2(new_n490), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n486), .A2(new_n488), .A3(new_n489), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT94), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n492), .A2(new_n493), .A3(new_n477), .A4(new_n482), .ZN(new_n494));
  INV_X1    g293(.A(new_n477), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n490), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n491), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(G1gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT16), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n254), .A2(G15gat), .ZN(new_n500));
  INV_X1    g299(.A(G15gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(G22gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n499), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(G1gat), .B1(new_n500), .B2(new_n502), .ZN(new_n505));
  OAI21_X1  g304(.A(G8gat), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n505), .ZN(new_n507));
  INV_X1    g306(.A(G8gat), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n507), .A2(new_n503), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n497), .A2(new_n510), .ZN(new_n511));
  AND2_X1   g310(.A1(G29gat), .A2(G36gat), .ZN(new_n512));
  NOR2_X1   g311(.A1(G29gat), .A2(G36gat), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n512), .B1(KEYINPUT14), .B2(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n514), .A2(new_n477), .A3(new_n482), .A4(new_n488), .ZN(new_n515));
  AOI22_X1  g314(.A1(new_n515), .A2(KEYINPUT94), .B1(new_n490), .B2(new_n495), .ZN(new_n516));
  AOI22_X1  g315(.A1(new_n516), .A2(new_n494), .B1(new_n506), .B2(new_n509), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n474), .B1(new_n511), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT12), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n520));
  XNOR2_X1  g319(.A(G169gat), .B(G197gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G113gat), .B(G141gat), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT93), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n522), .A2(new_n525), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n519), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n520), .B(new_n521), .Z(new_n530));
  XNOR2_X1  g329(.A(new_n523), .B(KEYINPUT93), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n532), .A2(KEYINPUT12), .A3(new_n526), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n497), .A2(new_n535), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n506), .A2(new_n509), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n516), .A2(KEYINPUT17), .A3(new_n494), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n497), .A2(new_n510), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n540), .A2(KEYINPUT18), .A3(new_n473), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n518), .B(new_n534), .C1(new_n539), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n473), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n536), .A2(new_n538), .A3(new_n537), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT18), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n472), .B1(new_n542), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT18), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n548), .B1(new_n539), .B2(new_n543), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n544), .A2(KEYINPUT18), .A3(new_n545), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n537), .A2(new_n494), .A3(new_n516), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(new_n540), .ZN(new_n552));
  AOI22_X1  g351(.A1(new_n552), .A2(new_n474), .B1(new_n529), .B2(new_n533), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n549), .A2(KEYINPUT95), .A3(new_n550), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n547), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n549), .A2(new_n550), .A3(new_n518), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n556), .A2(new_n533), .A3(new_n529), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n471), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G134gat), .B(G162gat), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G85gat), .A2(G92gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT7), .ZN(new_n563));
  XNOR2_X1  g362(.A(G99gat), .B(G106gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(G99gat), .A2(G106gat), .ZN(new_n565));
  INV_X1    g364(.A(G85gat), .ZN(new_n566));
  AOI22_X1  g365(.A1(KEYINPUT8), .A2(new_n565), .B1(new_n566), .B2(new_n405), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n563), .A2(new_n564), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n564), .B1(new_n563), .B2(new_n567), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n536), .A2(new_n538), .A3(new_n572), .ZN(new_n573));
  AND2_X1   g372(.A1(G232gat), .A2(G233gat), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n497), .A2(new_n571), .B1(KEYINPUT41), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT98), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT98), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n573), .A2(new_n578), .A3(new_n575), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n561), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n574), .A2(KEYINPUT41), .ZN(new_n582));
  XNOR2_X1  g381(.A(G190gat), .B(G218gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n577), .A2(new_n561), .A3(new_n579), .ZN(new_n585));
  AND3_X1   g384(.A1(new_n581), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n584), .B1(new_n581), .B2(new_n585), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G57gat), .B(G64gat), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  OR2_X1    g390(.A1(G71gat), .A2(G78gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(G71gat), .A2(G78gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT9), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n591), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n593), .B(new_n592), .C1(new_n590), .C2(new_n595), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n600), .A2(KEYINPUT21), .ZN(new_n601));
  XNOR2_X1  g400(.A(G127gat), .B(G155gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G183gat), .B(G211gat), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n603), .B(new_n604), .Z(new_n605));
  AOI21_X1  g404(.A(new_n510), .B1(new_n600), .B2(KEYINPUT21), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT97), .ZN(new_n607));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT96), .ZN(new_n609));
  XNOR2_X1  g408(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n607), .B(new_n611), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n605), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n605), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n599), .B1(new_n569), .B2(new_n570), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n563), .A2(new_n567), .ZN(new_n618));
  INV_X1    g417(.A(new_n564), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n620), .A2(new_n598), .A3(new_n597), .A4(new_n568), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT10), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n617), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n571), .A2(KEYINPUT10), .A3(new_n600), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G230gat), .A2(G233gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n617), .A2(new_n621), .ZN(new_n628));
  INV_X1    g427(.A(new_n626), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G120gat), .B(G148gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(G176gat), .ZN(new_n632));
  INV_X1    g431(.A(G204gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n627), .A2(new_n630), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(KEYINPUT99), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT99), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n627), .A2(new_n630), .A3(new_n637), .A4(new_n634), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n634), .B1(new_n627), .B2(new_n630), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(KEYINPUT100), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n640), .A2(KEYINPUT100), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n639), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n589), .A2(new_n616), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n559), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n387), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n455), .ZN(new_n652));
  NOR2_X1   g451(.A1(KEYINPUT101), .A2(KEYINPUT42), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT16), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  OR2_X1    g454(.A1(new_n655), .A2(G8gat), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n652), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n655), .A2(G8gat), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n656), .A2(new_n658), .A3(new_n659), .ZN(G1325gat));
  INV_X1    g459(.A(new_n648), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n467), .A2(KEYINPUT102), .A3(new_n469), .ZN(new_n662));
  AOI21_X1  g461(.A(KEYINPUT102), .B1(new_n467), .B2(new_n469), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(G15gat), .B1(new_n661), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n648), .A2(new_n501), .A3(new_n356), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(G1326gat));
  NAND2_X1  g466(.A1(new_n648), .A2(new_n268), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT43), .B(G22gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(G1327gat));
  NAND2_X1  g469(.A1(new_n615), .A2(new_n645), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n671), .A2(new_n589), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n559), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n673), .A2(new_n484), .A3(new_n649), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT45), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n471), .A2(KEYINPUT44), .A3(new_n588), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n555), .A2(KEYINPUT103), .A3(new_n557), .ZN(new_n677));
  AOI21_X1  g476(.A(KEYINPUT103), .B1(new_n555), .B2(new_n557), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n680), .A2(new_n671), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n457), .A2(new_n464), .ZN(new_n682));
  INV_X1    g481(.A(new_n438), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT104), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n268), .A2(new_n685), .A3(new_n416), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n685), .B1(new_n268), .B2(new_n416), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n664), .A2(new_n684), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n589), .B1(new_n690), .B2(new_n424), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n676), .B(new_n681), .C1(new_n691), .C2(KEYINPUT44), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n692), .A2(KEYINPUT105), .A3(new_n387), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT105), .B1(new_n692), .B2(new_n387), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(G29gat), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n675), .B1(new_n693), .B2(new_n695), .ZN(G1328gat));
  NAND3_X1  g495(.A1(new_n673), .A2(new_n485), .A3(new_n455), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n697), .B(KEYINPUT46), .Z(new_n698));
  INV_X1    g497(.A(new_n455), .ZN(new_n699));
  OAI21_X1  g498(.A(G36gat), .B1(new_n692), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(G1329gat));
  INV_X1    g500(.A(KEYINPUT47), .ZN(new_n702));
  OAI21_X1  g501(.A(G43gat), .B1(new_n692), .B2(new_n664), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n559), .A2(new_n478), .A3(new_n356), .A4(new_n672), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n704), .B(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n702), .A2(KEYINPUT106), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n707), .B1(new_n703), .B2(new_n708), .ZN(new_n709));
  OAI211_X1 g508(.A(KEYINPUT106), .B(G43gat), .C1(new_n692), .C2(new_n664), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n705), .B1(new_n709), .B2(new_n710), .ZN(G1330gat));
  OAI21_X1  g510(.A(G50gat), .B1(new_n692), .B2(new_n269), .ZN(new_n712));
  NOR2_X1   g511(.A1(KEYINPUT108), .A2(KEYINPUT48), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n269), .A2(G50gat), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n713), .B1(new_n673), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(KEYINPUT108), .A2(KEYINPUT48), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(G1331gat));
  INV_X1    g517(.A(new_n424), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n466), .A2(KEYINPUT104), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n686), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n721), .A2(new_n465), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n719), .B1(new_n722), .B2(new_n664), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n589), .A2(new_n616), .A3(new_n644), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n723), .A2(new_n679), .A3(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n387), .B(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g528(.A(KEYINPUT110), .B(G57gat), .Z(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1332gat));
  NAND2_X1  g530(.A1(new_n725), .A2(new_n455), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT49), .B(G64gat), .Z(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n732), .B2(new_n734), .ZN(G1333gat));
  INV_X1    g534(.A(KEYINPUT102), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n354), .A2(new_n355), .A3(KEYINPUT36), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n468), .B1(new_n421), .B2(new_n353), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n467), .A2(KEYINPUT102), .A3(new_n469), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n356), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(G71gat), .ZN(new_n744));
  AOI22_X1  g543(.A1(new_n742), .A2(G71gat), .B1(new_n725), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g545(.A1(new_n725), .A2(new_n268), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g547(.A1(new_n616), .A2(new_n679), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n644), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n676), .B(new_n751), .C1(new_n691), .C2(KEYINPUT44), .ZN(new_n752));
  OAI21_X1  g551(.A(G85gat), .B1(new_n752), .B2(new_n387), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n754));
  INV_X1    g553(.A(new_n749), .ZN(new_n755));
  NOR4_X1   g554(.A1(new_n723), .A2(new_n754), .A3(new_n589), .A4(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(KEYINPUT51), .B1(new_n691), .B2(new_n749), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n644), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n649), .A2(new_n566), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n753), .B1(new_n758), .B2(new_n759), .ZN(G1336gat));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n761));
  OAI21_X1  g560(.A(G92gat), .B1(new_n752), .B2(new_n699), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n699), .A2(G92gat), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n644), .B(new_n765), .C1(new_n756), .C2(new_n757), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n762), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n764), .B(new_n767), .ZN(G1337gat));
  INV_X1    g567(.A(G99gat), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n752), .A2(new_n769), .A3(new_n664), .ZN(new_n770));
  OR2_X1    g569(.A1(new_n758), .A2(new_n743), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(new_n771), .B2(new_n769), .ZN(G1338gat));
  OAI21_X1  g571(.A(G106gat), .B1(new_n752), .B2(new_n269), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT53), .B1(new_n773), .B2(KEYINPUT112), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n269), .A2(G106gat), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n644), .B(new_n775), .C1(new_n756), .C2(new_n757), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n773), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n776), .B(new_n773), .C1(KEYINPUT112), .C2(KEYINPUT53), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n778), .A2(new_n779), .ZN(G1339gat));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n625), .A2(new_n626), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n629), .B1(new_n623), .B2(new_n624), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n634), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n786), .B1(new_n627), .B2(KEYINPUT54), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n781), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n634), .B1(new_n783), .B2(new_n784), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n627), .A2(KEYINPUT54), .ZN(new_n790));
  OAI211_X1 g589(.A(KEYINPUT55), .B(new_n789), .C1(new_n790), .C2(new_n782), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n788), .A2(new_n639), .A3(new_n791), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n677), .A2(new_n678), .A3(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n473), .B1(new_n545), .B2(new_n540), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n552), .A2(new_n474), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n532), .B(new_n526), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n555), .A2(new_n796), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n797), .A2(new_n644), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n589), .B1(new_n793), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n792), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n588), .A2(new_n797), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n616), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n646), .A2(new_n679), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT113), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n678), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n555), .A2(KEYINPUT103), .A3(new_n557), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n805), .A2(new_n806), .A3(new_n800), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n797), .A2(new_n644), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n588), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n801), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n615), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n647), .A2(new_n680), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n804), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n815), .A2(new_n422), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n727), .A2(new_n455), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(G113gat), .B1(new_n818), .B2(new_n679), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n455), .A2(new_n387), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  XOR2_X1   g620(.A(new_n821), .B(KEYINPUT114), .Z(new_n822));
  INV_X1    g621(.A(new_n558), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(new_n311), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n819), .B1(new_n822), .B2(new_n824), .ZN(G1340gat));
  AOI21_X1  g624(.A(G120gat), .B1(new_n818), .B2(new_n644), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n645), .A2(new_n312), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n826), .B1(new_n822), .B2(new_n827), .ZN(G1341gat));
  INV_X1    g627(.A(new_n822), .ZN(new_n829));
  OAI21_X1  g628(.A(G127gat), .B1(new_n829), .B2(new_n615), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n818), .A2(new_n317), .A3(new_n616), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(G1342gat));
  OAI21_X1  g631(.A(G134gat), .B1(new_n829), .B2(new_n589), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n818), .A2(new_n315), .A3(new_n588), .ZN(new_n834));
  XOR2_X1   g633(.A(new_n834), .B(KEYINPUT56), .Z(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n836), .B(new_n837), .ZN(G1343gat));
  INV_X1    g637(.A(new_n815), .ZN(new_n839));
  AND4_X1   g638(.A1(new_n268), .A2(new_n664), .A3(new_n839), .A4(new_n817), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n823), .A2(G141gat), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT58), .ZN(new_n843));
  INV_X1    g642(.A(G141gat), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n268), .A2(KEYINPUT57), .ZN(new_n845));
  AOI22_X1  g644(.A1(new_n800), .A2(new_n558), .B1(new_n797), .B2(new_n644), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n801), .B1(new_n846), .B2(new_n588), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n803), .B1(new_n847), .B2(new_n615), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n804), .A2(new_n268), .A3(new_n814), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n739), .A2(new_n740), .A3(new_n820), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n852), .A2(new_n823), .A3(new_n853), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n842), .B(new_n843), .C1(new_n844), .C2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT118), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n850), .A2(new_n851), .ZN(new_n857));
  INV_X1    g656(.A(new_n849), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n853), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(KEYINPUT116), .A3(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n862), .B1(new_n852), .B2(new_n853), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n861), .A2(new_n679), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(G141gat), .ZN(new_n865));
  AOI22_X1  g664(.A1(new_n865), .A2(KEYINPUT117), .B1(new_n840), .B2(new_n841), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n864), .A2(new_n867), .A3(G141gat), .ZN(new_n868));
  AOI211_X1 g667(.A(new_n856), .B(new_n843), .C1(new_n866), .C2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n865), .A2(KEYINPUT117), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(new_n868), .A3(new_n842), .ZN(new_n871));
  AOI21_X1  g670(.A(KEYINPUT118), .B1(new_n871), .B2(KEYINPUT58), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n855), .B1(new_n869), .B2(new_n872), .ZN(G1344gat));
  NAND2_X1  g672(.A1(new_n840), .A2(new_n644), .ZN(new_n874));
  INV_X1    g673(.A(G148gat), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(KEYINPUT59), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n861), .A2(new_n644), .A3(new_n863), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n847), .A2(new_n615), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n646), .A2(new_n558), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n268), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n851), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n882), .B(new_n883), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n815), .A2(new_n845), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n645), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n853), .A2(new_n878), .ZN(new_n887));
  AOI22_X1  g686(.A1(new_n877), .A2(new_n878), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n876), .B1(new_n888), .B2(new_n875), .ZN(new_n889));
  XOR2_X1   g688(.A(new_n889), .B(KEYINPUT120), .Z(G1345gat));
  NAND3_X1  g689(.A1(new_n861), .A2(new_n616), .A3(new_n863), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n213), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n615), .A2(new_n213), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n840), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n894), .ZN(G1346gat));
  INV_X1    g694(.A(G162gat), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n840), .A2(new_n896), .A3(new_n588), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n861), .A2(new_n588), .A3(new_n863), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n897), .B1(new_n898), .B2(new_n896), .ZN(new_n899));
  XOR2_X1   g698(.A(new_n899), .B(KEYINPUT121), .Z(G1347gat));
  NAND3_X1  g699(.A1(new_n816), .A2(new_n455), .A3(new_n727), .ZN(new_n901));
  OAI21_X1  g700(.A(G169gat), .B1(new_n901), .B2(new_n823), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT122), .ZN(new_n903));
  NOR4_X1   g702(.A1(new_n815), .A2(new_n649), .A3(new_n699), .A4(new_n422), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(new_n282), .A3(new_n679), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(G1348gat));
  OAI21_X1  g705(.A(G176gat), .B1(new_n901), .B2(new_n645), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n904), .A2(new_n283), .A3(new_n644), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1349gat));
  OAI21_X1  g708(.A(G183gat), .B1(new_n901), .B2(new_n615), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n904), .A2(new_n303), .A3(new_n616), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT60), .ZN(new_n912));
  AOI22_X1  g711(.A1(new_n910), .A2(new_n911), .B1(KEYINPUT123), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n912), .A2(KEYINPUT123), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n913), .B(new_n914), .ZN(G1350gat));
  OAI21_X1  g714(.A(G190gat), .B1(new_n901), .B2(new_n589), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT61), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n904), .A2(new_n274), .A3(new_n588), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT124), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(G1351gat));
  NOR2_X1   g719(.A1(new_n815), .A2(new_n649), .ZN(new_n921));
  AND4_X1   g720(.A1(new_n455), .A2(new_n921), .A3(new_n664), .A4(new_n268), .ZN(new_n922));
  INV_X1    g721(.A(G197gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n922), .A2(new_n923), .A3(new_n679), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n884), .A2(new_n885), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n741), .A2(new_n699), .A3(new_n728), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n925), .B1(new_n928), .B2(new_n823), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(G197gat), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n928), .A2(new_n925), .A3(new_n823), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n924), .B1(new_n930), .B2(new_n931), .ZN(G1352gat));
  AOI21_X1  g731(.A(new_n633), .B1(new_n886), .B2(new_n927), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n922), .A2(new_n633), .A3(new_n644), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT126), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  XOR2_X1   g736(.A(new_n934), .B(KEYINPUT126), .Z(new_n938));
  AND3_X1   g737(.A1(new_n938), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n939));
  AOI21_X1  g738(.A(KEYINPUT127), .B1(new_n938), .B2(KEYINPUT62), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(G1353gat));
  NAND3_X1  g740(.A1(new_n922), .A2(new_n220), .A3(new_n616), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n926), .A2(new_n616), .A3(new_n927), .ZN(new_n943));
  AND3_X1   g742(.A1(new_n943), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n944));
  AOI21_X1  g743(.A(KEYINPUT63), .B1(new_n943), .B2(G211gat), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(G1354gat));
  NOR3_X1   g745(.A1(new_n928), .A2(new_n221), .A3(new_n589), .ZN(new_n947));
  AOI21_X1  g746(.A(G218gat), .B1(new_n922), .B2(new_n588), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n947), .A2(new_n948), .ZN(G1355gat));
endmodule


