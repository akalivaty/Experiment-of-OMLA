//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 1 0 1 1 0 1 0 1 1 0 0 1 1 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G58), .ZN(new_n209));
  INV_X1    g0009(.A(G232), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  OAI22_X1  g0012(.A1(new_n209), .A2(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n213), .B1(G107), .B2(G264), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  OAI22_X1  g0017(.A1(new_n202), .A2(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n218), .B1(G116), .B2(G270), .ZN(new_n219));
  AND2_X1   g0019(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  XNOR2_X1  g0021(.A(KEYINPUT64), .B(G238), .ZN(new_n222));
  INV_X1    g0022(.A(G257), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n205), .C2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G20), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT1), .Z(new_n227));
  NOR2_X1   g0027(.A1(new_n225), .A2(G13), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT0), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  INV_X1    g0031(.A(G20), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  INV_X1    g0034(.A(new_n201), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n235), .A2(G50), .ZN(new_n236));
  OAI211_X1 g0036(.A(new_n227), .B(new_n230), .C1(new_n234), .C2(new_n236), .ZN(new_n237));
  INV_X1    g0037(.A(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  INV_X1    g0043(.A(G264), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT65), .B(G270), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n242), .B(new_n247), .ZN(G358));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XOR2_X1   g0049(.A(G50), .B(G58), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n251), .B(KEYINPUT67), .Z(new_n252));
  XOR2_X1   g0052(.A(G87), .B(G97), .Z(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(KEYINPUT66), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G107), .B(G116), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n252), .B(new_n256), .ZN(G351));
  XNOR2_X1  g0057(.A(G58), .B(G68), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n258), .A2(G20), .B1(G159), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT3), .B(G33), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT7), .ZN(new_n262));
  NOR3_X1   g0062(.A1(new_n261), .A2(new_n262), .A3(G20), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G33), .ZN(new_n267));
  AOI21_X1  g0067(.A(G20), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(KEYINPUT75), .B1(new_n268), .B2(KEYINPUT7), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT75), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n270), .B(new_n262), .C1(new_n261), .C2(G20), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n263), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  OAI211_X1 g0072(.A(KEYINPUT16), .B(new_n260), .C1(new_n272), .C2(new_n221), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT16), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n262), .B1(new_n261), .B2(G20), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n265), .A2(new_n267), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(KEYINPUT7), .A3(new_n232), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n221), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n260), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n274), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n231), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n273), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT8), .B(G58), .ZN(new_n284));
  INV_X1    g0084(.A(G1), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G20), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n285), .A2(G13), .A3(G20), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(new_n282), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n288), .A2(new_n291), .B1(new_n290), .B2(new_n284), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n283), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G274), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(G1), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G45), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT69), .ZN(new_n297));
  XNOR2_X1  g0097(.A(KEYINPUT68), .B(G41), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n285), .A2(G274), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n296), .B(new_n297), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  AND2_X1   g0100(.A1(KEYINPUT68), .A2(G41), .ZN(new_n301));
  NOR2_X1   g0101(.A1(KEYINPUT68), .A2(G41), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI211_X1 g0103(.A(KEYINPUT69), .B(new_n295), .C1(new_n303), .C2(G45), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G41), .ZN(new_n306));
  OAI211_X1 g0106(.A(G1), .B(G13), .C1(new_n264), .C2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n215), .A2(G1698), .ZN(new_n309));
  OR2_X1    g0109(.A1(G223), .A2(G1698), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n261), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n264), .A2(new_n211), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n308), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n285), .B1(G41), .B2(G45), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n307), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G232), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n305), .A2(new_n313), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G169), .ZN(new_n319));
  INV_X1    g0119(.A(G179), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n319), .B1(new_n320), .B2(new_n318), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n293), .A2(new_n321), .A3(KEYINPUT18), .ZN(new_n322));
  AOI21_X1  g0122(.A(KEYINPUT18), .B1(new_n293), .B2(new_n321), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT17), .ZN(new_n326));
  INV_X1    g0126(.A(G190), .ZN(new_n327));
  OR2_X1    g0127(.A1(new_n318), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n318), .A2(G200), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n283), .A2(new_n328), .A3(new_n292), .A4(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT76), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n326), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  AND3_X1   g0132(.A1(new_n283), .A2(new_n292), .A3(new_n329), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n333), .A2(KEYINPUT76), .A3(KEYINPUT17), .A4(new_n328), .ZN(new_n334));
  INV_X1    g0134(.A(new_n259), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT15), .B(G87), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n264), .A2(G20), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  OAI22_X1  g0138(.A1(new_n335), .A2(new_n284), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n232), .A2(new_n216), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n282), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n341), .B(KEYINPUT71), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n291), .A2(G77), .A3(new_n286), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G1698), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G232), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n261), .B(new_n346), .C1(new_n222), .C2(new_n345), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n347), .B(new_n308), .C1(G107), .C2(new_n261), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n316), .A2(G244), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n305), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G190), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(G200), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n290), .A2(new_n216), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n344), .A2(new_n352), .A3(new_n353), .A4(new_n354), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n325), .A2(new_n332), .A3(new_n334), .A4(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n305), .B1(new_n215), .B2(new_n315), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT70), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n345), .A2(G222), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G223), .A2(G1698), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n261), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n362), .B(new_n308), .C1(G77), .C2(new_n261), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n305), .B(KEYINPUT70), .C1(new_n215), .C2(new_n315), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n359), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(G169), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n203), .A2(G20), .ZN(new_n368));
  INV_X1    g0168(.A(G150), .ZN(new_n369));
  OAI221_X1 g0169(.A(new_n368), .B1(new_n369), .B2(new_n335), .C1(new_n284), .C2(new_n338), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n282), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n290), .A2(new_n202), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n291), .A2(G50), .A3(new_n286), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n359), .A2(new_n320), .A3(new_n363), .A4(new_n364), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n367), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n365), .A2(G200), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT72), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT9), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n371), .A2(new_n372), .A3(new_n373), .A4(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n379), .A2(new_n380), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n382), .B(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n359), .A2(G190), .A3(new_n363), .A4(new_n364), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n378), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT10), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT10), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n378), .A2(new_n384), .A3(new_n388), .A4(new_n385), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n377), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n210), .A2(G1698), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n261), .B(new_n392), .C1(G226), .C2(G1698), .ZN(new_n393));
  NAND2_X1  g0193(.A1(G33), .A2(G97), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n308), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT13), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n316), .A2(G238), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n396), .A2(new_n305), .A3(new_n397), .A4(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G238), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n300), .B(new_n304), .C1(new_n400), .C2(new_n315), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n307), .B1(new_n393), .B2(new_n394), .ZN(new_n402));
  OAI21_X1  g0202(.A(KEYINPUT13), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(G169), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT14), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT14), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n404), .A2(new_n407), .A3(G169), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n406), .B(new_n408), .C1(new_n320), .C2(new_n404), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT73), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n290), .A2(new_n410), .A3(new_n221), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT73), .B1(new_n289), .B2(G68), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(KEYINPUT12), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n291), .A2(G68), .A3(new_n286), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT12), .ZN(new_n415));
  OAI211_X1 g0215(.A(KEYINPUT73), .B(new_n415), .C1(new_n289), .C2(G68), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n413), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  XNOR2_X1  g0217(.A(new_n417), .B(KEYINPUT74), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n337), .A2(G77), .B1(new_n259), .B2(G50), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n232), .B2(G68), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n282), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n421), .B(KEYINPUT11), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n409), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n404), .A2(new_n327), .ZN(new_n425));
  INV_X1    g0225(.A(G200), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n426), .B1(new_n399), .B2(new_n403), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n423), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n344), .A2(new_n354), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n350), .A2(new_n366), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n351), .A2(new_n320), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n424), .A2(new_n429), .A3(new_n433), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n356), .A2(new_n391), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n212), .A2(new_n345), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n223), .A2(G1698), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n265), .A2(new_n436), .A3(new_n267), .A4(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(G294), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n438), .B1(new_n264), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(G45), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n441), .A2(G1), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT5), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(new_n301), .B2(new_n302), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n444), .A2(new_n306), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n443), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n440), .A2(new_n308), .B1(new_n448), .B2(G274), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n445), .A2(new_n447), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n308), .B1(new_n450), .B2(new_n442), .ZN(new_n451));
  AOI21_X1  g0251(.A(KEYINPUT88), .B1(new_n451), .B2(G264), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT88), .ZN(new_n453));
  NOR4_X1   g0253(.A1(new_n448), .A2(new_n453), .A3(new_n244), .A4(new_n308), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n449), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G169), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n456), .B1(new_n320), .B2(new_n455), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT24), .ZN(new_n458));
  AND4_X1   g0258(.A1(new_n232), .A2(new_n265), .A3(new_n267), .A4(G87), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT22), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(KEYINPUT84), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT84), .ZN(new_n463));
  OAI21_X1  g0263(.A(KEYINPUT85), .B1(new_n463), .B2(KEYINPUT22), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT85), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n465), .A2(new_n460), .A3(KEYINPUT84), .ZN(new_n466));
  AND2_X1   g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n459), .A2(new_n462), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n464), .A2(new_n466), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n265), .A2(new_n267), .A3(new_n232), .A4(G87), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n469), .B1(new_n470), .B2(new_n461), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT23), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n473), .B1(new_n232), .B2(G107), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G116), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT78), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT78), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G116), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n476), .B1(new_n481), .B2(new_n338), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n458), .B1(new_n472), .B2(new_n483), .ZN(new_n484));
  AOI211_X1 g0284(.A(KEYINPUT24), .B(new_n482), .C1(new_n468), .C2(new_n471), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n282), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n290), .A2(new_n206), .B1(KEYINPUT86), .B2(KEYINPUT25), .ZN(new_n487));
  NOR2_X1   g0287(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n488));
  XNOR2_X1  g0288(.A(new_n487), .B(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n264), .A2(G1), .ZN(new_n490));
  NOR3_X1   g0290(.A1(new_n290), .A2(new_n282), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(G107), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n486), .A2(KEYINPUT87), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT87), .B1(new_n486), .B2(new_n494), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n457), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n455), .A2(G200), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n449), .B(G190), .C1(new_n452), .C2(new_n454), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n498), .A2(new_n486), .A3(new_n494), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G33), .A2(G283), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n501), .B(new_n232), .C1(G33), .C2(new_n205), .ZN(new_n502));
  XNOR2_X1  g0302(.A(KEYINPUT78), .B(G116), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n282), .B(new_n502), .C1(new_n503), .C2(new_n232), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT83), .ZN(new_n506));
  OR2_X1    g0306(.A1(new_n506), .A2(KEYINPUT20), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(KEYINPUT20), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n505), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n491), .A2(G116), .B1(new_n290), .B2(new_n481), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n504), .A2(new_n506), .A3(KEYINPUT20), .ZN(new_n511));
  AND3_X1   g0311(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n446), .B1(new_n298), .B2(new_n444), .ZN(new_n513));
  OAI211_X1 g0313(.A(G270), .B(new_n307), .C1(new_n513), .C2(new_n443), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n345), .A2(G257), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G264), .A2(G1698), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n261), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n517), .B(new_n308), .C1(G303), .C2(new_n261), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n448), .A2(G274), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n514), .A2(G179), .A3(new_n518), .A4(new_n519), .ZN(new_n520));
  OR2_X1    g0320(.A1(new_n512), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n514), .A2(new_n519), .A3(new_n518), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(G169), .A3(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT21), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n523), .A2(G200), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n512), .B(new_n527), .C1(new_n327), .C2(new_n523), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n522), .A2(new_n523), .A3(KEYINPUT21), .A4(G169), .ZN(new_n529));
  AND4_X1   g0329(.A1(new_n521), .A2(new_n526), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n497), .A2(new_n500), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n400), .A2(new_n345), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n217), .A2(G1698), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n265), .A2(new_n532), .A3(new_n267), .A4(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n478), .A2(new_n480), .A3(G33), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(KEYINPUT79), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT79), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n534), .A2(new_n538), .A3(new_n535), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n308), .A3(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n308), .A2(new_n442), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n541), .A2(G250), .B1(G45), .B2(new_n295), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n540), .A2(KEYINPUT80), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(KEYINPUT80), .B1(new_n540), .B2(new_n542), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n320), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n540), .A2(new_n542), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT80), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n540), .A2(KEYINPUT80), .A3(new_n542), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n548), .A2(new_n366), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n232), .A2(G33), .A3(G97), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT19), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT81), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n265), .A2(new_n267), .A3(new_n232), .A4(G68), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n232), .B1(new_n394), .B2(new_n552), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n211), .A2(new_n205), .A3(new_n206), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT81), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n551), .A2(new_n559), .A3(new_n552), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n554), .A2(new_n555), .A3(new_n558), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n282), .ZN(new_n562));
  INV_X1    g0362(.A(new_n336), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n491), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n336), .A2(new_n290), .ZN(new_n565));
  AND4_X1   g0365(.A1(KEYINPUT82), .A2(new_n562), .A3(new_n564), .A4(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n561), .A2(new_n282), .B1(new_n290), .B2(new_n336), .ZN(new_n567));
  AOI21_X1  g0367(.A(KEYINPUT82), .B1(new_n567), .B2(new_n564), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n545), .A2(new_n550), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(G190), .B1(new_n543), .B2(new_n544), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n548), .A2(G200), .A3(new_n549), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n491), .A2(G87), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n567), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n571), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n265), .A2(new_n267), .A3(G244), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT4), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n577), .A2(G1698), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n261), .A2(G244), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n580), .A3(new_n501), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n261), .A2(G250), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n345), .B1(new_n582), .B2(KEYINPUT4), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n308), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n451), .A2(G257), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n584), .A2(new_n585), .A3(new_n519), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n366), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n584), .A2(new_n320), .A3(new_n585), .A4(new_n519), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT77), .ZN(new_n589));
  NAND2_X1  g0389(.A1(KEYINPUT6), .A2(G97), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n589), .B1(new_n590), .B2(G107), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n206), .A2(KEYINPUT77), .A3(KEYINPUT6), .A4(G97), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(G97), .A2(G107), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT6), .B1(new_n207), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(G20), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n259), .A2(G77), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n206), .B1(new_n275), .B2(new_n277), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n282), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n289), .A2(G97), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n491), .A2(G97), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n587), .A2(new_n588), .A3(new_n604), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n586), .A2(G200), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n584), .A2(G190), .A3(new_n585), .A4(new_n519), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n570), .A2(new_n575), .A3(new_n605), .A4(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n531), .A2(new_n610), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n435), .A2(new_n611), .ZN(G372));
  NAND2_X1  g0412(.A1(new_n609), .A2(new_n605), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n521), .A2(new_n526), .A3(new_n529), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n486), .A2(new_n494), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n457), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n613), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n546), .A2(G200), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT89), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n546), .A2(KEYINPUT89), .A3(G200), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n571), .A2(new_n574), .A3(new_n621), .A4(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n546), .A2(new_n366), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n545), .A2(new_n569), .A3(new_n624), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n623), .A2(new_n500), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n618), .A2(new_n626), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n623), .A2(new_n625), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT90), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n604), .A2(new_n588), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n576), .A2(new_n577), .B1(G33), .B2(G283), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n577), .B1(new_n261), .B2(G250), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n631), .B(new_n580), .C1(new_n345), .C2(new_n632), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n633), .A2(new_n308), .B1(G257), .B2(new_n451), .ZN(new_n634));
  AOI21_X1  g0434(.A(G169), .B1(new_n634), .B2(new_n519), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n629), .B1(new_n630), .B2(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n587), .A2(KEYINPUT90), .A3(new_n588), .A4(new_n604), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n628), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n625), .ZN(new_n642));
  INV_X1    g0442(.A(new_n605), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n570), .A2(new_n575), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n642), .B1(new_n644), .B2(KEYINPUT26), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n627), .A2(new_n641), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n435), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n433), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n648), .A2(new_n429), .B1(new_n423), .B2(new_n409), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n334), .A2(new_n332), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n325), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n387), .A2(new_n389), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n377), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n647), .A2(new_n653), .ZN(G369));
  INV_X1    g0454(.A(G13), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(G20), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n285), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(G213), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(G343), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n512), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n614), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n530), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n665), .B1(new_n666), .B2(new_n664), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT91), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT91), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT92), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT92), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n668), .A2(new_n673), .A3(new_n670), .ZN(new_n674));
  INV_X1    g0474(.A(new_n500), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT87), .ZN(new_n676));
  INV_X1    g0476(.A(new_n282), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n467), .B1(new_n459), .B2(new_n462), .ZN(new_n678));
  NOR3_X1   g0478(.A1(new_n470), .A2(new_n469), .A3(new_n461), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n483), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(KEYINPUT24), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n472), .A2(new_n458), .A3(new_n483), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n677), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n676), .B1(new_n683), .B2(new_n493), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n486), .A2(KEYINPUT87), .A3(new_n494), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n675), .B1(new_n686), .B2(new_n457), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n662), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n686), .A2(new_n457), .A3(new_n662), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n672), .A2(G330), .A3(new_n674), .A4(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n614), .A2(new_n663), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n687), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n617), .A2(new_n662), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n692), .A2(new_n697), .ZN(G399));
  INV_X1    g0498(.A(new_n228), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(new_n303), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n557), .A2(G116), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(G1), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n236), .B2(new_n701), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT28), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT29), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n497), .A2(new_n615), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n613), .A2(KEYINPUT97), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT97), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n609), .A2(new_n605), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n707), .A2(new_n711), .A3(new_n626), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT98), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n623), .A2(new_n625), .ZN(new_n715));
  OAI21_X1  g0515(.A(KEYINPUT26), .B1(new_n715), .B2(new_n638), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n570), .A2(new_n575), .A3(new_n640), .A4(new_n643), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n716), .A2(new_n625), .A3(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n707), .A2(new_n711), .A3(KEYINPUT98), .A4(new_n626), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n714), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n706), .B1(new_n720), .B2(new_n663), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n646), .A2(new_n663), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(KEYINPUT29), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  AND4_X1   g0524(.A1(new_n570), .A2(new_n575), .A3(new_n605), .A4(new_n609), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n725), .A2(new_n687), .A3(new_n530), .A4(new_n663), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT96), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n497), .A2(new_n500), .A3(new_n530), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n729), .A2(KEYINPUT96), .A3(new_n725), .A4(new_n663), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT30), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n440), .A2(new_n308), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n519), .ZN(new_n734));
  OAI211_X1 g0534(.A(G264), .B(new_n307), .C1(new_n513), .C2(new_n443), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n453), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n451), .A2(KEYINPUT88), .A3(G264), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n734), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n634), .B(new_n738), .C1(new_n543), .C2(new_n544), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n520), .B(KEYINPUT94), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n732), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n738), .A2(G179), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n742), .A2(new_n546), .A3(new_n586), .A4(new_n523), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT94), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n520), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n584), .A2(new_n585), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n455), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n548), .A2(new_n549), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n745), .A2(new_n747), .A3(new_n748), .A4(KEYINPUT30), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n741), .A2(new_n743), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n662), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT31), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(KEYINPUT95), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT95), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n751), .A2(new_n755), .A3(new_n752), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  XOR2_X1   g0557(.A(KEYINPUT93), .B(KEYINPUT31), .Z(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n751), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n731), .A2(new_n757), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G330), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n724), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n705), .B1(new_n765), .B2(G1), .ZN(G364));
  AOI21_X1  g0566(.A(new_n231), .B1(G20), .B2(new_n366), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G179), .A2(G200), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT101), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G190), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G20), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n772), .A2(KEYINPUT102), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(KEYINPUT102), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n205), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n772), .A2(new_n769), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G159), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(KEYINPUT32), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n232), .A2(G179), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n781), .A2(new_n327), .A3(G200), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n206), .ZN(new_n783));
  NAND2_X1  g0583(.A1(G20), .A2(G179), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT99), .ZN(new_n785));
  AND3_X1   g0585(.A1(new_n785), .A2(new_n327), .A3(G200), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n781), .A2(G190), .A3(G200), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n786), .A2(G68), .B1(G87), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n785), .A2(G190), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n426), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n789), .B1(new_n202), .B2(new_n792), .ZN(new_n793));
  OR4_X1    g0593(.A1(new_n276), .A2(new_n780), .A3(new_n783), .A4(new_n793), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n776), .B(new_n794), .C1(KEYINPUT32), .C2(new_n779), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n790), .A2(G200), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n785), .A2(new_n327), .A3(new_n426), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(G58), .A2(new_n796), .B1(new_n798), .B2(G77), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT100), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(G326), .A2(new_n791), .B1(new_n798), .B2(G311), .ZN(new_n802));
  INV_X1    g0602(.A(G322), .ZN(new_n803));
  INV_X1    g0603(.A(new_n796), .ZN(new_n804));
  INV_X1    g0604(.A(new_n786), .ZN(new_n805));
  XOR2_X1   g0605(.A(KEYINPUT33), .B(G317), .Z(new_n806));
  OAI221_X1 g0606(.A(new_n802), .B1(new_n803), .B2(new_n804), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G303), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n276), .B1(new_n787), .B2(new_n808), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT103), .Z(new_n810));
  INV_X1    g0610(.A(G329), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n810), .B1(new_n439), .B2(new_n772), .C1(new_n777), .C2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n782), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n807), .B(new_n812), .C1(G283), .C2(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n767), .B1(new_n801), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n251), .A2(G45), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n699), .A2(new_n261), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n816), .B(new_n817), .C1(G45), .C2(new_n236), .ZN(new_n818));
  NAND3_X1  g0618(.A1(G355), .A2(new_n261), .A3(new_n228), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n818), .B(new_n819), .C1(G116), .C2(new_n228), .ZN(new_n820));
  NOR2_X1   g0620(.A1(G13), .A2(G33), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(G20), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(new_n767), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n815), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n672), .A2(new_n674), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n826), .B1(new_n827), .B2(new_n823), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n285), .B1(new_n656), .B2(G45), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n700), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n672), .A2(G330), .A3(new_n674), .ZN(new_n833));
  INV_X1    g0633(.A(new_n831), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(G330), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n827), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n832), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(G396));
  NOR2_X1   g0640(.A1(new_n433), .A2(new_n662), .ZN(new_n841));
  INV_X1    g0641(.A(new_n430), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n355), .B1(new_n842), .B2(new_n663), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n841), .B1(new_n843), .B2(new_n433), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n722), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n646), .A2(new_n844), .A3(new_n663), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n763), .B(new_n848), .Z(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n834), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n804), .A2(new_n439), .B1(new_n211), .B2(new_n782), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n851), .B(new_n776), .C1(G311), .C2(new_n778), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n261), .B1(new_n788), .B2(G107), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n791), .A2(G303), .B1(new_n786), .B2(G283), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n481), .B2(new_n797), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT104), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n855), .A2(new_n856), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n852), .A2(new_n853), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n796), .A2(G143), .B1(new_n786), .B2(G150), .ZN(new_n860));
  INV_X1    g0660(.A(G137), .ZN(new_n861));
  INV_X1    g0661(.A(G159), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n860), .B1(new_n861), .B2(new_n792), .C1(new_n862), .C2(new_n797), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT34), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n813), .A2(G68), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n772), .A2(new_n209), .B1(new_n202), .B2(new_n787), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n778), .B2(G132), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n864), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n859), .B1(new_n868), .B2(new_n276), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n834), .B1(new_n869), .B2(new_n767), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n767), .A2(new_n821), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n870), .B1(G77), .B2(new_n872), .C1(new_n822), .C2(new_n844), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n850), .A2(new_n873), .ZN(G384));
  NAND2_X1  g0674(.A1(new_n423), .A2(new_n662), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n424), .A2(new_n429), .A3(new_n875), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n423), .B(new_n662), .C1(new_n409), .C2(new_n428), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n844), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n751), .A2(new_n759), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n750), .A2(KEYINPUT31), .A3(new_n662), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n879), .B1(new_n731), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n260), .B1(new_n272), .B2(new_n221), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n274), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n885), .A2(new_n282), .A3(new_n273), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n660), .B1(new_n886), .B2(new_n292), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n650), .B2(new_n324), .ZN(new_n888));
  INV_X1    g0688(.A(new_n321), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n889), .A2(new_n660), .B1(new_n886), .B2(new_n292), .ZN(new_n890));
  INV_X1    g0690(.A(new_n330), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT37), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n293), .A2(new_n321), .ZN(new_n893));
  INV_X1    g0693(.A(new_n660), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n293), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT37), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n893), .A2(new_n895), .A3(new_n896), .A4(new_n330), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n892), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT38), .B1(new_n888), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n888), .A2(KEYINPUT38), .A3(new_n898), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n883), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT40), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n895), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n650), .B2(new_n324), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n893), .A2(new_n895), .A3(new_n330), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT37), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n897), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  XOR2_X1   g0711(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n901), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n883), .A2(KEYINPUT40), .A3(new_n914), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n905), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT106), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT96), .B1(new_n611), .B2(new_n663), .ZN(new_n918));
  NOR4_X1   g0718(.A1(new_n531), .A2(new_n610), .A3(new_n727), .A4(new_n662), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n882), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n435), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n917), .B(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(G330), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n435), .B1(new_n721), .B2(new_n723), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n653), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n900), .A2(KEYINPUT39), .A3(new_n901), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT39), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n888), .A2(KEYINPUT38), .A3(new_n898), .ZN(new_n928));
  INV_X1    g0728(.A(new_n912), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(new_n907), .B2(new_n910), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n927), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n424), .A2(new_n662), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n926), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n324), .A2(new_n660), .ZN(new_n934));
  INV_X1    g0734(.A(new_n878), .ZN(new_n935));
  INV_X1    g0735(.A(new_n841), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n935), .B1(new_n847), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n902), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n933), .A2(new_n934), .A3(new_n938), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n925), .B(new_n939), .Z(new_n940));
  XNOR2_X1  g0740(.A(new_n923), .B(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n285), .B2(new_n656), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n593), .A2(new_n595), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n477), .B1(new_n943), .B2(KEYINPUT35), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n944), .B(new_n233), .C1(KEYINPUT35), .C2(new_n943), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT36), .ZN(new_n946));
  OAI21_X1  g0746(.A(G77), .B1(new_n209), .B2(new_n221), .ZN(new_n947));
  OAI22_X1  g0747(.A1(new_n236), .A2(new_n947), .B1(G50), .B2(new_n221), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n948), .A2(G1), .A3(new_n655), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n942), .A2(new_n946), .A3(new_n949), .ZN(G367));
  NOR2_X1   g0750(.A1(new_n574), .A2(new_n663), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n642), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n715), .B2(new_n951), .ZN(new_n953));
  INV_X1    g0753(.A(new_n823), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n831), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(G283), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n804), .A2(new_n808), .B1(new_n956), .B2(new_n797), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n813), .A2(G97), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT46), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n787), .B2(new_n481), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NOR3_X1   g0761(.A1(new_n787), .A2(new_n959), .A3(new_n477), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n961), .A2(new_n261), .A3(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(G317), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n963), .B1(new_n206), .B2(new_n772), .C1(new_n777), .C2(new_n964), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n957), .B(new_n965), .C1(G311), .C2(new_n791), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n439), .B2(new_n805), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT109), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n775), .A2(new_n221), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n805), .A2(new_n862), .B1(new_n202), .B2(new_n797), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT110), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n261), .B1(new_n209), .B2(new_n787), .C1(new_n804), .C2(new_n369), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n791), .A2(G143), .B1(G77), .B2(new_n813), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n777), .B2(new_n861), .ZN(new_n974));
  OR4_X1    g0774(.A1(new_n969), .A2(new_n971), .A3(new_n972), .A4(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n968), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT111), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT47), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n955), .B1(new_n978), .B2(new_n767), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n247), .A2(new_n817), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n980), .B(new_n824), .C1(new_n228), .C2(new_n336), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(KEYINPUT108), .Z(new_n982));
  NAND2_X1  g0782(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n692), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n708), .A2(new_n710), .B1(new_n604), .B2(new_n662), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n605), .A2(new_n663), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n697), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT45), .ZN(new_n990));
  INV_X1    g0790(.A(new_n697), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT107), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT44), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n991), .A2(new_n992), .A3(new_n993), .A4(new_n987), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n992), .A2(new_n993), .ZN(new_n995));
  NAND2_X1  g0795(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n995), .B(new_n996), .C1(new_n697), .C2(new_n988), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n984), .B1(new_n990), .B2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT45), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n989), .B(new_n1000), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n1001), .A2(new_n692), .A3(new_n994), .A4(new_n997), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n695), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n691), .B2(new_n694), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n833), .B(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n765), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n700), .B(KEYINPUT41), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n830), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n692), .A2(new_n987), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n953), .A2(KEYINPUT43), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n695), .A2(new_n985), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT42), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n985), .A2(new_n686), .A3(new_n457), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n662), .B1(new_n1014), .B2(new_n605), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1011), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1010), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1010), .A2(new_n1016), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n953), .A2(KEYINPUT43), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1017), .A2(new_n1020), .A3(new_n1018), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n983), .B1(new_n1009), .B2(new_n1024), .ZN(G387));
  AOI21_X1  g0825(.A(new_n701), .B1(new_n1006), .B2(new_n764), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n764), .B2(new_n1006), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n778), .A2(G326), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n796), .A2(G317), .B1(new_n786), .B2(G311), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n808), .B2(new_n797), .C1(new_n803), .C2(new_n792), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT48), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n1031), .B1(new_n956), .B2(new_n772), .C1(new_n439), .C2(new_n787), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT49), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n261), .B(new_n1028), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n1033), .B2(new_n1032), .C1(new_n481), .C2(new_n782), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n775), .A2(new_n336), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n958), .B1(new_n202), .B2(new_n804), .C1(new_n777), .C2(new_n369), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n791), .A2(G159), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT112), .ZN(new_n1039));
  NOR3_X1   g0839(.A1(new_n1036), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n805), .A2(new_n284), .B1(new_n221), .B2(new_n797), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT113), .Z(new_n1042));
  OAI211_X1 g0842(.A(new_n1040), .B(new_n1042), .C1(new_n216), .C2(new_n787), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1035), .B1(new_n276), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n834), .B1(new_n1044), .B2(new_n767), .ZN(new_n1045));
  OR3_X1    g0845(.A1(new_n284), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1046));
  OAI21_X1  g0846(.A(KEYINPUT50), .B1(new_n284), .B2(G50), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1046), .A2(new_n1047), .A3(new_n441), .A4(new_n702), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(G68), .B2(G77), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n242), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n817), .B1(new_n1050), .B2(new_n441), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n261), .B(new_n228), .C1(G116), .C2(new_n557), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1049), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n228), .A2(G107), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n824), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1045), .B(new_n1055), .C1(new_n691), .C2(new_n954), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1027), .B(new_n1056), .C1(new_n829), .C2(new_n1006), .ZN(G393));
  AND2_X1   g0857(.A1(new_n999), .A2(new_n1002), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1006), .A2(new_n764), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1003), .B1(new_n764), .B2(new_n1006), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1060), .A2(new_n1061), .A3(new_n700), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1058), .A2(new_n830), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n772), .A2(new_n481), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n783), .B1(new_n798), .B2(G294), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1065), .B(new_n276), .C1(new_n956), .C2(new_n787), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1064), .B(new_n1066), .C1(G322), .C2(new_n778), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G311), .A2(new_n796), .B1(new_n791), .B2(G317), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT52), .Z(new_n1069));
  OAI211_X1 g0869(.A(new_n1067), .B(new_n1069), .C1(new_n808), .C2(new_n805), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n782), .A2(new_n211), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G150), .A2(new_n791), .B1(new_n796), .B2(G159), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n261), .B1(new_n221), .B2(new_n787), .C1(new_n1072), .C2(KEYINPUT51), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1071), .B(new_n1073), .C1(G143), .C2(new_n778), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(KEYINPUT51), .ZN(new_n1075));
  OAI21_X1  g0875(.A(G77), .B1(new_n774), .B2(new_n773), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n805), .A2(new_n202), .B1(new_n284), .B2(new_n797), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT114), .Z(new_n1079));
  OAI21_X1  g0879(.A(new_n1070), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n767), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n817), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n824), .B1(new_n205), .B2(new_n228), .C1(new_n256), .C2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1081), .A2(new_n831), .A3(new_n1083), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT115), .Z(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n954), .B2(new_n988), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1062), .A2(new_n1063), .A3(new_n1086), .ZN(G390));
  NAND2_X1  g0887(.A1(new_n844), .A2(G330), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n920), .A2(new_n878), .A3(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1090), .A2(KEYINPUT116), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n932), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n914), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n843), .A2(new_n433), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n720), .A2(new_n663), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n936), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1093), .B1(new_n1096), .B2(new_n878), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n847), .A2(new_n936), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n878), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n1099), .A2(new_n1092), .B1(new_n926), .B2(new_n931), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1091), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n920), .A2(KEYINPUT116), .A3(new_n1089), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n760), .B1(new_n754), .B2(new_n756), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1088), .B1(new_n1103), .B2(new_n731), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1102), .A2(new_n878), .A3(new_n1104), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n928), .A2(new_n899), .A3(new_n927), .ZN(new_n1106));
  AOI21_X1  g0906(.A(KEYINPUT39), .B1(new_n913), .B2(new_n901), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n1106), .A2(new_n1107), .B1(new_n937), .B2(new_n932), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n935), .B1(new_n1095), .B2(new_n936), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1105), .B(new_n1108), .C1(new_n1109), .C2(new_n1093), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1101), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n920), .A2(new_n435), .A3(G330), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n924), .A2(new_n653), .A3(new_n1112), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n728), .A2(new_n730), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n755), .B1(new_n751), .B2(new_n752), .ZN(new_n1115));
  AOI211_X1 g0915(.A(KEYINPUT95), .B(KEYINPUT31), .C1(new_n750), .C2(new_n662), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n761), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1089), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n935), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1119), .A2(new_n1090), .B1(new_n936), .B2(new_n847), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n935), .B(new_n1088), .C1(new_n1103), .C2(new_n731), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n878), .B1(new_n920), .B2(new_n1089), .ZN(new_n1122));
  NOR3_X1   g0922(.A1(new_n1121), .A2(new_n1122), .A3(new_n1096), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1113), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1111), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n878), .B1(new_n762), .B2(new_n1089), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n880), .A2(new_n881), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(new_n728), .B2(new_n730), .ZN(new_n1128));
  NOR3_X1   g0928(.A1(new_n1128), .A2(new_n935), .A3(new_n1088), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1098), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1095), .A2(new_n936), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n878), .B(new_n1089), .C1(new_n1114), .C2(new_n1117), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n935), .B1(new_n1128), .B2(new_n1088), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1130), .A2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1101), .A2(new_n1135), .A3(new_n1110), .A4(new_n1113), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1125), .A2(new_n700), .A3(new_n1136), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n1101), .A2(new_n1110), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n830), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n821), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n787), .A2(new_n369), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT118), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT53), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(G128), .A2(new_n791), .B1(new_n796), .B2(G132), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1144), .B1(new_n861), .B2(new_n805), .ZN(new_n1145));
  XOR2_X1   g0945(.A(KEYINPUT54), .B(G143), .Z(new_n1146));
  AOI21_X1  g0946(.A(new_n276), .B1(new_n798), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(G125), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1147), .B1(new_n777), .B2(new_n1148), .ZN(new_n1149));
  NOR3_X1   g0949(.A1(new_n1143), .A2(new_n1145), .A3(new_n1149), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1150), .B1(new_n202), .B2(new_n782), .C1(new_n862), .C2(new_n775), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1151), .B(KEYINPUT119), .Z(new_n1152));
  OAI21_X1  g0952(.A(new_n865), .B1(new_n777), .B2(new_n439), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT120), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n276), .B1(new_n805), .B2(new_n206), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n477), .A2(new_n804), .B1(new_n792), .B2(new_n956), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1155), .B(new_n1156), .C1(G87), .C2(new_n788), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1154), .A2(new_n1076), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(G97), .B2(new_n798), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n767), .B1(new_n1152), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n834), .B1(new_n284), .B2(new_n871), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n1161), .B(KEYINPUT117), .Z(new_n1162));
  NAND3_X1  g0962(.A1(new_n1140), .A2(new_n1160), .A3(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1137), .A2(new_n1139), .A3(new_n1163), .ZN(G378));
  INV_X1    g0964(.A(G124), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n264), .B(new_n306), .C1(new_n777), .C2(new_n1165), .ZN(new_n1166));
  AND2_X1   g0966(.A1(new_n786), .A2(G132), .ZN(new_n1167));
  INV_X1    g0967(.A(G128), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n1148), .A2(new_n792), .B1(new_n804), .B2(new_n1168), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1167), .B(new_n1169), .C1(new_n788), .C2(new_n1146), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1170), .B1(new_n861), .B2(new_n797), .C1(new_n369), .C2(new_n775), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1166), .B1(new_n1171), .B2(KEYINPUT59), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1172), .B1(KEYINPUT59), .B2(new_n1171), .C1(new_n862), .C2(new_n782), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n303), .A2(new_n261), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1173), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n796), .A2(G107), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n798), .A2(new_n563), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n786), .A2(G97), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1177), .A2(new_n1178), .A3(new_n1174), .A4(new_n1179), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n782), .A2(new_n209), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n791), .A2(G116), .B1(G77), .B2(new_n788), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n777), .B2(new_n956), .ZN(new_n1183));
  NOR4_X1   g0983(.A1(new_n969), .A2(new_n1180), .A3(new_n1181), .A4(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT58), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n767), .B1(new_n1176), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(new_n831), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT121), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n390), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n390), .A2(new_n1190), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n374), .A2(new_n894), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  NOR3_X1   g0995(.A1(new_n1192), .A2(new_n1193), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n391), .A2(KEYINPUT121), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1194), .B1(new_n1197), .B2(new_n1191), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1189), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1195), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1197), .A2(new_n1191), .A3(new_n1194), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1200), .A2(new_n1188), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1199), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1204), .A2(new_n822), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1187), .B(new_n1205), .C1(new_n202), .C2(new_n871), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n928), .A2(new_n899), .ZN(new_n1207));
  NOR3_X1   g1007(.A1(new_n1207), .A2(new_n1128), .A3(new_n879), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n915), .B(G330), .C1(new_n1208), .C2(KEYINPUT40), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n1204), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n939), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n905), .A2(new_n1203), .A3(G330), .A4(new_n915), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1211), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1206), .B1(new_n1215), .B2(new_n830), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n924), .A2(new_n653), .A3(new_n1112), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT122), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n924), .A2(KEYINPUT122), .A3(new_n653), .A4(new_n1112), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1136), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1215), .A2(KEYINPUT57), .A3(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n700), .ZN(new_n1223));
  AOI21_X1  g1023(.A(KEYINPUT57), .B1(new_n1215), .B2(new_n1221), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1216), .B1(new_n1223), .B2(new_n1224), .ZN(G375));
  NAND3_X1  g1025(.A1(new_n1217), .A2(new_n1130), .A3(new_n1134), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT123), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1217), .A2(new_n1130), .A3(new_n1134), .A4(KEYINPUT123), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1230), .A2(new_n1008), .A3(new_n1124), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n261), .B1(new_n862), .B2(new_n787), .C1(new_n777), .C2(new_n1168), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n1181), .B(new_n1232), .C1(G150), .C2(new_n798), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n791), .A2(G132), .B1(new_n786), .B2(new_n1146), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n1235), .B1(new_n202), .B2(new_n775), .C1(new_n861), .C2(new_n804), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1036), .B1(G283), .B2(new_n796), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1237), .B(KEYINPUT125), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n786), .A2(new_n503), .B1(G97), .B2(new_n788), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1239), .B1(new_n206), .B2(new_n797), .C1(new_n439), .C2(new_n792), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(G303), .B2(new_n778), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n276), .B1(new_n782), .B2(new_n216), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1242), .B(KEYINPUT124), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1238), .A2(new_n1241), .A3(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1236), .A2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n834), .B1(new_n1245), .B2(new_n767), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n871), .A2(new_n221), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n935), .A2(new_n821), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1090), .B1(new_n1104), .B2(new_n878), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1250), .A2(new_n1131), .B1(new_n1251), .B2(new_n1098), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1249), .B1(new_n1252), .B2(new_n829), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1231), .A2(new_n1254), .ZN(G381));
  INV_X1    g1055(.A(KEYINPUT57), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1214), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1252), .A2(new_n1217), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1260), .B1(new_n1138), .B2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1256), .B1(new_n1259), .B2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1263), .A2(new_n700), .A3(new_n1222), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1205), .A2(new_n1187), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(G50), .B2(new_n872), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1266), .B1(new_n1259), .B2(new_n829), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1267), .A2(G378), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1264), .A2(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1269), .A2(G381), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n982), .ZN(new_n1271));
  AOI211_X1 g1071(.A(new_n955), .B(new_n1271), .C1(new_n978), .C2(new_n767), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n829), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1024), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1272), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  NOR4_X1   g1076(.A1(G390), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1270), .A2(new_n1276), .A3(new_n1277), .ZN(G407));
  OAI211_X1 g1078(.A(G407), .B(G213), .C1(G343), .C2(new_n1269), .ZN(G409));
  INV_X1    g1079(.A(KEYINPUT126), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(new_n1276), .B2(G390), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(G393), .B(new_n839), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1276), .A2(G390), .ZN(new_n1283));
  INV_X1    g1083(.A(G390), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1284), .A2(G387), .ZN(new_n1285));
  OAI22_X1  g1085(.A1(new_n1281), .A2(new_n1282), .B1(new_n1283), .B2(new_n1285), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(G396), .B(G393), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1276), .A2(G390), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1284), .A2(G387), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1287), .A2(new_n1288), .A3(new_n1280), .A4(new_n1289), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1286), .A2(new_n1290), .A3(KEYINPUT127), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT127), .B1(new_n1286), .B2(new_n1290), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT61), .ZN(new_n1294));
  INV_X1    g1094(.A(G378), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1295), .B1(new_n1264), .B2(new_n1216), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1137), .A2(new_n1163), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1215), .A2(new_n1008), .A3(new_n1221), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1297), .A2(new_n1216), .A3(new_n1139), .A4(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n661), .A2(G213), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(G384), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT60), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1226), .A2(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(KEYINPUT60), .B1(new_n1252), .B2(new_n1217), .ZN(new_n1305));
  AOI211_X1 g1105(.A(new_n701), .B(new_n1304), .C1(new_n1230), .C2(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1302), .B1(new_n1306), .B2(new_n1253), .ZN(new_n1307));
  AOI21_X1  g1107(.A(KEYINPUT123), .B1(new_n1252), .B2(new_n1217), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1229), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1305), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1304), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1310), .A2(new_n700), .A3(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1312), .A2(G384), .A3(new_n1254), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1307), .A2(new_n1313), .ZN(new_n1314));
  NOR3_X1   g1114(.A1(new_n1296), .A2(new_n1301), .A3(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT62), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1294), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n661), .A2(G213), .A3(G2897), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1304), .B1(new_n1230), .B2(new_n1305), .ZN(new_n1320));
  AOI211_X1 g1120(.A(new_n1302), .B(new_n1253), .C1(new_n1320), .C2(new_n700), .ZN(new_n1321));
  AOI21_X1  g1121(.A(G384), .B1(new_n1312), .B2(new_n1254), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1319), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1307), .A2(new_n1313), .A3(new_n1318), .ZN(new_n1324));
  OAI211_X1 g1124(.A(new_n1323), .B(new_n1324), .C1(new_n1296), .C2(new_n1301), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(G375), .A2(G378), .ZN(new_n1326));
  AOI22_X1  g1126(.A1(new_n1268), .A2(new_n1298), .B1(G213), .B2(new_n661), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1326), .A2(new_n1327), .A3(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(KEYINPUT62), .B1(new_n1325), .B2(new_n1329), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1293), .B1(new_n1317), .B2(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(KEYINPUT61), .B1(new_n1286), .B2(new_n1290), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1315), .A2(KEYINPUT63), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT63), .ZN(new_n1334));
  NOR3_X1   g1134(.A1(new_n1321), .A2(new_n1322), .A3(new_n1319), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1318), .B1(new_n1307), .B2(new_n1313), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1334), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1339));
  OAI211_X1 g1139(.A(new_n1332), .B(new_n1333), .C1(new_n1339), .C2(new_n1315), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1331), .A2(new_n1340), .ZN(G405));
  INV_X1    g1141(.A(new_n1269), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1328), .B1(new_n1342), .B2(new_n1296), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1326), .A2(new_n1269), .A3(new_n1314), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1286), .A2(new_n1290), .ZN(new_n1346));
  XNOR2_X1  g1146(.A(new_n1345), .B(new_n1346), .ZN(G402));
endmodule


