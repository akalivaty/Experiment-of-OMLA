//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT9), .B(G234), .Z(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n187), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(G110), .B(G140), .ZN(new_n192));
  INV_X1    g006(.A(G953), .ZN(new_n193));
  AND2_X1   g007(.A1(new_n193), .A2(G227), .ZN(new_n194));
  XOR2_X1   g008(.A(new_n192), .B(new_n194), .Z(new_n195));
  INV_X1    g009(.A(G137), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G134), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(G134), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n197), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(KEYINPUT65), .A2(G137), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g016(.A1(KEYINPUT65), .A2(G137), .ZN(new_n203));
  OAI211_X1 g017(.A(KEYINPUT11), .B(G134), .C1(new_n202), .C2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G131), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n200), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n205), .B1(new_n200), .B2(new_n204), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT77), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n200), .A2(new_n204), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G131), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT77), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(new_n206), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n209), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT10), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(KEYINPUT64), .A3(G143), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n218));
  INV_X1    g032(.A(G143), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n218), .B1(new_n219), .B2(G146), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n219), .A2(G146), .ZN(new_n221));
  OAI211_X1 g035(.A(G128), .B(new_n217), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT1), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT1), .B1(new_n219), .B2(G146), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT75), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI211_X1 g041(.A(KEYINPUT75), .B(KEYINPUT1), .C1(new_n219), .C2(G146), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(G128), .A3(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n217), .B1(new_n220), .B2(new_n221), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n223), .A2(new_n224), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G104), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT3), .B1(new_n232), .B2(G107), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n234));
  INV_X1    g048(.A(G107), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n235), .A3(G104), .ZN(new_n236));
  INV_X1    g050(.A(G101), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n232), .A2(G107), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n233), .A2(new_n236), .A3(new_n237), .A4(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n235), .A2(G104), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n232), .A2(G107), .ZN(new_n241));
  OAI21_X1  g055(.A(G101), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n215), .B1(new_n231), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G128), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n216), .A2(G143), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n245), .B1(new_n246), .B2(new_n221), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n222), .A2(KEYINPUT0), .A3(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(G128), .B1(new_n246), .B2(new_n221), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT0), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n233), .A2(new_n236), .A3(new_n238), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n254), .A3(G101), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(G101), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(KEYINPUT4), .A3(new_n239), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n252), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT64), .B1(new_n216), .B2(G143), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n216), .A2(G143), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n261), .A2(new_n224), .A3(G128), .A4(new_n217), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n224), .B1(G143), .B2(new_n216), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n246), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n262), .A2(new_n264), .A3(new_n247), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT76), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n239), .A2(new_n242), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n266), .B1(new_n239), .B2(new_n242), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n265), .B(KEYINPUT10), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n214), .A2(new_n244), .A3(new_n258), .A4(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n244), .A2(new_n258), .A3(new_n269), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT79), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n211), .A2(new_n206), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n272), .B1(new_n271), .B2(new_n273), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n195), .B(new_n270), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n263), .A2(KEYINPUT75), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n228), .A2(G128), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n230), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n262), .ZN(new_n280));
  INV_X1    g094(.A(new_n243), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n243), .A2(new_n262), .A3(new_n264), .A4(new_n247), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT78), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT12), .B1(new_n284), .B2(new_n273), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT78), .ZN(new_n286));
  AND4_X1   g100(.A1(new_n243), .A2(new_n262), .A3(new_n264), .A4(new_n247), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n243), .B1(new_n279), .B2(new_n262), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n286), .B(new_n273), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT12), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n270), .B1(new_n285), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n195), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT80), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n276), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n295), .B1(new_n276), .B2(new_n294), .ZN(new_n298));
  INV_X1    g112(.A(G469), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  XOR2_X1   g114(.A(KEYINPUT70), .B(G902), .Z(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n248), .A2(new_n251), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n257), .A2(new_n255), .ZN(new_n304));
  OAI22_X1  g118(.A1(new_n303), .A2(new_n304), .B1(new_n288), .B2(KEYINPUT10), .ZN(new_n305));
  INV_X1    g119(.A(new_n269), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n273), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT79), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n195), .B1(new_n310), .B2(new_n270), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n292), .A2(new_n293), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n299), .B(new_n302), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n299), .A2(new_n189), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n191), .B1(new_n300), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT81), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n276), .A2(new_n294), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT80), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(G469), .A3(new_n296), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n322), .A2(new_n313), .A3(new_n315), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(KEYINPUT81), .A3(new_n191), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT89), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n326), .B1(new_n219), .B2(G128), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n245), .A2(KEYINPUT89), .A3(G143), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n219), .A2(G128), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT91), .ZN(new_n332));
  AOI22_X1  g146(.A1(new_n327), .A2(new_n328), .B1(G128), .B2(new_n219), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT91), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G134), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G116), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT87), .B1(new_n339), .B2(G122), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT87), .ZN(new_n341));
  INV_X1    g155(.A(G122), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n342), .A3(G116), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n339), .A2(G122), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(KEYINPUT14), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n347), .A3(G107), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n332), .A2(G134), .A3(new_n335), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n344), .B(new_n345), .C1(KEYINPUT14), .C2(new_n235), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n338), .A2(new_n348), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  OR2_X1    g165(.A1(KEYINPUT88), .A2(KEYINPUT13), .ZN(new_n352));
  NAND2_X1  g166(.A1(KEYINPUT88), .A2(KEYINPUT13), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n329), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n333), .B1(new_n354), .B2(G134), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n352), .A2(new_n353), .ZN(new_n356));
  AND4_X1   g170(.A1(G134), .A2(new_n329), .A3(new_n330), .A4(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n346), .A2(G107), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n235), .B1(new_n344), .B2(new_n345), .ZN(new_n359));
  OAI22_X1  g173(.A1(new_n355), .A2(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n360), .A2(KEYINPUT90), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT90), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n356), .B1(new_n327), .B2(new_n328), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n331), .B1(new_n363), .B2(new_n337), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n354), .A2(G134), .A3(new_n333), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n346), .B(G107), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n362), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n351), .B1(new_n361), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n188), .A2(G217), .A3(new_n193), .ZN(new_n370));
  XOR2_X1   g184(.A(new_n370), .B(KEYINPUT92), .Z(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n360), .A2(KEYINPUT90), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n366), .A2(new_n362), .A3(new_n367), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(new_n351), .A3(new_n371), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n373), .A2(new_n302), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(KEYINPUT93), .ZN(new_n379));
  INV_X1    g193(.A(G478), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n380), .A2(KEYINPUT15), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT93), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n373), .A2(new_n382), .A3(new_n302), .A4(new_n377), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n379), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n378), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n385), .B1(KEYINPUT15), .B2(new_n380), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G237), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(new_n193), .A3(G214), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n219), .ZN(new_n391));
  NOR2_X1   g205(.A1(G237), .A2(G953), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(G143), .A3(G214), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n205), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT18), .ZN(new_n395));
  XNOR2_X1  g209(.A(G125), .B(G140), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(new_n216), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n391), .A2(new_n393), .ZN(new_n398));
  AND2_X1   g212(.A1(KEYINPUT18), .A2(G131), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n395), .B(new_n397), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n393), .ZN(new_n401));
  AOI21_X1  g215(.A(G143), .B1(new_n392), .B2(G214), .ZN(new_n402));
  OAI21_X1  g216(.A(G131), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT17), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n391), .A2(new_n205), .A3(new_n393), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n394), .A2(KEYINPUT17), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G125), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n409), .A2(KEYINPUT16), .A3(G140), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n410), .B1(new_n396), .B2(KEYINPUT16), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT72), .B1(new_n411), .B2(G146), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(G146), .ZN(new_n413));
  INV_X1    g227(.A(new_n410), .ZN(new_n414));
  AND2_X1   g228(.A1(G125), .A2(G140), .ZN(new_n415));
  NOR2_X1   g229(.A1(G125), .A2(G140), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT16), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT72), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n419), .A3(new_n216), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n412), .A2(new_n413), .A3(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n400), .B1(new_n408), .B2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(G113), .B(G122), .ZN(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT84), .B(G104), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n423), .B(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n400), .B(new_n425), .C1(new_n408), .C2(new_n421), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n189), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT86), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT86), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n432), .B(new_n189), .C1(new_n427), .C2(new_n429), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n431), .A2(G475), .A3(new_n433), .ZN(new_n434));
  XOR2_X1   g248(.A(new_n396), .B(KEYINPUT19), .Z(new_n435));
  OAI21_X1  g249(.A(new_n413), .B1(new_n435), .B2(G146), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n403), .A2(new_n405), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n400), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n426), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n428), .ZN(new_n440));
  NOR2_X1   g254(.A1(G475), .A2(G902), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT20), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n439), .A2(KEYINPUT85), .A3(new_n428), .ZN(new_n445));
  AOI21_X1  g259(.A(KEYINPUT85), .B1(new_n439), .B2(new_n428), .ZN(new_n446));
  OAI211_X1 g260(.A(KEYINPUT20), .B(new_n441), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n434), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G952), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n449), .A2(G953), .ZN(new_n450));
  NAND2_X1  g264(.A1(G234), .A2(G237), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n301), .A2(G953), .A3(new_n451), .ZN(new_n453));
  XOR2_X1   g267(.A(KEYINPUT21), .B(G898), .Z(new_n454));
  OAI21_X1  g268(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(G214), .B1(G237), .B2(G902), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n456), .B(KEYINPUT82), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n252), .A2(G125), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n265), .A2(new_n409), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G224), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n462), .A2(G953), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n463), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n459), .A2(new_n465), .A3(new_n460), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT7), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n464), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  NOR3_X1   g283(.A1(new_n339), .A2(KEYINPUT5), .A3(G119), .ZN(new_n470));
  XNOR2_X1  g284(.A(G116), .B(G119), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n470), .B1(new_n471), .B2(KEYINPUT5), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G113), .ZN(new_n473));
  XOR2_X1   g287(.A(KEYINPUT2), .B(G113), .Z(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n471), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT83), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n243), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(G110), .B(G122), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n480), .B(KEYINPUT8), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n472), .A2(G113), .B1(new_n471), .B2(new_n474), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n482), .B1(KEYINPUT83), .B2(new_n281), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n479), .B(new_n481), .C1(new_n483), .C2(new_n478), .ZN(new_n484));
  INV_X1    g298(.A(new_n471), .ZN(new_n485));
  XNOR2_X1  g299(.A(KEYINPUT2), .B(G113), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(new_n475), .A3(KEYINPUT66), .ZN(new_n488));
  OR3_X1    g302(.A1(new_n474), .A2(KEYINPUT66), .A3(new_n471), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n257), .A2(new_n488), .A3(new_n255), .A4(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n482), .B1(new_n267), .B2(new_n268), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n491), .A3(new_n480), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n484), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n459), .A2(new_n467), .A3(new_n465), .A4(new_n460), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n469), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n490), .A2(new_n491), .ZN(new_n496));
  INV_X1    g310(.A(new_n480), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(KEYINPUT6), .A3(new_n492), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n459), .A2(new_n465), .A3(new_n460), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n465), .B1(new_n459), .B2(new_n460), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT6), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n496), .A2(new_n503), .A3(new_n497), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n499), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n495), .A2(new_n505), .A3(new_n189), .ZN(new_n506));
  OAI21_X1  g320(.A(G210), .B1(G237), .B2(G902), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n495), .A2(new_n505), .A3(new_n189), .A4(new_n507), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n458), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n388), .A2(new_n448), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT74), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n245), .A2(G119), .ZN(new_n514));
  INV_X1    g328(.A(G119), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(G128), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT24), .B(G110), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT71), .ZN(new_n520));
  OR2_X1    g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT23), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n522), .B1(new_n515), .B2(G128), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n245), .A2(KEYINPUT23), .A3(G119), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n516), .A3(new_n524), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n519), .A2(new_n520), .B1(G110), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n421), .A2(new_n521), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(G110), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n523), .A2(new_n524), .A3(new_n528), .A4(new_n516), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT73), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n517), .A2(new_n518), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n529), .A2(new_n530), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n396), .A2(new_n216), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n535), .A3(new_n413), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n527), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT22), .B(G137), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n193), .A2(G221), .A3(G234), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n538), .B(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n527), .A2(new_n536), .A3(new_n540), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n513), .B(KEYINPUT25), .C1(new_n544), .C2(new_n301), .ZN(new_n545));
  INV_X1    g359(.A(new_n543), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n540), .B1(new_n527), .B2(new_n536), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT25), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n549), .A2(KEYINPUT74), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(KEYINPUT74), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n548), .A2(new_n302), .A3(new_n551), .A4(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(G217), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n554), .B1(new_n302), .B2(G234), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n545), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n555), .A2(G902), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n548), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NOR3_X1   g373(.A1(new_n202), .A2(new_n203), .A3(G134), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n337), .A2(G137), .ZN(new_n561));
  OAI21_X1  g375(.A(G131), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n562), .A2(new_n206), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n252), .A2(new_n273), .B1(new_n563), .B2(new_n265), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n488), .A2(new_n489), .ZN(new_n565));
  AOI21_X1  g379(.A(KEYINPUT28), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n565), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n265), .A2(new_n206), .A3(new_n562), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n211), .A2(new_n206), .B1(new_n248), .B2(new_n251), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n273), .A2(new_n252), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n265), .A2(new_n206), .A3(new_n562), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(new_n565), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n566), .B1(KEYINPUT28), .B2(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(KEYINPUT26), .B(G101), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n392), .A2(G210), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT29), .B1(new_n575), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT69), .ZN(new_n582));
  INV_X1    g396(.A(new_n573), .ZN(new_n583));
  OAI21_X1  g397(.A(KEYINPUT30), .B1(new_n568), .B2(new_n569), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT30), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n571), .A2(new_n585), .A3(new_n572), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n583), .B1(new_n587), .B2(new_n567), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n582), .B1(new_n588), .B2(new_n580), .ZN(new_n589));
  INV_X1    g403(.A(new_n580), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n565), .B1(new_n584), .B2(new_n586), .ZN(new_n591));
  OAI211_X1 g405(.A(KEYINPUT69), .B(new_n590), .C1(new_n591), .C2(new_n583), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n581), .A2(new_n589), .A3(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n575), .A2(KEYINPUT29), .A3(new_n580), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(new_n302), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n586), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n585), .B1(new_n571), .B2(new_n572), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n567), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n573), .A2(new_n580), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(KEYINPUT68), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT68), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n573), .A2(new_n601), .A3(new_n580), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n598), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT31), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n574), .A2(KEYINPUT28), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n590), .B1(new_n605), .B2(new_n566), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT31), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n598), .A2(new_n600), .A3(new_n607), .A4(new_n602), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n604), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(G472), .A2(G902), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT32), .ZN(new_n612));
  AOI22_X1  g426(.A1(G472), .A2(new_n595), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n609), .A2(KEYINPUT32), .A3(new_n610), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n559), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n325), .A2(new_n512), .A3(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT94), .B(G101), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G3));
  INV_X1    g432(.A(new_n559), .ZN(new_n619));
  INV_X1    g433(.A(G472), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(new_n609), .B2(new_n302), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n610), .B2(new_n609), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n325), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n373), .A2(KEYINPUT33), .A3(new_n377), .ZN(new_n624));
  AOI21_X1  g438(.A(KEYINPUT33), .B1(new_n373), .B2(new_n377), .ZN(new_n625));
  OAI211_X1 g439(.A(G478), .B(new_n302), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(KEYINPUT95), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n379), .A2(new_n380), .A3(new_n383), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT33), .ZN(new_n629));
  INV_X1    g443(.A(new_n377), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n371), .B1(new_n376), .B2(new_n351), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n373), .A2(KEYINPUT33), .A3(new_n377), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT95), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n634), .A2(new_n635), .A3(G478), .A4(new_n302), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n627), .A2(new_n628), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n434), .A2(new_n444), .A3(new_n447), .ZN(new_n638));
  INV_X1    g452(.A(new_n456), .ZN(new_n639));
  INV_X1    g453(.A(new_n455), .ZN(new_n640));
  AOI211_X1 g454(.A(new_n639), .B(new_n640), .C1(new_n509), .C2(new_n510), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n637), .A2(new_n638), .A3(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n623), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT34), .B(G104), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  OAI21_X1  g460(.A(new_n441), .B1(new_n445), .B2(new_n446), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n443), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n648), .A2(new_n434), .A3(new_n447), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n641), .A2(new_n387), .A3(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n623), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT35), .B(G107), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  NOR2_X1   g468(.A1(new_n541), .A2(KEYINPUT36), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n537), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n557), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n556), .A2(KEYINPUT96), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(KEYINPUT96), .B1(new_n556), .B2(new_n657), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n325), .A2(new_n512), .A3(new_n622), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G110), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT97), .B(KEYINPUT37), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G12));
  AOI21_X1  g479(.A(new_n660), .B1(new_n613), .B2(new_n614), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n452), .B1(new_n453), .B2(G900), .ZN(new_n667));
  AND4_X1   g481(.A1(new_n447), .A2(new_n648), .A3(new_n434), .A4(new_n667), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n668), .A2(new_n387), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n639), .B1(new_n509), .B2(new_n510), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n325), .A2(new_n666), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G128), .ZN(G30));
  NAND2_X1  g487(.A1(new_n556), .A2(new_n657), .ZN(new_n674));
  INV_X1    g488(.A(new_n574), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n603), .B1(new_n675), .B2(new_n580), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n620), .B1(new_n676), .B2(new_n189), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n677), .B1(new_n611), .B2(new_n612), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n674), .B1(new_n678), .B2(new_n614), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n509), .A2(new_n510), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT38), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n387), .A2(new_n638), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n682), .A2(new_n639), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n667), .B(KEYINPUT39), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n325), .A2(KEYINPUT40), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(KEYINPUT40), .B1(new_n325), .B2(new_n685), .ZN(new_n687));
  OAI211_X1 g501(.A(new_n679), .B(new_n684), .C1(new_n686), .C2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G143), .ZN(G45));
  AND3_X1   g503(.A1(new_n637), .A2(new_n638), .A3(new_n667), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n325), .A2(new_n670), .A3(new_n666), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G146), .ZN(G48));
  NAND2_X1  g506(.A1(new_n595), .A2(G472), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n611), .A2(new_n612), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n693), .A2(new_n694), .A3(new_n614), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n311), .A2(new_n312), .ZN(new_n696));
  OAI21_X1  g510(.A(G469), .B1(new_n696), .B2(new_n301), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n697), .A2(new_n191), .A3(new_n313), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n642), .A2(new_n619), .A3(new_n695), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT41), .B(G113), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G15));
  NAND4_X1  g515(.A1(new_n650), .A2(new_n698), .A3(new_n695), .A4(new_n619), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G116), .ZN(G18));
  AND4_X1   g517(.A1(new_n191), .A2(new_n697), .A3(new_n313), .A4(new_n670), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n387), .A2(new_n638), .A3(new_n640), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n704), .A2(new_n695), .A3(new_n661), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G119), .ZN(G21));
  XNOR2_X1  g521(.A(new_n610), .B(KEYINPUT98), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n609), .A2(new_n708), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n709), .A2(new_n621), .A3(new_n559), .ZN(new_n710));
  INV_X1    g524(.A(new_n670), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n683), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n710), .A2(new_n698), .A3(new_n712), .A4(new_n455), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT99), .B(G122), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G24));
  INV_X1    g529(.A(new_n674), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n709), .A2(new_n621), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n690), .A2(new_n704), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G125), .ZN(G27));
  INV_X1    g533(.A(KEYINPUT100), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n294), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n292), .A2(KEYINPUT100), .A3(new_n293), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n721), .A2(G469), .A3(new_n276), .A4(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n313), .A2(new_n723), .A3(new_n315), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT101), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n313), .A2(new_n723), .A3(KEYINPUT101), .A4(new_n315), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n509), .A2(new_n510), .A3(new_n456), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT102), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT102), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n509), .A2(new_n731), .A3(new_n510), .A4(new_n456), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n730), .A2(new_n191), .A3(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n615), .A2(new_n690), .A3(new_n728), .A4(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT42), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT103), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n614), .B(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n559), .B1(new_n739), .B2(new_n613), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n733), .B1(new_n726), .B2(new_n727), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n740), .A2(KEYINPUT42), .A3(new_n690), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n737), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G131), .ZN(G33));
  AND3_X1   g558(.A1(new_n741), .A2(new_n615), .A3(new_n669), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n337), .ZN(G36));
  NAND2_X1  g560(.A1(new_n637), .A2(new_n448), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT43), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(KEYINPUT43), .B1(new_n637), .B2(new_n448), .ZN(new_n750));
  OR2_X1    g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n622), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n751), .A2(KEYINPUT44), .A3(new_n752), .A4(new_n674), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n752), .B(new_n674), .C1(new_n749), .C2(new_n750), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT44), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n730), .A2(new_n732), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n753), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT105), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n321), .A2(new_n296), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n299), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n721), .A2(KEYINPUT45), .A3(new_n276), .A4(new_n722), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n314), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OR3_X1    g578(.A1(new_n764), .A2(KEYINPUT104), .A3(KEYINPUT46), .ZN(new_n765));
  OAI21_X1  g579(.A(KEYINPUT104), .B1(new_n764), .B2(KEYINPUT46), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n764), .A2(KEYINPUT46), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n765), .A2(new_n766), .A3(new_n313), .A4(new_n767), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n768), .A2(new_n191), .A3(new_n685), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT105), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n753), .A2(new_n756), .A3(new_n770), .A4(new_n757), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n759), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G137), .ZN(G39));
  INV_X1    g587(.A(new_n695), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n637), .A2(new_n638), .ZN(new_n775));
  INV_X1    g589(.A(new_n667), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n775), .A2(new_n619), .A3(new_n776), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n768), .A2(KEYINPUT47), .A3(new_n191), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT47), .B1(new_n768), .B2(new_n191), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n774), .B(new_n777), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n757), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G140), .ZN(G42));
  NOR2_X1   g597(.A1(new_n778), .A2(new_n779), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n697), .A2(new_n313), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n190), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(KEYINPUT112), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n751), .A2(new_n451), .A3(new_n450), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(new_n710), .A3(new_n757), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT112), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n784), .A2(new_n792), .A3(new_n786), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n788), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n785), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(new_n733), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n678), .A2(new_n614), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n452), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n796), .A2(new_n619), .A3(new_n798), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n799), .A2(new_n638), .A3(new_n637), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n789), .A2(new_n796), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n800), .B1(new_n802), .B2(new_n717), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n794), .A2(KEYINPUT51), .A3(new_n803), .ZN(new_n804));
  OR2_X1    g618(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n698), .A2(KEYINPUT110), .A3(new_n639), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT110), .B1(new_n698), .B2(new_n639), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n807), .A2(new_n681), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n789), .A2(new_n710), .A3(new_n806), .A4(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT50), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  AOI22_X1  g626(.A1(new_n804), .A2(new_n805), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n787), .A2(new_n791), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n812), .A2(KEYINPUT111), .A3(new_n811), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(new_n815), .A3(new_n803), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT51), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n683), .A2(new_n711), .A3(new_n776), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n679), .A2(new_n728), .A3(new_n820), .A4(new_n191), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n691), .A2(new_n672), .A3(new_n718), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT52), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n690), .A2(new_n704), .A3(new_n717), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n661), .A2(new_n695), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n825), .B1(new_n319), .B2(new_n324), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n824), .B1(new_n826), .B2(new_n671), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n827), .A2(new_n828), .A3(new_n691), .A4(new_n821), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n823), .A2(new_n829), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n730), .A2(new_n668), .A3(new_n732), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n270), .B1(new_n274), .B2(new_n275), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(new_n293), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n292), .A2(new_n293), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n301), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n314), .B1(new_n835), .B2(new_n299), .ZN(new_n836));
  AOI211_X1 g650(.A(new_n318), .B(new_n190), .C1(new_n836), .C2(new_n322), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT81), .B1(new_n323), .B2(new_n191), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n666), .B(new_n831), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n387), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n699), .A2(new_n702), .A3(new_n706), .A4(new_n713), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n745), .B1(new_n737), .B2(new_n742), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n690), .A2(new_n728), .A3(new_n734), .A4(new_n717), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT109), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT109), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n741), .A2(new_n847), .A3(new_n690), .A4(new_n717), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n637), .A2(new_n638), .A3(new_n511), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n387), .A2(new_n448), .A3(new_n511), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT108), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT108), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n387), .A2(new_n448), .A3(new_n511), .A4(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n850), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n325), .A2(new_n619), .A3(new_n622), .A4(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n849), .A2(new_n616), .A3(new_n662), .A4(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n844), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT53), .B1(new_n830), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n823), .A2(new_n829), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n662), .A2(new_n856), .A3(new_n616), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(new_n842), .A3(new_n843), .A4(new_n849), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n860), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n819), .B1(new_n859), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n830), .A2(new_n858), .A3(KEYINPUT53), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n863), .B1(new_n860), .B2(new_n862), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n866), .A2(new_n867), .A3(KEYINPUT54), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n740), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT114), .ZN(new_n871));
  OAI22_X1  g685(.A1(new_n801), .A2(new_n870), .B1(new_n871), .B2(KEYINPUT48), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(KEYINPUT48), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n871), .A2(KEYINPUT48), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n789), .A2(new_n740), .A3(new_n796), .A4(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n450), .A2(KEYINPUT113), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n789), .A2(new_n704), .A3(new_n710), .ZN(new_n878));
  OAI22_X1  g692(.A1(new_n799), .A2(new_n775), .B1(KEYINPUT113), .B2(new_n450), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n876), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n881), .A2(KEYINPUT115), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n881), .A2(KEYINPUT115), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n818), .B(new_n869), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  OAI22_X1  g698(.A1(new_n813), .A2(new_n884), .B1(G952), .B2(G953), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n619), .A2(new_n457), .A3(new_n191), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(KEYINPUT106), .Z(new_n887));
  AOI21_X1  g701(.A(new_n747), .B1(new_n795), .B2(KEYINPUT49), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n887), .A2(KEYINPUT107), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n682), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT107), .B1(new_n887), .B2(new_n888), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n795), .A2(KEYINPUT49), .ZN(new_n892));
  OR4_X1    g706(.A1(new_n797), .A2(new_n890), .A3(new_n891), .A4(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n885), .A2(new_n893), .ZN(G75));
  NAND2_X1  g708(.A1(new_n449), .A2(G953), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT118), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT56), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n866), .A2(new_n867), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n301), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n898), .B1(new_n900), .B2(new_n507), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n499), .A2(new_n504), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(new_n502), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT116), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT55), .Z(new_n905));
  AOI21_X1  g719(.A(new_n905), .B1(KEYINPUT117), .B2(new_n898), .ZN(new_n906));
  OR2_X1    g720(.A1(new_n901), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n901), .A2(new_n906), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n897), .B1(new_n907), .B2(new_n908), .ZN(G51));
  XNOR2_X1  g723(.A(new_n314), .B(KEYINPUT57), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n865), .A2(new_n868), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n696), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n911), .A2(KEYINPUT119), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(KEYINPUT119), .B1(new_n911), .B2(new_n912), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n900), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n916), .A2(new_n763), .A3(new_n762), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n897), .B1(new_n915), .B2(new_n917), .ZN(G54));
  NAND2_X1  g732(.A1(KEYINPUT58), .A2(G475), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(KEYINPUT120), .ZN(new_n920));
  OR2_X1    g734(.A1(new_n919), .A2(KEYINPUT120), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n916), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n445), .A2(new_n446), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n922), .A2(new_n923), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n924), .A2(new_n925), .A3(new_n897), .ZN(G60));
  NAND2_X1  g740(.A1(G478), .A2(G902), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT59), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n865), .A2(new_n634), .A3(new_n868), .A4(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT121), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n929), .A2(new_n930), .A3(new_n896), .ZN(new_n931));
  INV_X1    g745(.A(new_n869), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n634), .B1(new_n932), .B2(new_n928), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n930), .B1(new_n929), .B2(new_n896), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n931), .A2(new_n933), .A3(new_n934), .ZN(G63));
  NAND2_X1  g749(.A1(G217), .A2(G902), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT60), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(new_n866), .B2(new_n867), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n656), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n939), .B(new_n896), .C1(new_n548), .C2(new_n938), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT61), .B1(new_n939), .B2(KEYINPUT122), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(G66));
  AOI21_X1  g756(.A(new_n193), .B1(new_n454), .B2(G224), .ZN(new_n943));
  INV_X1    g757(.A(new_n861), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n944), .A2(new_n841), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n943), .B1(new_n946), .B2(new_n193), .ZN(new_n947));
  INV_X1    g761(.A(G898), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n902), .B1(new_n948), .B2(G953), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n947), .B(new_n949), .ZN(G69));
  NAND2_X1  g764(.A1(G900), .A2(G953), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n587), .B(new_n435), .Z(new_n952));
  INV_X1    g766(.A(new_n843), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n769), .A2(new_n740), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n953), .B1(new_n954), .B2(new_n712), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n827), .A2(new_n691), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n772), .A2(KEYINPUT125), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(KEYINPUT125), .B1(new_n772), .B2(new_n956), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n782), .B(new_n955), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n951), .B(new_n952), .C1(new_n959), .C2(G953), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n775), .B1(new_n638), .B2(new_n388), .ZN(new_n961));
  AOI211_X1 g775(.A(new_n559), .B(new_n774), .C1(new_n961), .C2(KEYINPUT124), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n961), .A2(KEYINPUT124), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n962), .A2(new_n325), .A3(new_n685), .A4(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n781), .B1(new_n780), .B2(new_n964), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n956), .A2(KEYINPUT62), .A3(new_n688), .ZN(new_n966));
  AOI21_X1  g780(.A(KEYINPUT62), .B1(new_n956), .B2(new_n688), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n772), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n193), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n952), .B(KEYINPUT123), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n960), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n193), .B1(G227), .B2(G900), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n973), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n960), .A2(new_n971), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n974), .A2(new_n976), .ZN(G72));
  NAND2_X1  g791(.A1(G472), .A2(G902), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT63), .Z(new_n979));
  OAI21_X1  g793(.A(new_n979), .B1(new_n959), .B2(new_n946), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n588), .A2(new_n590), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT127), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n897), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n965), .ZN(new_n984));
  OR2_X1    g798(.A1(new_n966), .A2(new_n967), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n984), .A2(new_n985), .A3(new_n772), .A4(new_n945), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT126), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n986), .A2(new_n987), .A3(new_n979), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n965), .A2(new_n968), .A3(new_n946), .ZN(new_n989));
  INV_X1    g803(.A(new_n979), .ZN(new_n990));
  OAI21_X1  g804(.A(KEYINPUT126), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n588), .A2(new_n590), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n988), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n589), .A2(new_n603), .A3(new_n592), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n899), .A2(new_n979), .A3(new_n994), .ZN(new_n995));
  AND3_X1   g809(.A1(new_n983), .A2(new_n993), .A3(new_n995), .ZN(G57));
endmodule


