

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753;

  XNOR2_X1 U379 ( .A(n382), .B(n472), .ZN(n531) );
  AND2_X1 U380 ( .A1(n572), .A2(n471), .ZN(n382) );
  XNOR2_X1 U381 ( .A(n452), .B(G119), .ZN(n454) );
  XNOR2_X1 U382 ( .A(G113), .B(G101), .ZN(n453) );
  NOR2_X1 U383 ( .A1(n528), .A2(n583), .ZN(n368) );
  XNOR2_X1 U384 ( .A(n422), .B(n421), .ZN(n511) );
  AND2_X1 U385 ( .A1(n511), .A2(n504), .ZN(n639) );
  AND2_X1 U386 ( .A1(n572), .A2(n571), .ZN(n355) );
  NOR2_X2 U387 ( .A1(n605), .A2(n611), .ZN(n548) );
  OR2_X2 U388 ( .A1(n625), .A2(G902), .ZN(n501) );
  NOR2_X2 U389 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X2 U390 ( .A(n444), .B(KEYINPUT73), .ZN(n476) );
  XNOR2_X2 U391 ( .A(n366), .B(n514), .ZN(n622) );
  XNOR2_X1 U392 ( .A(n551), .B(n363), .ZN(n696) );
  INV_X1 U393 ( .A(n594), .ZN(n583) );
  INV_X1 U394 ( .A(n558), .ZN(n677) );
  OR2_X1 U395 ( .A1(n609), .A2(n730), .ZN(n660) );
  XNOR2_X1 U396 ( .A(n358), .B(n357), .ZN(n750) );
  NAND2_X1 U397 ( .A1(n696), .A2(n571), .ZN(n358) );
  NOR2_X1 U398 ( .A1(n715), .A2(n725), .ZN(n716) );
  AND2_X1 U399 ( .A1(n742), .A2(n605), .ZN(n403) );
  AND2_X1 U400 ( .A1(n370), .A2(n602), .ZN(n742) );
  OR2_X1 U401 ( .A1(n750), .A2(n753), .ZN(n383) );
  OR2_X1 U402 ( .A1(n666), .A2(n665), .ZN(n551) );
  XNOR2_X1 U403 ( .A(n388), .B(n387), .ZN(n674) );
  XNOR2_X1 U404 ( .A(n400), .B(G146), .ZN(n448) );
  XNOR2_X1 U405 ( .A(n559), .B(KEYINPUT106), .ZN(n357) );
  INV_X1 U406 ( .A(KEYINPUT3), .ZN(n452) );
  XNOR2_X1 U407 ( .A(G143), .B(G128), .ZN(n460) );
  XNOR2_X1 U408 ( .A(KEYINPUT71), .B(G131), .ZN(n485) );
  XNOR2_X2 U409 ( .A(n356), .B(KEYINPUT16), .ZN(n458) );
  XNOR2_X1 U410 ( .A(n356), .B(n493), .ZN(n496) );
  XNOR2_X2 U411 ( .A(n454), .B(n453), .ZN(n356) );
  XNOR2_X2 U412 ( .A(n458), .B(n457), .ZN(n726) );
  XNOR2_X1 U413 ( .A(n369), .B(G104), .ZN(n455) );
  INV_X1 U414 ( .A(G122), .ZN(n369) );
  OR2_X1 U415 ( .A1(n575), .A2(n376), .ZN(n375) );
  NAND2_X1 U416 ( .A1(n355), .A2(KEYINPUT81), .ZN(n374) );
  NAND2_X1 U417 ( .A1(n392), .A2(n360), .ZN(n577) );
  NAND2_X1 U418 ( .A1(n393), .A2(KEYINPUT47), .ZN(n392) );
  XNOR2_X1 U419 ( .A(n389), .B(KEYINPUT20), .ZN(n443) );
  NAND2_X1 U420 ( .A1(n418), .A2(G234), .ZN(n389) );
  XNOR2_X1 U421 ( .A(n448), .B(n399), .ZN(n428) );
  INV_X1 U422 ( .A(KEYINPUT10), .ZN(n399) );
  XNOR2_X1 U423 ( .A(n487), .B(n486), .ZN(n741) );
  XNOR2_X1 U424 ( .A(n726), .B(n461), .ZN(n462) );
  XNOR2_X1 U425 ( .A(n593), .B(n592), .ZN(n370) );
  NAND2_X1 U426 ( .A1(n580), .A2(n397), .ZN(n396) );
  NOR2_X1 U427 ( .A1(n558), .A2(n398), .ZN(n397) );
  INV_X1 U428 ( .A(n674), .ZN(n398) );
  INV_X1 U429 ( .A(KEYINPUT28), .ZN(n395) );
  INV_X1 U430 ( .A(KEYINPUT38), .ZN(n549) );
  NOR2_X1 U431 ( .A1(n557), .A2(n560), .ZN(n580) );
  XNOR2_X1 U432 ( .A(n371), .B(n361), .ZN(n534) );
  OR2_X1 U433 ( .A1(n712), .A2(G902), .ZN(n371) );
  INV_X1 U434 ( .A(n511), .ZN(n557) );
  XNOR2_X1 U435 ( .A(n475), .B(n474), .ZN(n507) );
  XNOR2_X1 U436 ( .A(n473), .B(KEYINPUT67), .ZN(n474) );
  NAND2_X1 U437 ( .A1(n381), .A2(n379), .ZN(n475) );
  INV_X1 U438 ( .A(KEYINPUT22), .ZN(n473) );
  XNOR2_X1 U439 ( .A(n545), .B(n544), .ZN(n730) );
  XOR2_X1 U440 ( .A(KEYINPUT11), .B(G140), .Z(n430) );
  XNOR2_X1 U441 ( .A(G113), .B(G143), .ZN(n429) );
  XNOR2_X1 U442 ( .A(n455), .B(n485), .ZN(n426) );
  INV_X1 U443 ( .A(KEYINPUT12), .ZN(n373) );
  XNOR2_X1 U444 ( .A(n741), .B(G146), .ZN(n498) );
  XNOR2_X1 U445 ( .A(G101), .B(G104), .ZN(n479) );
  INV_X1 U446 ( .A(G107), .ZN(n481) );
  XNOR2_X1 U447 ( .A(n368), .B(KEYINPUT33), .ZN(n698) );
  OR2_X1 U448 ( .A1(n531), .A2(n698), .ZN(n513) );
  OR2_X1 U449 ( .A1(n573), .A2(n667), .ZN(n393) );
  INV_X1 U450 ( .A(G125), .ZN(n400) );
  XNOR2_X1 U451 ( .A(n460), .B(n459), .ZN(n487) );
  XNOR2_X1 U452 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n459) );
  INV_X1 U453 ( .A(n487), .ZN(n461) );
  NOR2_X1 U454 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U455 ( .A1(n375), .A2(n374), .ZN(n576) );
  INV_X1 U456 ( .A(KEYINPUT46), .ZN(n570) );
  XNOR2_X1 U457 ( .A(n417), .B(G902), .ZN(n605) );
  INV_X1 U458 ( .A(KEYINPUT15), .ZN(n417) );
  AND2_X1 U459 ( .A1(n550), .A2(n380), .ZN(n379) );
  INV_X1 U460 ( .A(n510), .ZN(n380) );
  XNOR2_X1 U461 ( .A(G137), .B(G116), .ZN(n492) );
  XOR2_X1 U462 ( .A(G137), .B(G140), .Z(n477) );
  INV_X1 U463 ( .A(KEYINPUT21), .ZN(n387) );
  NAND2_X1 U464 ( .A1(n443), .A2(G221), .ZN(n388) );
  XOR2_X1 U465 ( .A(KEYINPUT8), .B(KEYINPUT70), .Z(n406) );
  XNOR2_X1 U466 ( .A(n405), .B(n404), .ZN(n407) );
  INV_X1 U467 ( .A(KEYINPUT83), .ZN(n404) );
  XNOR2_X1 U468 ( .A(G128), .B(KEYINPUT24), .ZN(n408) );
  INV_X1 U469 ( .A(KEYINPUT79), .ZN(n410) );
  XNOR2_X1 U470 ( .A(G119), .B(G110), .ZN(n411) );
  XOR2_X1 U471 ( .A(G116), .B(G107), .Z(n456) );
  XOR2_X1 U472 ( .A(G134), .B(G122), .Z(n435) );
  XNOR2_X1 U473 ( .A(n384), .B(KEYINPUT86), .ZN(n609) );
  AND2_X1 U474 ( .A1(n394), .A2(n552), .ZN(n571) );
  XNOR2_X1 U475 ( .A(n396), .B(n395), .ZN(n394) );
  XNOR2_X1 U476 ( .A(n568), .B(n567), .ZN(n600) );
  INV_X1 U477 ( .A(KEYINPUT39), .ZN(n567) );
  AND2_X1 U478 ( .A1(n565), .A2(n385), .ZN(n568) );
  XNOR2_X1 U479 ( .A(n377), .B(n509), .ZN(n520) );
  NAND2_X1 U480 ( .A1(n508), .A2(n583), .ZN(n378) );
  NOR2_X1 U481 ( .A1(G902), .A2(n721), .ZN(n422) );
  INV_X1 U482 ( .A(KEYINPUT25), .ZN(n419) );
  XNOR2_X1 U483 ( .A(n432), .B(n372), .ZN(n712) );
  XNOR2_X1 U484 ( .A(n431), .B(n401), .ZN(n432) );
  XNOR2_X1 U485 ( .A(n427), .B(n373), .ZN(n372) );
  BUF_X1 U486 ( .A(n711), .Z(n720) );
  XNOR2_X1 U487 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U488 ( .A(n480), .B(n479), .ZN(n484) );
  XNOR2_X1 U489 ( .A(n569), .B(KEYINPUT40), .ZN(n753) );
  AND2_X1 U490 ( .A1(n644), .A2(n600), .ZN(n569) );
  NAND2_X1 U491 ( .A1(n367), .A2(n359), .ZN(n366) );
  XNOR2_X1 U492 ( .A(n513), .B(n512), .ZN(n367) );
  NAND2_X1 U493 ( .A1(n359), .A2(n391), .ZN(n390) );
  AND2_X1 U494 ( .A1(n534), .A2(n535), .ZN(n359) );
  NOR2_X1 U495 ( .A1(n643), .A2(n365), .ZN(n360) );
  XNOR2_X1 U496 ( .A(n558), .B(KEYINPUT6), .ZN(n594) );
  XOR2_X1 U497 ( .A(n434), .B(n433), .Z(n361) );
  INV_X1 U498 ( .A(n531), .ZN(n381) );
  XNOR2_X1 U499 ( .A(n548), .B(n547), .ZN(n598) );
  AND2_X1 U500 ( .A1(n602), .A2(KEYINPUT2), .ZN(n362) );
  XOR2_X1 U501 ( .A(KEYINPUT105), .B(KEYINPUT41), .Z(n363) );
  XNOR2_X1 U502 ( .A(KEYINPUT47), .B(KEYINPUT69), .ZN(n364) );
  AND2_X1 U503 ( .A1(KEYINPUT81), .A2(n574), .ZN(n365) );
  XNOR2_X1 U504 ( .A(n622), .B(KEYINPUT68), .ZN(n515) );
  NAND2_X1 U505 ( .A1(n370), .A2(n362), .ZN(n384) );
  NAND2_X1 U506 ( .A1(n355), .A2(n364), .ZN(n376) );
  XNOR2_X1 U507 ( .A(n667), .B(KEYINPUT82), .ZN(n575) );
  NOR2_X1 U508 ( .A1(n507), .A2(n378), .ZN(n377) );
  XNOR2_X1 U509 ( .A(n383), .B(n570), .ZN(n591) );
  XNOR2_X2 U510 ( .A(n552), .B(KEYINPUT1), .ZN(n680) );
  NOR2_X1 U511 ( .A1(n639), .A2(n752), .ZN(n516) );
  NAND2_X1 U512 ( .A1(n565), .A2(n564), .ZN(n386) );
  AND2_X1 U513 ( .A1(n564), .A2(n663), .ZN(n385) );
  NOR2_X1 U514 ( .A1(n386), .A2(n390), .ZN(n643) );
  INV_X1 U515 ( .A(n598), .ZN(n391) );
  XNOR2_X2 U516 ( .A(G110), .B(KEYINPUT74), .ZN(n444) );
  NOR2_X2 U517 ( .A1(n511), .A2(n510), .ZN(n681) );
  XNOR2_X2 U518 ( .A(n490), .B(G469), .ZN(n552) );
  XNOR2_X2 U519 ( .A(n501), .B(n500), .ZN(n558) );
  XOR2_X1 U520 ( .A(n430), .B(n429), .Z(n401) );
  OR2_X1 U521 ( .A1(G902), .A2(n717), .ZN(n402) );
  INV_X1 U522 ( .A(KEYINPUT76), .ZN(n578) );
  INV_X1 U523 ( .A(KEYINPUT80), .ZN(n445) );
  INV_X1 U524 ( .A(n652), .ZN(n588) );
  XNOR2_X1 U525 ( .A(n446), .B(n445), .ZN(n447) );
  NOR2_X1 U526 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U527 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U528 ( .A(n407), .B(n406), .ZN(n438) );
  XNOR2_X1 U529 ( .A(n484), .B(n483), .ZN(n488) );
  INV_X1 U530 ( .A(KEYINPUT42), .ZN(n559) );
  INV_X1 U531 ( .A(n546), .ZN(n547) );
  XNOR2_X1 U532 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U533 ( .A(n618), .B(KEYINPUT56), .ZN(n619) );
  INV_X2 U534 ( .A(G953), .ZN(n743) );
  NAND2_X1 U535 ( .A1(G234), .A2(n743), .ZN(n405) );
  AND2_X1 U536 ( .A1(n438), .A2(G221), .ZN(n415) );
  XOR2_X1 U537 ( .A(KEYINPUT23), .B(KEYINPUT92), .Z(n409) );
  XNOR2_X1 U538 ( .A(n409), .B(n408), .ZN(n413) );
  XNOR2_X1 U539 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U540 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U541 ( .A(n428), .B(n477), .Z(n740) );
  XNOR2_X1 U542 ( .A(n416), .B(n740), .ZN(n721) );
  INV_X1 U543 ( .A(n605), .ZN(n418) );
  NAND2_X1 U544 ( .A1(n443), .A2(G217), .ZN(n420) );
  NOR2_X1 U545 ( .A1(G953), .A2(G237), .ZN(n424) );
  INV_X1 U546 ( .A(KEYINPUT77), .ZN(n423) );
  XNOR2_X1 U547 ( .A(n424), .B(n423), .ZN(n494) );
  NAND2_X1 U548 ( .A1(G214), .A2(n494), .ZN(n425) );
  XNOR2_X1 U549 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U550 ( .A(n428), .B(KEYINPUT98), .ZN(n431) );
  XNOR2_X1 U551 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n434) );
  INV_X1 U552 ( .A(G475), .ZN(n433) );
  XNOR2_X1 U553 ( .A(n456), .B(KEYINPUT7), .ZN(n437) );
  XNOR2_X1 U554 ( .A(n460), .B(n435), .ZN(n436) );
  XNOR2_X1 U555 ( .A(n437), .B(n436), .ZN(n442) );
  XOR2_X1 U556 ( .A(KEYINPUT9), .B(KEYINPUT101), .Z(n440) );
  NAND2_X1 U557 ( .A1(G217), .A2(n438), .ZN(n439) );
  XNOR2_X1 U558 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U559 ( .A(n442), .B(n441), .ZN(n717) );
  XNOR2_X1 U560 ( .A(G478), .B(n402), .ZN(n535) );
  NOR2_X1 U561 ( .A1(n534), .A2(n535), .ZN(n550) );
  XNOR2_X1 U562 ( .A(KEYINPUT93), .B(n674), .ZN(n510) );
  NAND2_X1 U563 ( .A1(G224), .A2(n743), .ZN(n446) );
  XNOR2_X1 U564 ( .A(n476), .B(n447), .ZN(n451) );
  XNOR2_X1 U565 ( .A(n448), .B(KEYINPUT18), .ZN(n449) );
  XNOR2_X1 U566 ( .A(n449), .B(KEYINPUT17), .ZN(n450) );
  XOR2_X1 U567 ( .A(n451), .B(n450), .Z(n463) );
  XOR2_X1 U568 ( .A(n456), .B(n455), .Z(n457) );
  XNOR2_X1 U569 ( .A(n463), .B(n462), .ZN(n611) );
  OR2_X1 U570 ( .A1(G237), .A2(G902), .ZN(n464) );
  NAND2_X1 U571 ( .A1(G210), .A2(n464), .ZN(n546) );
  XNOR2_X1 U572 ( .A(n548), .B(n546), .ZN(n465) );
  NAND2_X1 U573 ( .A1(G214), .A2(n464), .ZN(n662) );
  NAND2_X1 U574 ( .A1(n465), .A2(n662), .ZN(n466) );
  XNOR2_X1 U575 ( .A(n466), .B(KEYINPUT19), .ZN(n572) );
  NAND2_X1 U576 ( .A1(G234), .A2(G237), .ZN(n467) );
  XNOR2_X1 U577 ( .A(n467), .B(KEYINPUT14), .ZN(n468) );
  NAND2_X1 U578 ( .A1(G952), .A2(n468), .ZN(n695) );
  NOR2_X1 U579 ( .A1(G953), .A2(n695), .ZN(n556) );
  NAND2_X1 U580 ( .A1(G902), .A2(n468), .ZN(n553) );
  INV_X1 U581 ( .A(G898), .ZN(n735) );
  NAND2_X1 U582 ( .A1(G953), .A2(n735), .ZN(n728) );
  NOR2_X1 U583 ( .A1(n553), .A2(n728), .ZN(n469) );
  NOR2_X1 U584 ( .A1(n556), .A2(n469), .ZN(n470) );
  XNOR2_X1 U585 ( .A(KEYINPUT91), .B(n470), .ZN(n471) );
  INV_X1 U586 ( .A(KEYINPUT0), .ZN(n472) );
  XNOR2_X1 U587 ( .A(n477), .B(n476), .ZN(n478) );
  INV_X1 U588 ( .A(n478), .ZN(n480) );
  NAND2_X1 U589 ( .A1(G227), .A2(n743), .ZN(n482) );
  XNOR2_X1 U590 ( .A(n485), .B(G134), .ZN(n486) );
  XNOR2_X1 U591 ( .A(n488), .B(n498), .ZN(n707) );
  INV_X1 U592 ( .A(G902), .ZN(n489) );
  NAND2_X1 U593 ( .A1(n707), .A2(n489), .ZN(n490) );
  NOR2_X1 U594 ( .A1(n507), .A2(n680), .ZN(n525) );
  XNOR2_X1 U595 ( .A(KEYINPUT95), .B(KEYINPUT5), .ZN(n491) );
  XNOR2_X1 U596 ( .A(n492), .B(n491), .ZN(n493) );
  NAND2_X1 U597 ( .A1(n494), .A2(G210), .ZN(n495) );
  XNOR2_X1 U598 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U599 ( .A(n498), .B(n497), .ZN(n625) );
  XNOR2_X1 U600 ( .A(G472), .B(KEYINPUT96), .ZN(n499) );
  XNOR2_X1 U601 ( .A(n499), .B(KEYINPUT75), .ZN(n500) );
  NAND2_X1 U602 ( .A1(n525), .A2(n558), .ZN(n503) );
  INV_X1 U603 ( .A(KEYINPUT66), .ZN(n502) );
  XNOR2_X1 U604 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U605 ( .A(KEYINPUT102), .B(n557), .ZN(n675) );
  XNOR2_X1 U606 ( .A(n680), .B(KEYINPUT90), .ZN(n586) );
  INV_X1 U607 ( .A(n586), .ZN(n505) );
  NOR2_X1 U608 ( .A1(n675), .A2(n505), .ZN(n506) );
  XNOR2_X1 U609 ( .A(n506), .B(KEYINPUT104), .ZN(n508) );
  INV_X1 U610 ( .A(KEYINPUT32), .ZN(n509) );
  INV_X1 U611 ( .A(n520), .ZN(n752) );
  NAND2_X1 U612 ( .A1(n681), .A2(n680), .ZN(n528) );
  INV_X1 U613 ( .A(KEYINPUT34), .ZN(n512) );
  INV_X1 U614 ( .A(KEYINPUT35), .ZN(n514) );
  NAND2_X1 U615 ( .A1(n516), .A2(n515), .ZN(n518) );
  INV_X1 U616 ( .A(KEYINPUT44), .ZN(n517) );
  NAND2_X1 U617 ( .A1(n518), .A2(n517), .ZN(n524) );
  AND2_X1 U618 ( .A1(KEYINPUT44), .A2(KEYINPUT68), .ZN(n519) );
  NAND2_X1 U619 ( .A1(n520), .A2(n519), .ZN(n521) );
  NOR2_X1 U620 ( .A1(n639), .A2(n521), .ZN(n522) );
  NAND2_X1 U621 ( .A1(n522), .A2(n622), .ZN(n523) );
  NAND2_X1 U622 ( .A1(n524), .A2(n523), .ZN(n542) );
  NAND2_X1 U623 ( .A1(n525), .A2(n583), .ZN(n526) );
  XNOR2_X1 U624 ( .A(n526), .B(KEYINPUT87), .ZN(n527) );
  NAND2_X1 U625 ( .A1(n527), .A2(n675), .ZN(n631) );
  NOR2_X1 U626 ( .A1(n528), .A2(n558), .ZN(n529) );
  XNOR2_X1 U627 ( .A(n529), .B(KEYINPUT97), .ZN(n686) );
  NOR2_X1 U628 ( .A1(n686), .A2(n531), .ZN(n530) );
  XNOR2_X1 U629 ( .A(n530), .B(KEYINPUT31), .ZN(n649) );
  NAND2_X1 U630 ( .A1(n681), .A2(n552), .ZN(n532) );
  XNOR2_X1 U631 ( .A(n532), .B(KEYINPUT94), .ZN(n561) );
  NOR2_X1 U632 ( .A1(n561), .A2(n677), .ZN(n533) );
  NAND2_X1 U633 ( .A1(n381), .A2(n533), .ZN(n634) );
  NAND2_X1 U634 ( .A1(n649), .A2(n634), .ZN(n538) );
  XOR2_X1 U635 ( .A(n534), .B(KEYINPUT100), .Z(n536) );
  NOR2_X1 U636 ( .A1(n536), .A2(n535), .ZN(n644) );
  AND2_X1 U637 ( .A1(n536), .A2(n535), .ZN(n640) );
  NOR2_X1 U638 ( .A1(n644), .A2(n640), .ZN(n667) );
  INV_X1 U639 ( .A(n575), .ZN(n537) );
  NAND2_X1 U640 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U641 ( .A1(n631), .A2(n539), .ZN(n540) );
  XNOR2_X1 U642 ( .A(n540), .B(KEYINPUT103), .ZN(n541) );
  NAND2_X1 U643 ( .A1(n542), .A2(n541), .ZN(n545) );
  INV_X1 U644 ( .A(KEYINPUT64), .ZN(n543) );
  XNOR2_X1 U645 ( .A(n543), .B(KEYINPUT45), .ZN(n544) );
  INV_X1 U646 ( .A(n730), .ZN(n603) );
  XNOR2_X1 U647 ( .A(n598), .B(n549), .ZN(n566) );
  INV_X1 U648 ( .A(n566), .ZN(n663) );
  NAND2_X1 U649 ( .A1(n663), .A2(n662), .ZN(n666) );
  INV_X1 U650 ( .A(n550), .ZN(n665) );
  OR2_X1 U651 ( .A1(n743), .A2(n553), .ZN(n554) );
  NOR2_X1 U652 ( .A1(G900), .A2(n554), .ZN(n555) );
  NOR2_X1 U653 ( .A1(n556), .A2(n555), .ZN(n560) );
  XNOR2_X1 U654 ( .A(n562), .B(KEYINPUT78), .ZN(n565) );
  NAND2_X1 U655 ( .A1(n677), .A2(n662), .ZN(n563) );
  XOR2_X1 U656 ( .A(KEYINPUT30), .B(n563), .Z(n564) );
  NOR2_X1 U657 ( .A1(KEYINPUT81), .A2(n355), .ZN(n573) );
  INV_X1 U658 ( .A(KEYINPUT47), .ZN(n574) );
  XNOR2_X1 U659 ( .A(n579), .B(n578), .ZN(n589) );
  NAND2_X1 U660 ( .A1(n674), .A2(n662), .ZN(n582) );
  NAND2_X1 U661 ( .A1(n644), .A2(n580), .ZN(n581) );
  NOR2_X1 U662 ( .A1(n582), .A2(n581), .ZN(n595) );
  NAND2_X1 U663 ( .A1(n595), .A2(n391), .ZN(n584) );
  NOR2_X1 U664 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U665 ( .A(KEYINPUT36), .B(n585), .ZN(n587) );
  NAND2_X1 U666 ( .A1(n587), .A2(n586), .ZN(n652) );
  NAND2_X1 U667 ( .A1(n591), .A2(n590), .ZN(n593) );
  XOR2_X1 U668 ( .A(KEYINPUT48), .B(KEYINPUT72), .Z(n592) );
  NAND2_X1 U669 ( .A1(n595), .A2(n594), .ZN(n596) );
  OR2_X1 U670 ( .A1(n596), .A2(n680), .ZN(n597) );
  XNOR2_X1 U671 ( .A(n597), .B(KEYINPUT43), .ZN(n599) );
  AND2_X1 U672 ( .A1(n599), .A2(n598), .ZN(n656) );
  INV_X1 U673 ( .A(n656), .ZN(n601) );
  NAND2_X1 U674 ( .A1(n640), .A2(n600), .ZN(n655) );
  AND2_X1 U675 ( .A1(n601), .A2(n655), .ZN(n602) );
  NAND2_X1 U676 ( .A1(n603), .A2(n403), .ZN(n608) );
  INV_X1 U677 ( .A(KEYINPUT85), .ZN(n604) );
  XNOR2_X1 U678 ( .A(n605), .B(n604), .ZN(n606) );
  NAND2_X1 U679 ( .A1(n606), .A2(KEYINPUT2), .ZN(n607) );
  NAND2_X1 U680 ( .A1(n608), .A2(n607), .ZN(n610) );
  AND2_X2 U681 ( .A1(n610), .A2(n660), .ZN(n711) );
  NAND2_X1 U682 ( .A1(n711), .A2(G210), .ZN(n615) );
  XOR2_X1 U683 ( .A(KEYINPUT118), .B(KEYINPUT54), .Z(n613) );
  XNOR2_X1 U684 ( .A(n611), .B(KEYINPUT55), .ZN(n612) );
  XNOR2_X1 U685 ( .A(n613), .B(n612), .ZN(n614) );
  XNOR2_X1 U686 ( .A(n615), .B(n614), .ZN(n617) );
  INV_X1 U687 ( .A(G952), .ZN(n616) );
  AND2_X1 U688 ( .A1(n616), .A2(G953), .ZN(n725) );
  NOR2_X1 U689 ( .A1(n617), .A2(n725), .ZN(n620) );
  INV_X1 U690 ( .A(KEYINPUT119), .ZN(n618) );
  XNOR2_X1 U691 ( .A(n620), .B(n619), .ZN(G51) );
  XOR2_X1 U692 ( .A(G122), .B(KEYINPUT125), .Z(n621) );
  XNOR2_X1 U693 ( .A(n622), .B(n621), .ZN(G24) );
  NAND2_X1 U694 ( .A1(n711), .A2(G472), .ZN(n627) );
  XNOR2_X1 U695 ( .A(KEYINPUT89), .B(KEYINPUT107), .ZN(n623) );
  XNOR2_X1 U696 ( .A(n623), .B(KEYINPUT62), .ZN(n624) );
  XNOR2_X1 U697 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U698 ( .A(n627), .B(n626), .ZN(n628) );
  NOR2_X1 U699 ( .A1(n628), .A2(n725), .ZN(n630) );
  XOR2_X1 U700 ( .A(KEYINPUT88), .B(KEYINPUT63), .Z(n629) );
  XNOR2_X1 U701 ( .A(n630), .B(n629), .ZN(G57) );
  XNOR2_X1 U702 ( .A(G101), .B(n631), .ZN(G3) );
  INV_X1 U703 ( .A(n644), .ZN(n647) );
  NOR2_X1 U704 ( .A1(n634), .A2(n647), .ZN(n632) );
  XOR2_X1 U705 ( .A(KEYINPUT108), .B(n632), .Z(n633) );
  XNOR2_X1 U706 ( .A(G104), .B(n633), .ZN(G6) );
  INV_X1 U707 ( .A(n640), .ZN(n650) );
  NOR2_X1 U708 ( .A1(n634), .A2(n650), .ZN(n638) );
  XOR2_X1 U709 ( .A(KEYINPUT26), .B(KEYINPUT27), .Z(n636) );
  XNOR2_X1 U710 ( .A(G107), .B(KEYINPUT109), .ZN(n635) );
  XNOR2_X1 U711 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U712 ( .A(n638), .B(n637), .ZN(G9) );
  XOR2_X1 U713 ( .A(G110), .B(n639), .Z(G12) );
  XOR2_X1 U714 ( .A(G128), .B(KEYINPUT29), .Z(n642) );
  NAND2_X1 U715 ( .A1(n355), .A2(n640), .ZN(n641) );
  XNOR2_X1 U716 ( .A(n642), .B(n641), .ZN(G30) );
  XOR2_X1 U717 ( .A(G143), .B(n643), .Z(G45) );
  NAND2_X1 U718 ( .A1(n355), .A2(n644), .ZN(n645) );
  XNOR2_X1 U719 ( .A(n645), .B(KEYINPUT110), .ZN(n646) );
  XNOR2_X1 U720 ( .A(G146), .B(n646), .ZN(G48) );
  NOR2_X1 U721 ( .A1(n647), .A2(n649), .ZN(n648) );
  XOR2_X1 U722 ( .A(G113), .B(n648), .Z(G15) );
  NOR2_X1 U723 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U724 ( .A(G116), .B(n651), .Z(G18) );
  XNOR2_X1 U725 ( .A(KEYINPUT111), .B(KEYINPUT37), .ZN(n653) );
  XNOR2_X1 U726 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U727 ( .A(G125), .B(n654), .ZN(G27) );
  XNOR2_X1 U728 ( .A(G134), .B(n655), .ZN(G36) );
  XOR2_X1 U729 ( .A(G140), .B(n656), .Z(G42) );
  NOR2_X1 U730 ( .A1(n603), .A2(KEYINPUT2), .ZN(n659) );
  NOR2_X1 U731 ( .A1(n742), .A2(KEYINPUT2), .ZN(n657) );
  XNOR2_X1 U732 ( .A(n657), .B(KEYINPUT84), .ZN(n658) );
  NOR2_X1 U733 ( .A1(n659), .A2(n658), .ZN(n661) );
  NAND2_X1 U734 ( .A1(n661), .A2(n660), .ZN(n702) );
  NOR2_X1 U735 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U736 ( .A1(n665), .A2(n664), .ZN(n670) );
  NOR2_X1 U737 ( .A1(n667), .A2(n666), .ZN(n668) );
  XOR2_X1 U738 ( .A(KEYINPUT115), .B(n668), .Z(n669) );
  NOR2_X1 U739 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U740 ( .A(n671), .B(KEYINPUT116), .ZN(n672) );
  NOR2_X1 U741 ( .A1(n672), .A2(n698), .ZN(n673) );
  XNOR2_X1 U742 ( .A(n673), .B(KEYINPUT117), .ZN(n692) );
  NOR2_X1 U743 ( .A1(n675), .A2(n674), .ZN(n676) );
  XOR2_X1 U744 ( .A(KEYINPUT49), .B(n676), .Z(n678) );
  NOR2_X1 U745 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U746 ( .A(n679), .B(KEYINPUT112), .Z(n684) );
  NOR2_X1 U747 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U748 ( .A(KEYINPUT50), .B(n682), .ZN(n683) );
  NOR2_X1 U749 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U750 ( .A(n685), .B(KEYINPUT113), .ZN(n687) );
  NAND2_X1 U751 ( .A1(n687), .A2(n686), .ZN(n689) );
  XOR2_X1 U752 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n688) );
  XNOR2_X1 U753 ( .A(n689), .B(n688), .ZN(n690) );
  NAND2_X1 U754 ( .A1(n690), .A2(n696), .ZN(n691) );
  NAND2_X1 U755 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U756 ( .A(KEYINPUT52), .B(n693), .Z(n694) );
  NOR2_X1 U757 ( .A1(n695), .A2(n694), .ZN(n700) );
  INV_X1 U758 ( .A(n696), .ZN(n697) );
  NOR2_X1 U759 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U760 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U761 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U762 ( .A1(n703), .A2(G953), .ZN(n704) );
  XNOR2_X1 U763 ( .A(n704), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U764 ( .A1(n720), .A2(G469), .ZN(n709) );
  XNOR2_X1 U765 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n705) );
  XNOR2_X1 U766 ( .A(n705), .B(KEYINPUT57), .ZN(n706) );
  XNOR2_X1 U767 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U768 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X1 U769 ( .A1(n725), .A2(n710), .ZN(G54) );
  NAND2_X1 U770 ( .A1(n711), .A2(G475), .ZN(n714) );
  XOR2_X1 U771 ( .A(n712), .B(KEYINPUT59), .Z(n713) );
  XNOR2_X1 U772 ( .A(n714), .B(n713), .ZN(n715) );
  XNOR2_X1 U773 ( .A(n716), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U774 ( .A1(n720), .A2(G478), .ZN(n718) );
  XNOR2_X1 U775 ( .A(n718), .B(n717), .ZN(n719) );
  NOR2_X1 U776 ( .A1(n725), .A2(n719), .ZN(G63) );
  NAND2_X1 U777 ( .A1(n720), .A2(G217), .ZN(n723) );
  XOR2_X1 U778 ( .A(n721), .B(KEYINPUT121), .Z(n722) );
  XNOR2_X1 U779 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U780 ( .A1(n725), .A2(n724), .ZN(G66) );
  XOR2_X1 U781 ( .A(n726), .B(G110), .Z(n727) );
  XNOR2_X1 U782 ( .A(KEYINPUT124), .B(n727), .ZN(n729) );
  NAND2_X1 U783 ( .A1(n729), .A2(n728), .ZN(n739) );
  NOR2_X1 U784 ( .A1(n730), .A2(G953), .ZN(n731) );
  XOR2_X1 U785 ( .A(KEYINPUT123), .B(n731), .Z(n737) );
  XOR2_X1 U786 ( .A(KEYINPUT122), .B(KEYINPUT61), .Z(n733) );
  NAND2_X1 U787 ( .A1(G224), .A2(G953), .ZN(n732) );
  XNOR2_X1 U788 ( .A(n733), .B(n732), .ZN(n734) );
  NOR2_X1 U789 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U790 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U791 ( .A(n739), .B(n738), .ZN(G69) );
  XNOR2_X1 U792 ( .A(n740), .B(n741), .ZN(n745) );
  XNOR2_X1 U793 ( .A(n742), .B(n745), .ZN(n744) );
  NAND2_X1 U794 ( .A1(n744), .A2(n743), .ZN(n749) );
  XOR2_X1 U795 ( .A(n745), .B(G227), .Z(n746) );
  NAND2_X1 U796 ( .A1(n746), .A2(G900), .ZN(n747) );
  NAND2_X1 U797 ( .A1(n747), .A2(G953), .ZN(n748) );
  NAND2_X1 U798 ( .A1(n749), .A2(n748), .ZN(G72) );
  XOR2_X1 U799 ( .A(G137), .B(n750), .Z(G39) );
  XOR2_X1 U800 ( .A(G119), .B(KEYINPUT126), .Z(n751) );
  XNOR2_X1 U801 ( .A(n752), .B(n751), .ZN(G21) );
  XOR2_X1 U802 ( .A(G131), .B(n753), .Z(G33) );
endmodule

