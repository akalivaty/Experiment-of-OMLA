//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 0 1 0 0 1 1 0 0 0 1 0 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n776, new_n777, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT83), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  XNOR2_X1  g003(.A(G116), .B(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT5), .ZN(new_n191));
  INV_X1    g005(.A(G113), .ZN(new_n192));
  INV_X1    g006(.A(G116), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G119), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT5), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n192), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n192), .A2(KEYINPUT2), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G113), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  AOI22_X1  g014(.A1(new_n191), .A2(new_n196), .B1(new_n190), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G104), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT3), .B1(new_n202), .B2(G107), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n204));
  INV_X1    g018(.A(G107), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(G104), .ZN(new_n206));
  INV_X1    g020(.A(G101), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n202), .A2(G107), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n203), .A2(new_n206), .A3(new_n207), .A4(new_n208), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n202), .A2(G107), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n205), .A2(G104), .ZN(new_n211));
  OAI21_X1  g025(.A(G101), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n201), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(G110), .B(G122), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n203), .A2(new_n206), .A3(new_n208), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n216), .A2(G101), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n209), .A2(KEYINPUT4), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G119), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n220), .A2(G116), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n197), .B(new_n199), .C1(new_n194), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n200), .A2(new_n190), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT4), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n216), .A2(new_n225), .A3(G101), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n214), .B(new_n215), .C1(new_n219), .C2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n209), .A2(new_n212), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n201), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n215), .B(KEYINPUT8), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n220), .A2(G116), .ZN(new_n232));
  OAI21_X1  g046(.A(G113), .B1(new_n232), .B2(KEYINPUT5), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT79), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n233), .A2(new_n234), .B1(new_n190), .B2(KEYINPUT5), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n196), .A2(KEYINPUT79), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n235), .A2(new_n236), .B1(new_n190), .B2(new_n200), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n230), .B(new_n231), .C1(new_n237), .C2(new_n229), .ZN(new_n238));
  INV_X1    g052(.A(G128), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(KEYINPUT1), .ZN(new_n240));
  INV_X1    g054(.A(G143), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G146), .ZN(new_n242));
  INV_X1    g056(.A(G146), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G143), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n240), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT67), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(G143), .B(G146), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(KEYINPUT67), .A3(new_n240), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT64), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(new_n243), .A3(G143), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT64), .B1(new_n241), .B2(G146), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n241), .A2(G146), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT1), .B1(new_n241), .B2(G146), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(G128), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n239), .A2(KEYINPUT68), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n256), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n255), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G125), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n250), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT0), .B(G128), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n251), .B1(new_n243), .B2(G143), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n244), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n264), .B1(new_n266), .B2(new_n252), .ZN(new_n267));
  AND2_X1   g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n248), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(G125), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G224), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n271), .A2(G953), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n263), .A2(new_n270), .A3(KEYINPUT7), .A4(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n238), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT80), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n263), .A2(new_n276), .A3(new_n270), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n250), .A2(new_n261), .A3(KEYINPUT80), .A4(new_n262), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n273), .A2(KEYINPUT7), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT81), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n278), .A2(new_n279), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT81), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n263), .A2(new_n270), .A3(new_n276), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n275), .B1(new_n281), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n228), .B1(new_n286), .B2(KEYINPUT82), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT82), .ZN(new_n288));
  AOI211_X1 g102(.A(new_n288), .B(new_n275), .C1(new_n281), .C2(new_n285), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n189), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n214), .B1(new_n219), .B2(new_n227), .ZN(new_n291));
  INV_X1    g105(.A(new_n215), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(KEYINPUT6), .A3(new_n228), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT6), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n291), .A2(new_n295), .A3(new_n292), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n263), .A2(new_n270), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n272), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n263), .A2(new_n273), .A3(new_n270), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n294), .A2(new_n296), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT78), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT78), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n294), .A2(new_n303), .A3(new_n300), .A4(new_n296), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n188), .B1(new_n290), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n228), .ZN(new_n307));
  INV_X1    g121(.A(new_n275), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n277), .A2(KEYINPUT81), .A3(new_n280), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n283), .B1(new_n282), .B2(new_n284), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n307), .B1(new_n311), .B2(new_n288), .ZN(new_n312));
  INV_X1    g126(.A(new_n289), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n302), .A2(new_n304), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n314), .A2(new_n189), .A3(new_n187), .A4(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n306), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(G214), .B1(G237), .B2(G902), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT9), .B(G234), .ZN(new_n319));
  OAI21_X1  g133(.A(G221), .B1(new_n319), .B2(G902), .ZN(new_n320));
  INV_X1    g134(.A(G469), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n239), .B1(new_n244), .B2(KEYINPUT1), .ZN(new_n322));
  OR2_X1    g136(.A1(new_n322), .A2(new_n248), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n229), .B1(new_n250), .B2(new_n323), .ZN(new_n324));
  XOR2_X1   g138(.A(KEYINPUT75), .B(KEYINPUT10), .Z(new_n325));
  OR2_X1    g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT11), .ZN(new_n327));
  INV_X1    g141(.A(G134), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n327), .B1(new_n328), .B2(G137), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(G137), .ZN(new_n330));
  INV_X1    g144(.A(G137), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(KEYINPUT11), .A3(G134), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n329), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G131), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT66), .ZN(new_n335));
  INV_X1    g149(.A(G131), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n329), .A2(new_n332), .A3(new_n336), .A4(new_n330), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n334), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n333), .A2(KEYINPUT66), .A3(G131), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n264), .ZN(new_n341));
  AOI22_X1  g155(.A1(new_n255), .A2(new_n341), .B1(new_n248), .B2(new_n268), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n342), .B(new_n226), .C1(new_n217), .C2(new_n218), .ZN(new_n343));
  AOI21_X1  g157(.A(KEYINPUT67), .B1(new_n248), .B2(new_n240), .ZN(new_n344));
  AND4_X1   g158(.A1(KEYINPUT67), .A2(new_n240), .A3(new_n242), .A4(new_n244), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n241), .A2(KEYINPUT64), .A3(G146), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n346), .B1(new_n244), .B2(new_n265), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n239), .A2(KEYINPUT68), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n257), .A2(G128), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n348), .A2(new_n349), .B1(new_n244), .B2(KEYINPUT1), .ZN(new_n350));
  OAI22_X1  g164(.A1(new_n344), .A2(new_n345), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(KEYINPUT10), .A3(new_n213), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n326), .A2(new_n340), .A3(new_n343), .A4(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(G110), .B(G140), .ZN(new_n354));
  INV_X1    g168(.A(G953), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n355), .A2(G227), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n354), .B(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n250), .A2(new_n323), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n213), .ZN(new_n361));
  AOI22_X1  g175(.A1(new_n247), .A2(new_n249), .B1(new_n255), .B2(new_n260), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n229), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n340), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT77), .B1(new_n364), .B2(KEYINPUT12), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n338), .A2(new_n339), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n351), .A2(new_n213), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n366), .B1(new_n367), .B2(new_n324), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT77), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT12), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  OAI211_X1 g186(.A(KEYINPUT12), .B(new_n366), .C1(new_n367), .C2(new_n324), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT76), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT76), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n364), .A2(new_n375), .A3(KEYINPUT12), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n359), .B1(new_n372), .B2(new_n377), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n352), .B(new_n343), .C1(new_n324), .C2(new_n325), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n366), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n358), .B1(new_n380), .B2(new_n353), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n321), .B(new_n189), .C1(new_n378), .C2(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n321), .A2(new_n189), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n359), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n380), .ZN(new_n386));
  INV_X1    g200(.A(new_n353), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n387), .B1(new_n372), .B2(new_n377), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n386), .B1(new_n388), .B2(new_n358), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n382), .B(new_n384), .C1(new_n389), .C2(new_n321), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n317), .A2(new_n318), .A3(new_n320), .A4(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(G475), .A2(G902), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT85), .ZN(new_n393));
  INV_X1    g207(.A(G237), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(new_n355), .A3(G214), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n241), .ZN(new_n396));
  NOR2_X1   g210(.A1(G237), .A2(G953), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(G143), .A3(G214), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n393), .B1(new_n399), .B2(G131), .ZN(new_n400));
  AOI211_X1 g214(.A(KEYINPUT85), .B(new_n336), .C1(new_n396), .C2(new_n398), .ZN(new_n401));
  OAI21_X1  g215(.A(KEYINPUT17), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AND4_X1   g216(.A1(G143), .A2(new_n394), .A3(new_n355), .A4(G214), .ZN(new_n403));
  AOI21_X1  g217(.A(G143), .B1(new_n397), .B2(G214), .ZN(new_n404));
  OAI21_X1  g218(.A(G131), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT85), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT17), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n393), .B(G131), .C1(new_n403), .C2(new_n404), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n396), .A2(new_n336), .A3(new_n398), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n406), .A2(new_n407), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n262), .A2(G140), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT16), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G140), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G125), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n262), .A2(G140), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n413), .B1(new_n417), .B2(new_n412), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n243), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n413), .B(G146), .C1(new_n417), .C2(new_n412), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n402), .A2(new_n410), .A3(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(G113), .B(G122), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n424), .B(new_n202), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n414), .A2(G125), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT84), .B1(new_n411), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT84), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n415), .A2(new_n416), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n427), .A2(G146), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n417), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n243), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(KEYINPUT18), .A2(G131), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n396), .A2(new_n398), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n434), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n436), .B1(new_n403), .B2(new_n404), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n433), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n423), .A2(new_n425), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n406), .A2(new_n408), .A3(new_n409), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n427), .A2(KEYINPUT19), .A3(new_n429), .ZN(new_n441));
  OR2_X1    g255(.A1(new_n417), .A2(KEYINPUT19), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n441), .A2(new_n243), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n440), .A2(new_n420), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n425), .B1(new_n444), .B2(new_n438), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT86), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n439), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n437), .A2(new_n435), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n448), .B1(new_n432), .B2(new_n430), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n443), .A2(new_n420), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n449), .B1(new_n450), .B2(new_n440), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n451), .A2(KEYINPUT86), .A3(new_n425), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n392), .B1(new_n447), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT20), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT87), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n453), .A2(KEYINPUT87), .A3(KEYINPUT20), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT20), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n458), .B(new_n392), .C1(new_n447), .C2(new_n452), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n456), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n423), .A2(new_n438), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n425), .A2(KEYINPUT88), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n189), .B1(new_n461), .B2(new_n462), .ZN(new_n465));
  OAI21_X1  g279(.A(G475), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT14), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(new_n193), .A3(G122), .ZN(new_n468));
  INV_X1    g282(.A(G122), .ZN(new_n469));
  AOI21_X1  g283(.A(KEYINPUT14), .B1(new_n469), .B2(G116), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n469), .A2(G116), .ZN(new_n471));
  OAI211_X1 g285(.A(KEYINPUT89), .B(new_n468), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n467), .B1(new_n193), .B2(G122), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT89), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n193), .A2(G122), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n472), .A2(G107), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT90), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n348), .A2(new_n349), .A3(G143), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n241), .A2(G128), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(G134), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n479), .A2(new_n328), .A3(new_n480), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(G116), .B(G122), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n205), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT90), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n472), .A2(new_n487), .A3(G107), .A4(new_n476), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n478), .A2(new_n484), .A3(new_n486), .A4(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT13), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n480), .B(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n479), .ZN(new_n492));
  OAI21_X1  g306(.A(G134), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n485), .B(new_n205), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n483), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n489), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G217), .ZN(new_n497));
  NOR3_X1   g311(.A1(new_n319), .A2(new_n497), .A3(G953), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n498), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n489), .A2(new_n495), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n499), .A2(new_n189), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT91), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(G478), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT92), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n506), .A2(KEYINPUT15), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(KEYINPUT15), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n499), .A2(KEYINPUT91), .A3(new_n189), .A4(new_n501), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n504), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  OR2_X1    g326(.A1(new_n502), .A2(new_n510), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(G234), .A2(G237), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n515), .A2(G952), .A3(new_n355), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT21), .B(G898), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(KEYINPUT93), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n515), .A2(G902), .A3(G953), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n516), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n514), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n460), .A2(new_n466), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT94), .B1(new_n391), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT71), .ZN(new_n525));
  NOR2_X1   g339(.A1(G472), .A2(G902), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT26), .B(G101), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n397), .A2(G210), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n530), .B(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT28), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT69), .ZN(new_n534));
  INV_X1    g348(.A(new_n330), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n328), .A2(G137), .ZN(new_n536));
  OAI21_X1  g350(.A(G131), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n337), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n351), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n338), .A2(new_n339), .A3(new_n342), .ZN(new_n541));
  INV_X1    g355(.A(new_n224), .ZN(new_n542));
  AND4_X1   g356(.A1(new_n534), .A2(new_n540), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n224), .B1(new_n351), .B2(new_n539), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n534), .B1(new_n544), .B2(new_n541), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT65), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n547), .B1(new_n267), .B2(new_n269), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n255), .A2(new_n341), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n248), .A2(new_n268), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(KEYINPUT65), .A3(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n548), .A2(new_n551), .A3(new_n339), .A4(new_n338), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n542), .B1(new_n552), .B2(new_n540), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n533), .B1(new_n546), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(KEYINPUT28), .B1(new_n544), .B2(new_n541), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n532), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n540), .A2(new_n541), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT30), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT30), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n552), .A2(new_n560), .A3(new_n540), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n224), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n338), .A2(new_n339), .A3(new_n342), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n542), .B1(new_n362), .B2(new_n538), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT69), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n544), .A2(new_n534), .A3(new_n541), .ZN(new_n567));
  INV_X1    g381(.A(new_n532), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n563), .A2(new_n569), .A3(KEYINPUT31), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT31), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n542), .B1(new_n559), .B2(new_n561), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n527), .B1(new_n557), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n525), .B1(new_n576), .B2(KEYINPUT32), .ZN(new_n577));
  INV_X1    g391(.A(new_n556), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT29), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n532), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n566), .A2(new_n567), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n542), .B1(new_n540), .B2(new_n541), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT72), .ZN(new_n583));
  OR2_X1    g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n583), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n581), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n578), .B(new_n580), .C1(new_n586), .C2(new_n533), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n189), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n552), .A2(new_n540), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n566), .B(new_n567), .C1(new_n589), .C2(new_n542), .ZN(new_n590));
  AOI211_X1 g404(.A(new_n556), .B(new_n532), .C1(new_n590), .C2(KEYINPUT28), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n532), .B1(new_n572), .B2(new_n581), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n579), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(G472), .B1(new_n588), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n576), .A2(KEYINPUT32), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT32), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT28), .B1(new_n581), .B2(new_n553), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n578), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n599), .A2(new_n532), .B1(new_n570), .B2(new_n574), .ZN(new_n600));
  OAI211_X1 g414(.A(KEYINPUT71), .B(new_n597), .C1(new_n600), .C2(new_n527), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n577), .A2(new_n595), .A3(new_n596), .A4(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n497), .B1(G234), .B2(new_n189), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n348), .A2(new_n349), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n605), .A2(KEYINPUT23), .A3(G119), .ZN(new_n606));
  AOI21_X1  g420(.A(KEYINPUT23), .B1(new_n239), .B2(G119), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n239), .A2(G119), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT24), .B(G110), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT73), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n608), .B1(new_n605), .B2(G119), .ZN(new_n613));
  OAI22_X1  g427(.A1(new_n610), .A2(G110), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n614), .A2(new_n420), .A3(new_n432), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n610), .A2(G110), .B1(new_n612), .B2(new_n613), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n421), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT22), .B(G137), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n355), .A2(G221), .A3(G234), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(KEYINPUT74), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n615), .A2(new_n617), .A3(new_n621), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(new_n189), .A3(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT25), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n624), .A2(KEYINPUT25), .A3(new_n189), .A4(new_n625), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n604), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n624), .A2(new_n625), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n603), .A2(G902), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n602), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n523), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n390), .A2(new_n320), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT94), .ZN(new_n638));
  INV_X1    g452(.A(new_n318), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n639), .B1(new_n306), .B2(new_n316), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n636), .A2(new_n637), .A3(new_n638), .A4(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n524), .A2(new_n635), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT95), .B(G101), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G3));
  INV_X1    g458(.A(new_n187), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n645), .B1(new_n290), .B2(new_n305), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n639), .B1(new_n646), .B2(new_n316), .ZN(new_n647));
  INV_X1    g461(.A(new_n521), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n460), .A2(new_n466), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n504), .A2(new_n505), .A3(new_n511), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(KEYINPUT98), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT98), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n504), .A2(new_n653), .A3(new_n505), .A4(new_n511), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g469(.A1(new_n500), .A2(KEYINPUT97), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n496), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n496), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n657), .A2(KEYINPUT33), .A3(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n505), .A2(G902), .ZN(new_n660));
  INV_X1    g474(.A(new_n501), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n500), .B1(new_n489), .B2(new_n495), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n661), .A2(KEYINPUT33), .A3(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT96), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR4_X1   g479(.A1(new_n661), .A2(new_n662), .A3(KEYINPUT96), .A4(KEYINPUT33), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n659), .B(new_n660), .C1(new_n665), .C2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n655), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n650), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n649), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n390), .A2(new_n634), .A3(new_n320), .ZN(new_n671));
  OAI21_X1  g485(.A(G472), .B1(new_n600), .B2(G902), .ZN(new_n672));
  INV_X1    g486(.A(new_n576), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n670), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT34), .B(G104), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G6));
  NAND3_X1  g492(.A1(new_n456), .A2(KEYINPUT99), .A3(new_n457), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT99), .ZN(new_n680));
  OAI21_X1  g494(.A(KEYINPUT86), .B1(new_n451), .B2(new_n425), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n445), .A2(new_n446), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(new_n682), .A3(new_n439), .ZN(new_n683));
  AOI211_X1 g497(.A(new_n455), .B(new_n458), .C1(new_n683), .C2(new_n392), .ZN(new_n684));
  AOI21_X1  g498(.A(KEYINPUT87), .B1(new_n453), .B2(KEYINPUT20), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n680), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n679), .A2(new_n686), .A3(new_n459), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n687), .A2(new_n466), .A3(new_n514), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n649), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n675), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT35), .B(G107), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G9));
  INV_X1    g506(.A(KEYINPUT36), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n622), .A2(new_n693), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n618), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n618), .A2(new_n694), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n697), .A2(new_n632), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n630), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n674), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n524), .A2(new_n641), .A3(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT37), .B(G110), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G12));
  INV_X1    g517(.A(new_n516), .ZN(new_n704));
  INV_X1    g518(.A(new_n520), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n704), .B1(new_n705), .B2(G900), .ZN(new_n706));
  AND4_X1   g520(.A1(new_n466), .A2(new_n687), .A3(new_n514), .A4(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n646), .A2(new_n316), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n318), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n630), .A2(new_n698), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n390), .A2(new_n710), .A3(new_n320), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n707), .A2(new_n602), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G128), .ZN(G30));
  NAND2_X1  g528(.A1(new_n390), .A2(new_n320), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n706), .B(KEYINPUT39), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(KEYINPUT40), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n577), .A2(new_n601), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n572), .A2(new_n573), .ZN(new_n721));
  OAI21_X1  g535(.A(KEYINPUT101), .B1(new_n586), .B2(new_n568), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT101), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n582), .B(KEYINPUT72), .ZN(new_n724));
  OAI211_X1 g538(.A(new_n723), .B(new_n532), .C1(new_n724), .C2(new_n581), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n721), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT102), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n189), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  AOI211_X1 g542(.A(KEYINPUT102), .B(new_n721), .C1(new_n722), .C2(new_n725), .ZN(new_n729));
  OAI21_X1  g543(.A(G472), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n720), .A2(new_n730), .A3(new_n596), .ZN(new_n731));
  XOR2_X1   g545(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n732));
  XNOR2_X1  g546(.A(new_n317), .B(new_n732), .ZN(new_n733));
  AOI22_X1  g547(.A1(new_n460), .A2(new_n466), .B1(new_n513), .B2(new_n512), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n734), .A2(new_n318), .A3(new_n699), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n719), .A2(new_n731), .A3(new_n733), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G143), .ZN(G45));
  INV_X1    g551(.A(new_n459), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n684), .A2(new_n685), .A3(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n466), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n668), .B(new_n706), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT103), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT103), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n650), .A2(new_n743), .A3(new_n668), .A4(new_n706), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n712), .A2(new_n742), .A3(new_n602), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G146), .ZN(G48));
  INV_X1    g560(.A(new_n649), .ZN(new_n747));
  INV_X1    g561(.A(new_n669), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n189), .B1(new_n378), .B2(new_n381), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(G469), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n751), .A2(new_n320), .A3(new_n382), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n602), .A2(new_n634), .A3(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  XOR2_X1   g568(.A(KEYINPUT41), .B(G113), .Z(new_n755));
  XNOR2_X1  g569(.A(new_n754), .B(new_n755), .ZN(G15));
  INV_X1    g570(.A(new_n753), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n689), .ZN(new_n758));
  XOR2_X1   g572(.A(KEYINPUT104), .B(G116), .Z(new_n759));
  XNOR2_X1  g573(.A(new_n758), .B(new_n759), .ZN(G18));
  AND2_X1   g574(.A1(new_n647), .A2(new_n752), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n523), .A2(new_n699), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(new_n602), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G119), .ZN(G21));
  INV_X1    g578(.A(new_n634), .ZN(new_n765));
  INV_X1    g579(.A(G472), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n557), .A2(new_n575), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n766), .B1(new_n767), .B2(new_n189), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n578), .B1(new_n586), .B2(new_n533), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n532), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n527), .B1(new_n770), .B2(new_n575), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n765), .A2(new_n768), .A3(new_n771), .ZN(new_n772));
  AND4_X1   g586(.A1(new_n648), .A2(new_n751), .A3(new_n320), .A4(new_n382), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n772), .A2(new_n734), .A3(new_n647), .A4(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G122), .ZN(G24));
  NOR3_X1   g589(.A1(new_n768), .A2(new_n771), .A3(new_n699), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n742), .A2(new_n761), .A3(new_n744), .A4(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G125), .ZN(G27));
  INV_X1    g592(.A(KEYINPUT42), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n742), .A2(new_n744), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n306), .A2(new_n318), .A3(new_n316), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n602), .A2(new_n634), .A3(new_n637), .A4(new_n781), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n779), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n595), .A2(new_n596), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n673), .A2(new_n597), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n765), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n306), .A2(new_n318), .A3(new_n316), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n715), .A2(new_n787), .A3(new_n779), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n786), .A2(new_n788), .A3(new_n744), .A4(new_n742), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n783), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G131), .ZN(G33));
  INV_X1    g605(.A(KEYINPUT105), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n715), .A2(new_n787), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n635), .A2(new_n707), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n687), .A2(new_n466), .A3(new_n514), .A4(new_n706), .ZN(new_n795));
  OAI21_X1  g609(.A(KEYINPUT105), .B1(new_n782), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G134), .ZN(G36));
  AOI21_X1  g612(.A(new_n650), .B1(new_n655), .B2(new_n667), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT43), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n699), .B1(new_n672), .B2(new_n673), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT44), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  XOR2_X1   g618(.A(new_n804), .B(KEYINPUT107), .Z(new_n805));
  INV_X1    g619(.A(KEYINPUT45), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n389), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n321), .B1(new_n389), .B2(new_n806), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n809), .A2(new_n383), .ZN(new_n810));
  OR3_X1    g624(.A1(new_n810), .A2(KEYINPUT106), .A3(KEYINPUT46), .ZN(new_n811));
  OAI21_X1  g625(.A(KEYINPUT106), .B1(new_n810), .B2(KEYINPUT46), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n810), .A2(KEYINPUT46), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n811), .A2(new_n382), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n320), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n717), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n787), .B1(new_n802), .B2(new_n803), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n805), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  XOR2_X1   g632(.A(KEYINPUT108), .B(G137), .Z(new_n819));
  XNOR2_X1  g633(.A(new_n818), .B(new_n819), .ZN(G39));
  NAND3_X1  g634(.A1(new_n814), .A2(KEYINPUT109), .A3(new_n320), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT109), .B1(new_n814), .B2(new_n320), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT47), .ZN(new_n824));
  OAI22_X1  g638(.A1(new_n822), .A2(new_n823), .B1(KEYINPUT110), .B2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n823), .ZN(new_n826));
  XNOR2_X1  g640(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n826), .A2(new_n821), .A3(new_n828), .ZN(new_n829));
  NOR4_X1   g643(.A1(new_n780), .A2(new_n602), .A3(new_n634), .A4(new_n787), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n825), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT111), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n831), .B(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(G140), .ZN(G42));
  NAND2_X1  g648(.A1(new_n781), .A2(new_n752), .ZN(new_n835));
  OR4_X1    g649(.A1(new_n765), .A2(new_n731), .A3(new_n704), .A4(new_n835), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n836), .A2(new_n650), .A3(new_n668), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n800), .A2(new_n516), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT118), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT118), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n800), .A2(new_n840), .A3(new_n516), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n835), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n837), .B1(new_n842), .B2(new_n776), .ZN(new_n843));
  INV_X1    g657(.A(new_n772), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n844), .B1(new_n839), .B2(new_n841), .ZN(new_n845));
  INV_X1    g659(.A(new_n752), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n733), .A2(new_n318), .A3(new_n846), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n845), .A2(KEYINPUT50), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT50), .B1(new_n845), .B2(new_n847), .ZN(new_n849));
  OAI211_X1 g663(.A(KEYINPUT51), .B(new_n843), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n751), .A2(new_n382), .ZN(new_n851));
  INV_X1    g665(.A(new_n320), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n825), .ZN(new_n854));
  INV_X1    g668(.A(new_n829), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n845), .A2(new_n781), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n850), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI211_X1 g672(.A(G952), .B(new_n355), .C1(new_n836), .C2(new_n669), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(new_n845), .B2(new_n761), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n842), .A2(new_n786), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n861), .A2(KEYINPUT48), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(KEYINPUT48), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n860), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n858), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n843), .B1(new_n848), .B2(new_n849), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n867), .B1(new_n854), .B2(new_n855), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n825), .A2(new_n829), .A3(KEYINPUT119), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n868), .A2(new_n869), .A3(new_n853), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n866), .B1(new_n870), .B2(new_n857), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n865), .B1(new_n871), .B2(KEYINPUT51), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n742), .A2(new_n744), .A3(new_n776), .ZN(new_n873));
  AND4_X1   g687(.A1(new_n513), .A2(new_n710), .A3(new_n512), .A4(new_n706), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(new_n602), .A3(new_n466), .A4(new_n687), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n793), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n790), .A2(new_n797), .A3(new_n877), .ZN(new_n878));
  AOI211_X1 g692(.A(new_n521), .B(new_n639), .C1(new_n306), .C2(new_n316), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n748), .A2(new_n675), .A3(new_n879), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n763), .A2(new_n880), .A3(new_n774), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n757), .B1(new_n689), .B2(new_n670), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n640), .A2(new_n648), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n460), .A2(new_n466), .A3(new_n514), .ZN(new_n884));
  OAI21_X1  g698(.A(KEYINPUT112), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT112), .ZN(new_n886));
  INV_X1    g700(.A(new_n650), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n879), .A2(new_n886), .A3(new_n887), .A4(new_n514), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n885), .A2(new_n888), .A3(new_n675), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n524), .B(new_n641), .C1(new_n635), .C2(new_n700), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n881), .A2(new_n882), .A3(new_n889), .A4(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n878), .A2(new_n891), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n712), .A2(new_n602), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n742), .A2(new_n744), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n893), .B1(new_n894), .B2(new_n707), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n734), .A2(new_n647), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n706), .B(KEYINPUT113), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT114), .B1(new_n710), .B2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT114), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n699), .A2(new_n900), .A3(new_n897), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n715), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n731), .A2(new_n896), .A3(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n895), .A2(KEYINPUT52), .A3(new_n777), .A4(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n713), .A2(new_n745), .A3(new_n903), .A4(new_n777), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT52), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT115), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n904), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  OR3_X1    g723(.A1(new_n905), .A2(new_n908), .A3(new_n906), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n892), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n904), .A2(new_n907), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n892), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g727(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n914));
  OAI22_X1  g728(.A1(new_n911), .A2(KEYINPUT53), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(KEYINPUT54), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n905), .B(KEYINPUT52), .ZN(new_n917));
  AOI22_X1  g731(.A1(new_n783), .A2(new_n789), .B1(new_n794), .B2(new_n796), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n890), .A2(new_n889), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n687), .A2(new_n466), .A3(new_n514), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n747), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n753), .B1(new_n921), .B2(new_n749), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n763), .A2(new_n880), .A3(new_n774), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n918), .A2(new_n919), .A3(new_n924), .A4(new_n877), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n914), .B1(new_n917), .B2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT117), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n913), .A2(KEYINPUT117), .A3(new_n914), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n892), .A2(new_n909), .A3(KEYINPUT53), .A4(new_n910), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n916), .B1(KEYINPUT54), .B2(new_n931), .ZN(new_n932));
  OAI22_X1  g746(.A1(new_n872), .A2(new_n932), .B1(G952), .B2(G953), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n851), .B(KEYINPUT49), .Z(new_n934));
  NOR4_X1   g748(.A1(new_n934), .A2(new_n765), .A3(new_n639), .A4(new_n852), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n799), .ZN(new_n936));
  OR3_X1    g750(.A1(new_n936), .A2(new_n731), .A3(new_n733), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n933), .A2(new_n937), .ZN(G75));
  AND2_X1   g752(.A1(new_n294), .A2(new_n296), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(new_n300), .ZN(new_n940));
  XOR2_X1   g754(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n931), .A2(G902), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(G210), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT56), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n355), .A2(G952), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n942), .A2(new_n945), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n948), .B1(new_n943), .B2(new_n188), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n946), .A2(new_n947), .A3(new_n949), .ZN(G51));
  NAND2_X1  g764(.A1(new_n943), .A2(new_n809), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT121), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n931), .B(KEYINPUT54), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n383), .B(KEYINPUT57), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n956), .B1(new_n381), .B2(new_n378), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n947), .B1(new_n953), .B2(new_n957), .ZN(G54));
  NAND3_X1  g772(.A1(new_n943), .A2(KEYINPUT58), .A3(G475), .ZN(new_n959));
  INV_X1    g773(.A(new_n683), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n959), .A2(new_n960), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n961), .A2(new_n962), .A3(new_n947), .ZN(G60));
  OR2_X1    g777(.A1(new_n665), .A2(new_n666), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n964), .A2(new_n659), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT122), .ZN(new_n966));
  NAND2_X1  g780(.A1(G478), .A2(G902), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT59), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n954), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n966), .B1(new_n932), .B2(new_n968), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n969), .A2(new_n947), .A3(new_n970), .ZN(G63));
  NAND2_X1  g785(.A1(G217), .A2(G902), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT60), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n914), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n975), .B1(new_n892), .B2(new_n912), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n930), .B1(new_n976), .B2(KEYINPUT117), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n926), .A2(new_n927), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n697), .B(new_n974), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n947), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n979), .A2(KEYINPUT61), .A3(new_n980), .ZN(new_n981));
  AOI211_X1 g795(.A(KEYINPUT123), .B(new_n631), .C1(new_n931), .C2(new_n974), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT123), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n974), .B1(new_n977), .B2(new_n978), .ZN(new_n984));
  INV_X1    g798(.A(new_n631), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NOR3_X1   g800(.A1(new_n981), .A2(new_n982), .A3(new_n986), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n979), .A2(new_n980), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n984), .A2(new_n985), .ZN(new_n989));
  AOI21_X1  g803(.A(KEYINPUT61), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(KEYINPUT124), .B1(new_n987), .B2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT124), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT61), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n979), .A2(new_n980), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n631), .B1(new_n931), .B2(new_n974), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n993), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(new_n986), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n995), .A2(new_n983), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n992), .B(new_n996), .C1(new_n999), .C2(new_n981), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n991), .A2(new_n1000), .ZN(G66));
  AOI21_X1  g815(.A(new_n355), .B1(new_n518), .B2(G224), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1002), .B1(new_n891), .B2(new_n355), .ZN(new_n1003));
  INV_X1    g817(.A(G898), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n939), .B1(new_n1004), .B2(G953), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1003), .B(new_n1005), .ZN(G69));
  NAND2_X1  g820(.A1(new_n441), .A2(new_n442), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n562), .B(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(G900), .B1(new_n1009), .B2(G227), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(G953), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1008), .A2(new_n355), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n895), .A2(new_n777), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1013), .A2(new_n736), .ZN(new_n1014));
  OR2_X1    g828(.A1(new_n1014), .A2(KEYINPUT62), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(KEYINPUT62), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n717), .B1(new_n669), .B2(new_n884), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n635), .A2(new_n1017), .A3(new_n793), .ZN(new_n1018));
  AND4_X1   g832(.A1(new_n818), .A2(new_n1015), .A3(new_n1016), .A4(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1012), .B1(new_n1019), .B2(new_n833), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n816), .A2(new_n896), .A3(new_n786), .ZN(new_n1021));
  AND4_X1   g835(.A1(new_n818), .A2(new_n1013), .A3(new_n918), .A4(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1022), .A2(new_n833), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1023), .A2(new_n355), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1020), .B1(new_n1024), .B2(new_n1009), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n355), .B1(G227), .B2(G900), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1026), .B(KEYINPUT125), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1011), .B1(new_n1025), .B2(new_n1027), .ZN(G72));
  NOR2_X1   g842(.A1(new_n572), .A2(new_n581), .ZN(new_n1029));
  XNOR2_X1  g843(.A(new_n1029), .B(KEYINPUT126), .ZN(new_n1030));
  INV_X1    g844(.A(new_n891), .ZN(new_n1031));
  AND3_X1   g845(.A1(new_n1019), .A2(new_n833), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g846(.A1(G472), .A2(G902), .ZN(new_n1033));
  XOR2_X1   g847(.A(new_n1033), .B(KEYINPUT63), .Z(new_n1034));
  INV_X1    g848(.A(new_n1034), .ZN(new_n1035));
  OAI211_X1 g849(.A(new_n568), .B(new_n1030), .C1(new_n1032), .C2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1034), .B1(new_n1023), .B2(new_n891), .ZN(new_n1037));
  NOR2_X1   g851(.A1(new_n1030), .A2(new_n568), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g853(.A(new_n592), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n1034), .B1(new_n1040), .B2(new_n721), .ZN(new_n1041));
  XNOR2_X1  g855(.A(new_n1041), .B(KEYINPUT127), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n947), .B1(new_n915), .B2(new_n1042), .ZN(new_n1043));
  AND3_X1   g857(.A1(new_n1036), .A2(new_n1039), .A3(new_n1043), .ZN(G57));
endmodule


