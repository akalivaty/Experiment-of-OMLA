

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U565 ( .A1(G2104), .A2(n560), .ZN(n898) );
  AND2_X1 U566 ( .A1(n560), .A2(G2104), .ZN(n901) );
  AND2_X1 U567 ( .A1(G2105), .A2(G2104), .ZN(n897) );
  NAND2_X1 U568 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X2 U569 ( .A1(n585), .A2(n584), .ZN(n982) );
  NOR2_X2 U570 ( .A1(n583), .A2(n582), .ZN(n585) );
  XNOR2_X2 U571 ( .A(n566), .B(KEYINPUT65), .ZN(G160) );
  NAND2_X1 U572 ( .A1(n690), .A2(n783), .ZN(n741) );
  NAND2_X1 U573 ( .A1(G160), .A2(G40), .ZN(n782) );
  NOR2_X2 U574 ( .A1(G2105), .A2(G2104), .ZN(n557) );
  AND2_X1 U575 ( .A1(n783), .A2(n690), .ZN(n721) );
  NOR2_X1 U576 ( .A1(n762), .A2(n988), .ZN(n763) );
  AND2_X1 U577 ( .A1(n779), .A2(n531), .ZN(n780) );
  XOR2_X1 U578 ( .A(n562), .B(KEYINPUT66), .Z(n530) );
  NAND2_X1 U579 ( .A1(n781), .A2(n780), .ZN(n815) );
  NOR2_X2 U580 ( .A1(n757), .A2(n756), .ZN(n772) );
  XOR2_X2 U581 ( .A(KEYINPUT17), .B(n557), .Z(n902) );
  OR2_X1 U582 ( .A1(n778), .A2(n777), .ZN(n531) );
  NOR2_X1 U583 ( .A1(n814), .A2(n821), .ZN(n532) );
  OR2_X1 U584 ( .A1(n750), .A2(n728), .ZN(n729) );
  XNOR2_X1 U585 ( .A(n730), .B(KEYINPUT30), .ZN(n731) );
  INV_X1 U586 ( .A(KEYINPUT99), .ZN(n739) );
  XOR2_X1 U587 ( .A(G543), .B(KEYINPUT0), .Z(n648) );
  XNOR2_X1 U588 ( .A(n595), .B(n594), .ZN(n694) );
  XNOR2_X1 U589 ( .A(KEYINPUT64), .B(n541), .ZN(n659) );
  NOR2_X1 U590 ( .A1(G651), .A2(G543), .ZN(n654) );
  NAND2_X1 U591 ( .A1(G89), .A2(n654), .ZN(n533) );
  XNOR2_X1 U592 ( .A(n533), .B(KEYINPUT76), .ZN(n534) );
  XNOR2_X1 U593 ( .A(KEYINPUT4), .B(n534), .ZN(n537) );
  INV_X1 U594 ( .A(G651), .ZN(n539) );
  NOR2_X1 U595 ( .A1(n648), .A2(n539), .ZN(n655) );
  NAND2_X1 U596 ( .A1(n655), .A2(G76), .ZN(n535) );
  XOR2_X1 U597 ( .A(KEYINPUT77), .B(n535), .Z(n536) );
  NAND2_X1 U598 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U599 ( .A(KEYINPUT5), .B(n538), .ZN(n547) );
  NOR2_X1 U600 ( .A1(G543), .A2(n539), .ZN(n540) );
  XOR2_X1 U601 ( .A(KEYINPUT1), .B(n540), .Z(n580) );
  NAND2_X1 U602 ( .A1(G63), .A2(n580), .ZN(n543) );
  NOR2_X1 U603 ( .A1(G651), .A2(n648), .ZN(n541) );
  NAND2_X1 U604 ( .A1(G51), .A2(n659), .ZN(n542) );
  NAND2_X1 U605 ( .A1(n543), .A2(n542), .ZN(n545) );
  XOR2_X1 U606 ( .A(KEYINPUT6), .B(KEYINPUT78), .Z(n544) );
  XNOR2_X1 U607 ( .A(n545), .B(n544), .ZN(n546) );
  NAND2_X1 U608 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U609 ( .A(KEYINPUT7), .B(n548), .ZN(G168) );
  XOR2_X1 U610 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U611 ( .A1(G64), .A2(n580), .ZN(n550) );
  NAND2_X1 U612 ( .A1(G52), .A2(n659), .ZN(n549) );
  NAND2_X1 U613 ( .A1(n550), .A2(n549), .ZN(n556) );
  NAND2_X1 U614 ( .A1(G90), .A2(n654), .ZN(n552) );
  NAND2_X1 U615 ( .A1(G77), .A2(n655), .ZN(n551) );
  NAND2_X1 U616 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U617 ( .A(KEYINPUT9), .B(n553), .Z(n554) );
  XNOR2_X1 U618 ( .A(KEYINPUT68), .B(n554), .ZN(n555) );
  NOR2_X1 U619 ( .A1(n556), .A2(n555), .ZN(G171) );
  AND2_X1 U620 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U621 ( .A(G57), .ZN(G237) );
  INV_X1 U622 ( .A(G132), .ZN(G219) );
  NAND2_X1 U623 ( .A1(G137), .A2(n902), .ZN(n559) );
  INV_X1 U624 ( .A(G2105), .ZN(n560) );
  NAND2_X1 U625 ( .A1(G125), .A2(n898), .ZN(n558) );
  AND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n565) );
  NAND2_X1 U627 ( .A1(G101), .A2(n901), .ZN(n561) );
  XNOR2_X1 U628 ( .A(KEYINPUT23), .B(n561), .ZN(n563) );
  NAND2_X1 U629 ( .A1(G113), .A2(n897), .ZN(n562) );
  NOR2_X1 U630 ( .A1(n563), .A2(n530), .ZN(n564) );
  NAND2_X1 U631 ( .A1(G102), .A2(n901), .ZN(n568) );
  NAND2_X1 U632 ( .A1(G138), .A2(n902), .ZN(n567) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n572) );
  NAND2_X1 U634 ( .A1(G114), .A2(n897), .ZN(n570) );
  NAND2_X1 U635 ( .A1(G126), .A2(n898), .ZN(n569) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U637 ( .A1(n572), .A2(n571), .ZN(G164) );
  NAND2_X1 U638 ( .A1(G7), .A2(G661), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U640 ( .A(G223), .ZN(n844) );
  NAND2_X1 U641 ( .A1(n844), .A2(G567), .ZN(n574) );
  XOR2_X1 U642 ( .A(KEYINPUT11), .B(n574), .Z(G234) );
  NAND2_X1 U643 ( .A1(n654), .A2(G81), .ZN(n575) );
  XNOR2_X1 U644 ( .A(n575), .B(KEYINPUT12), .ZN(n577) );
  NAND2_X1 U645 ( .A1(G68), .A2(n655), .ZN(n576) );
  NAND2_X1 U646 ( .A1(n577), .A2(n576), .ZN(n579) );
  XOR2_X1 U647 ( .A(KEYINPUT13), .B(KEYINPUT72), .Z(n578) );
  XNOR2_X1 U648 ( .A(n579), .B(n578), .ZN(n583) );
  NAND2_X1 U649 ( .A1(n580), .A2(G56), .ZN(n581) );
  XOR2_X1 U650 ( .A(KEYINPUT14), .B(n581), .Z(n582) );
  NAND2_X1 U651 ( .A1(G43), .A2(n659), .ZN(n584) );
  INV_X1 U652 ( .A(G860), .ZN(n625) );
  OR2_X1 U653 ( .A1(n982), .A2(n625), .ZN(G153) );
  INV_X1 U654 ( .A(G868), .ZN(n674) );
  NAND2_X1 U655 ( .A1(n659), .A2(G54), .ZN(n586) );
  XNOR2_X1 U656 ( .A(n586), .B(KEYINPUT74), .ZN(n593) );
  NAND2_X1 U657 ( .A1(G79), .A2(n655), .ZN(n588) );
  NAND2_X1 U658 ( .A1(G66), .A2(n580), .ZN(n587) );
  NAND2_X1 U659 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U660 ( .A1(G92), .A2(n654), .ZN(n589) );
  XNOR2_X1 U661 ( .A(KEYINPUT73), .B(n589), .ZN(n590) );
  NOR2_X1 U662 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U663 ( .A1(n593), .A2(n592), .ZN(n595) );
  INV_X1 U664 ( .A(KEYINPUT15), .ZN(n594) );
  INV_X1 U665 ( .A(n694), .ZN(n989) );
  NAND2_X1 U666 ( .A1(n674), .A2(n989), .ZN(n597) );
  NAND2_X1 U667 ( .A1(G171), .A2(G868), .ZN(n596) );
  NAND2_X1 U668 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U669 ( .A(n598), .B(KEYINPUT75), .ZN(G284) );
  NAND2_X1 U670 ( .A1(n659), .A2(G53), .ZN(n599) );
  XNOR2_X1 U671 ( .A(n599), .B(KEYINPUT70), .ZN(n606) );
  NAND2_X1 U672 ( .A1(G91), .A2(n654), .ZN(n601) );
  NAND2_X1 U673 ( .A1(G78), .A2(n655), .ZN(n600) );
  NAND2_X1 U674 ( .A1(n601), .A2(n600), .ZN(n604) );
  NAND2_X1 U675 ( .A1(G65), .A2(n580), .ZN(n602) );
  XNOR2_X1 U676 ( .A(KEYINPUT69), .B(n602), .ZN(n603) );
  NOR2_X1 U677 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U678 ( .A1(n606), .A2(n605), .ZN(G299) );
  NOR2_X1 U679 ( .A1(G286), .A2(n674), .ZN(n608) );
  NOR2_X1 U680 ( .A1(G868), .A2(G299), .ZN(n607) );
  NOR2_X1 U681 ( .A1(n608), .A2(n607), .ZN(G297) );
  NAND2_X1 U682 ( .A1(n625), .A2(G559), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n609), .A2(n989), .ZN(n610) );
  XNOR2_X1 U684 ( .A(n610), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U685 ( .A1(G868), .A2(n982), .ZN(n613) );
  NAND2_X1 U686 ( .A1(G868), .A2(n989), .ZN(n611) );
  NOR2_X1 U687 ( .A1(G559), .A2(n611), .ZN(n612) );
  NOR2_X1 U688 ( .A1(n613), .A2(n612), .ZN(G282) );
  NAND2_X1 U689 ( .A1(G111), .A2(n897), .ZN(n620) );
  NAND2_X1 U690 ( .A1(G99), .A2(n901), .ZN(n615) );
  NAND2_X1 U691 ( .A1(G135), .A2(n902), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U693 ( .A1(n898), .A2(G123), .ZN(n616) );
  XOR2_X1 U694 ( .A(KEYINPUT18), .B(n616), .Z(n617) );
  NOR2_X1 U695 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U696 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U697 ( .A(n621), .B(KEYINPUT79), .ZN(n953) );
  XNOR2_X1 U698 ( .A(G2096), .B(n953), .ZN(n623) );
  INV_X1 U699 ( .A(G2100), .ZN(n622) );
  NAND2_X1 U700 ( .A1(n623), .A2(n622), .ZN(G156) );
  NAND2_X1 U701 ( .A1(G559), .A2(n989), .ZN(n624) );
  XOR2_X1 U702 ( .A(n982), .B(n624), .Z(n671) );
  NAND2_X1 U703 ( .A1(n625), .A2(n671), .ZN(n632) );
  NAND2_X1 U704 ( .A1(G93), .A2(n654), .ZN(n627) );
  NAND2_X1 U705 ( .A1(G80), .A2(n655), .ZN(n626) );
  NAND2_X1 U706 ( .A1(n627), .A2(n626), .ZN(n631) );
  NAND2_X1 U707 ( .A1(G67), .A2(n580), .ZN(n629) );
  NAND2_X1 U708 ( .A1(G55), .A2(n659), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U710 ( .A1(n631), .A2(n630), .ZN(n673) );
  XOR2_X1 U711 ( .A(n632), .B(n673), .Z(G145) );
  XOR2_X1 U712 ( .A(KEYINPUT80), .B(KEYINPUT2), .Z(n634) );
  NAND2_X1 U713 ( .A1(G73), .A2(n655), .ZN(n633) );
  XNOR2_X1 U714 ( .A(n634), .B(n633), .ZN(n638) );
  NAND2_X1 U715 ( .A1(G86), .A2(n654), .ZN(n636) );
  NAND2_X1 U716 ( .A1(G61), .A2(n580), .ZN(n635) );
  NAND2_X1 U717 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U718 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U719 ( .A1(G48), .A2(n659), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n640), .A2(n639), .ZN(G305) );
  NAND2_X1 U721 ( .A1(G60), .A2(n580), .ZN(n642) );
  NAND2_X1 U722 ( .A1(G47), .A2(n659), .ZN(n641) );
  NAND2_X1 U723 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U724 ( .A(KEYINPUT67), .B(n643), .ZN(n647) );
  NAND2_X1 U725 ( .A1(G85), .A2(n654), .ZN(n645) );
  NAND2_X1 U726 ( .A1(G72), .A2(n655), .ZN(n644) );
  AND2_X1 U727 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U728 ( .A1(n647), .A2(n646), .ZN(G290) );
  NAND2_X1 U729 ( .A1(n648), .A2(G87), .ZN(n650) );
  NAND2_X1 U730 ( .A1(G49), .A2(n659), .ZN(n649) );
  NAND2_X1 U731 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U732 ( .A1(n580), .A2(n651), .ZN(n653) );
  NAND2_X1 U733 ( .A1(G651), .A2(G74), .ZN(n652) );
  NAND2_X1 U734 ( .A1(n653), .A2(n652), .ZN(G288) );
  NAND2_X1 U735 ( .A1(G88), .A2(n654), .ZN(n657) );
  NAND2_X1 U736 ( .A1(G75), .A2(n655), .ZN(n656) );
  NAND2_X1 U737 ( .A1(n657), .A2(n656), .ZN(n663) );
  NAND2_X1 U738 ( .A1(G62), .A2(n580), .ZN(n658) );
  XOR2_X1 U739 ( .A(KEYINPUT81), .B(n658), .Z(n661) );
  NAND2_X1 U740 ( .A1(G50), .A2(n659), .ZN(n660) );
  NAND2_X1 U741 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U742 ( .A1(n663), .A2(n662), .ZN(G166) );
  INV_X1 U743 ( .A(G299), .ZN(n711) );
  XNOR2_X1 U744 ( .A(n711), .B(G305), .ZN(n664) );
  XNOR2_X1 U745 ( .A(n664), .B(G290), .ZN(n668) );
  XNOR2_X1 U746 ( .A(KEYINPUT83), .B(KEYINPUT82), .ZN(n666) );
  XNOR2_X1 U747 ( .A(G288), .B(KEYINPUT19), .ZN(n665) );
  XNOR2_X1 U748 ( .A(n666), .B(n665), .ZN(n667) );
  XOR2_X1 U749 ( .A(n668), .B(n667), .Z(n670) );
  XNOR2_X1 U750 ( .A(G166), .B(n673), .ZN(n669) );
  XNOR2_X1 U751 ( .A(n670), .B(n669), .ZN(n913) );
  XOR2_X1 U752 ( .A(n913), .B(n671), .Z(n672) );
  NOR2_X1 U753 ( .A1(n674), .A2(n672), .ZN(n676) );
  AND2_X1 U754 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U755 ( .A1(n676), .A2(n675), .ZN(G295) );
  NAND2_X1 U756 ( .A1(G2078), .A2(G2084), .ZN(n677) );
  XOR2_X1 U757 ( .A(KEYINPUT20), .B(n677), .Z(n678) );
  NAND2_X1 U758 ( .A1(G2090), .A2(n678), .ZN(n679) );
  XNOR2_X1 U759 ( .A(KEYINPUT21), .B(n679), .ZN(n680) );
  NAND2_X1 U760 ( .A1(n680), .A2(G2072), .ZN(n681) );
  XNOR2_X1 U761 ( .A(KEYINPUT84), .B(n681), .ZN(G158) );
  XNOR2_X1 U762 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U763 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  NOR2_X1 U764 ( .A1(G219), .A2(G220), .ZN(n682) );
  XOR2_X1 U765 ( .A(KEYINPUT22), .B(n682), .Z(n683) );
  NOR2_X1 U766 ( .A1(G218), .A2(n683), .ZN(n684) );
  NAND2_X1 U767 ( .A1(G96), .A2(n684), .ZN(n848) );
  NAND2_X1 U768 ( .A1(n848), .A2(G2106), .ZN(n688) );
  NAND2_X1 U769 ( .A1(G69), .A2(G120), .ZN(n685) );
  NOR2_X1 U770 ( .A1(G237), .A2(n685), .ZN(n686) );
  NAND2_X1 U771 ( .A1(G108), .A2(n686), .ZN(n849) );
  NAND2_X1 U772 ( .A1(n849), .A2(G567), .ZN(n687) );
  NAND2_X1 U773 ( .A1(n688), .A2(n687), .ZN(n871) );
  NAND2_X1 U774 ( .A1(G661), .A2(G483), .ZN(n689) );
  NOR2_X1 U775 ( .A1(n871), .A2(n689), .ZN(n847) );
  NAND2_X1 U776 ( .A1(n847), .A2(G36), .ZN(G176) );
  XNOR2_X1 U777 ( .A(KEYINPUT85), .B(G166), .ZN(G303) );
  XNOR2_X1 U778 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n833) );
  INV_X1 U779 ( .A(n782), .ZN(n690) );
  NOR2_X1 U780 ( .A1(G164), .A2(G1384), .ZN(n783) );
  NOR2_X1 U781 ( .A1(G2067), .A2(n741), .ZN(n692) );
  NOR2_X1 U782 ( .A1(n721), .A2(G1348), .ZN(n691) );
  NOR2_X1 U783 ( .A1(n692), .A2(n691), .ZN(n693) );
  OR2_X1 U784 ( .A1(n693), .A2(n694), .ZN(n704) );
  NAND2_X1 U785 ( .A1(n694), .A2(n693), .ZN(n702) );
  NAND2_X1 U786 ( .A1(n783), .A2(G1996), .ZN(n695) );
  NOR2_X1 U787 ( .A1(n695), .A2(n782), .ZN(n696) );
  XNOR2_X1 U788 ( .A(n696), .B(KEYINPUT26), .ZN(n700) );
  NAND2_X1 U789 ( .A1(n741), .A2(G1341), .ZN(n698) );
  INV_X1 U790 ( .A(n982), .ZN(n697) );
  NAND2_X1 U791 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U792 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U793 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U794 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U795 ( .A(n705), .B(KEYINPUT97), .ZN(n710) );
  NAND2_X1 U796 ( .A1(n721), .A2(G2072), .ZN(n706) );
  XNOR2_X1 U797 ( .A(n706), .B(KEYINPUT27), .ZN(n708) );
  AND2_X1 U798 ( .A1(G1956), .A2(n741), .ZN(n707) );
  NOR2_X1 U799 ( .A1(n708), .A2(n707), .ZN(n712) );
  NAND2_X1 U800 ( .A1(n712), .A2(n711), .ZN(n709) );
  NAND2_X1 U801 ( .A1(n710), .A2(n709), .ZN(n716) );
  NOR2_X1 U802 ( .A1(n712), .A2(n711), .ZN(n714) );
  XOR2_X1 U803 ( .A(KEYINPUT28), .B(KEYINPUT96), .Z(n713) );
  XNOR2_X1 U804 ( .A(n714), .B(n713), .ZN(n715) );
  NAND2_X1 U805 ( .A1(n716), .A2(n715), .ZN(n718) );
  XOR2_X1 U806 ( .A(KEYINPUT29), .B(KEYINPUT98), .Z(n717) );
  XNOR2_X1 U807 ( .A(n718), .B(n717), .ZN(n727) );
  XOR2_X1 U808 ( .A(G2078), .B(KEYINPUT25), .Z(n719) );
  XNOR2_X1 U809 ( .A(KEYINPUT93), .B(n719), .ZN(n928) );
  NAND2_X1 U810 ( .A1(n721), .A2(n928), .ZN(n720) );
  XNOR2_X1 U811 ( .A(KEYINPUT94), .B(n720), .ZN(n724) );
  NOR2_X1 U812 ( .A1(n721), .A2(G1961), .ZN(n722) );
  XOR2_X1 U813 ( .A(KEYINPUT92), .B(n722), .Z(n723) );
  NAND2_X1 U814 ( .A1(n724), .A2(n723), .ZN(n732) );
  AND2_X1 U815 ( .A1(n732), .A2(G171), .ZN(n725) );
  XNOR2_X1 U816 ( .A(KEYINPUT95), .B(n725), .ZN(n726) );
  NAND2_X1 U817 ( .A1(n727), .A2(n726), .ZN(n738) );
  NAND2_X1 U818 ( .A1(G8), .A2(n741), .ZN(n778) );
  NOR2_X1 U819 ( .A1(n778), .A2(G1966), .ZN(n755) );
  NOR2_X1 U820 ( .A1(G2084), .A2(n741), .ZN(n750) );
  INV_X1 U821 ( .A(G8), .ZN(n728) );
  OR2_X1 U822 ( .A1(n755), .A2(n729), .ZN(n730) );
  NOR2_X1 U823 ( .A1(n731), .A2(G168), .ZN(n734) );
  NOR2_X1 U824 ( .A1(G171), .A2(n732), .ZN(n733) );
  NOR2_X1 U825 ( .A1(n734), .A2(n733), .ZN(n736) );
  INV_X1 U826 ( .A(KEYINPUT31), .ZN(n735) );
  XNOR2_X1 U827 ( .A(n736), .B(n735), .ZN(n737) );
  NAND2_X1 U828 ( .A1(n738), .A2(n737), .ZN(n752) );
  NAND2_X1 U829 ( .A1(n752), .A2(G286), .ZN(n740) );
  XNOR2_X1 U830 ( .A(n740), .B(n739), .ZN(n747) );
  NOR2_X1 U831 ( .A1(G1971), .A2(n778), .ZN(n743) );
  NOR2_X1 U832 ( .A1(G2090), .A2(n741), .ZN(n742) );
  NOR2_X1 U833 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U834 ( .A1(n744), .A2(G303), .ZN(n745) );
  XNOR2_X1 U835 ( .A(KEYINPUT100), .B(n745), .ZN(n746) );
  NAND2_X1 U836 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U837 ( .A1(n748), .A2(G8), .ZN(n749) );
  XOR2_X1 U838 ( .A(KEYINPUT32), .B(n749), .Z(n757) );
  NAND2_X1 U839 ( .A1(G8), .A2(n750), .ZN(n751) );
  XOR2_X1 U840 ( .A(KEYINPUT91), .B(n751), .Z(n753) );
  NAND2_X1 U841 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U842 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n981) );
  NOR2_X1 U844 ( .A1(G1971), .A2(G303), .ZN(n758) );
  NOR2_X1 U845 ( .A1(n981), .A2(n758), .ZN(n759) );
  XNOR2_X1 U846 ( .A(n759), .B(KEYINPUT101), .ZN(n760) );
  NOR2_X1 U847 ( .A1(n772), .A2(n760), .ZN(n762) );
  NAND2_X1 U848 ( .A1(G288), .A2(G1976), .ZN(n761) );
  XOR2_X1 U849 ( .A(KEYINPUT102), .B(n761), .Z(n988) );
  XNOR2_X1 U850 ( .A(n763), .B(KEYINPUT103), .ZN(n764) );
  NOR2_X1 U851 ( .A1(n764), .A2(n778), .ZN(n765) );
  NOR2_X1 U852 ( .A1(KEYINPUT33), .A2(n765), .ZN(n768) );
  NAND2_X1 U853 ( .A1(n981), .A2(KEYINPUT33), .ZN(n766) );
  NOR2_X1 U854 ( .A1(n766), .A2(n778), .ZN(n767) );
  NOR2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U856 ( .A(G1981), .B(G305), .Z(n973) );
  NAND2_X1 U857 ( .A1(n769), .A2(n973), .ZN(n781) );
  NOR2_X1 U858 ( .A1(G2090), .A2(G303), .ZN(n770) );
  XNOR2_X1 U859 ( .A(n770), .B(KEYINPUT104), .ZN(n771) );
  NAND2_X1 U860 ( .A1(n771), .A2(G8), .ZN(n774) );
  INV_X1 U861 ( .A(n772), .ZN(n773) );
  NAND2_X1 U862 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U863 ( .A1(n775), .A2(n778), .ZN(n779) );
  NOR2_X1 U864 ( .A1(G1981), .A2(G305), .ZN(n776) );
  XOR2_X1 U865 ( .A(n776), .B(KEYINPUT24), .Z(n777) );
  NOR2_X1 U866 ( .A1(n783), .A2(n782), .ZN(n784) );
  XOR2_X1 U867 ( .A(KEYINPUT86), .B(n784), .Z(n828) );
  XOR2_X1 U868 ( .A(G2067), .B(KEYINPUT37), .Z(n816) );
  NAND2_X1 U869 ( .A1(G104), .A2(n901), .ZN(n786) );
  NAND2_X1 U870 ( .A1(G140), .A2(n902), .ZN(n785) );
  NAND2_X1 U871 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U872 ( .A(KEYINPUT34), .B(n787), .ZN(n792) );
  NAND2_X1 U873 ( .A1(G116), .A2(n897), .ZN(n789) );
  NAND2_X1 U874 ( .A1(G128), .A2(n898), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U876 ( .A(n790), .B(KEYINPUT35), .Z(n791) );
  NOR2_X1 U877 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U878 ( .A(KEYINPUT87), .B(n793), .Z(n795) );
  XOR2_X1 U879 ( .A(KEYINPUT88), .B(KEYINPUT36), .Z(n794) );
  XNOR2_X1 U880 ( .A(n795), .B(n794), .ZN(n896) );
  NAND2_X1 U881 ( .A1(n816), .A2(n896), .ZN(n796) );
  XNOR2_X1 U882 ( .A(KEYINPUT89), .B(n796), .ZN(n966) );
  XNOR2_X1 U883 ( .A(G1986), .B(G290), .ZN(n991) );
  NOR2_X1 U884 ( .A1(n966), .A2(n991), .ZN(n797) );
  NOR2_X1 U885 ( .A1(n828), .A2(n797), .ZN(n814) );
  NAND2_X1 U886 ( .A1(G95), .A2(n901), .ZN(n799) );
  NAND2_X1 U887 ( .A1(G131), .A2(n902), .ZN(n798) );
  NAND2_X1 U888 ( .A1(n799), .A2(n798), .ZN(n803) );
  NAND2_X1 U889 ( .A1(G107), .A2(n897), .ZN(n801) );
  NAND2_X1 U890 ( .A1(G119), .A2(n898), .ZN(n800) );
  NAND2_X1 U891 ( .A1(n801), .A2(n800), .ZN(n802) );
  NOR2_X1 U892 ( .A1(n803), .A2(n802), .ZN(n880) );
  INV_X1 U893 ( .A(G1991), .ZN(n818) );
  NOR2_X1 U894 ( .A1(n880), .A2(n818), .ZN(n813) );
  XOR2_X1 U895 ( .A(KEYINPUT90), .B(KEYINPUT38), .Z(n805) );
  NAND2_X1 U896 ( .A1(G105), .A2(n901), .ZN(n804) );
  XNOR2_X1 U897 ( .A(n805), .B(n804), .ZN(n809) );
  NAND2_X1 U898 ( .A1(G141), .A2(n902), .ZN(n807) );
  NAND2_X1 U899 ( .A1(G129), .A2(n898), .ZN(n806) );
  NAND2_X1 U900 ( .A1(n807), .A2(n806), .ZN(n808) );
  NOR2_X1 U901 ( .A1(n809), .A2(n808), .ZN(n811) );
  NAND2_X1 U902 ( .A1(n897), .A2(G117), .ZN(n810) );
  NAND2_X1 U903 ( .A1(n811), .A2(n810), .ZN(n890) );
  AND2_X1 U904 ( .A1(n890), .A2(G1996), .ZN(n812) );
  NOR2_X1 U905 ( .A1(n813), .A2(n812), .ZN(n960) );
  NOR2_X1 U906 ( .A1(n960), .A2(n828), .ZN(n821) );
  NAND2_X1 U907 ( .A1(n815), .A2(n532), .ZN(n831) );
  NOR2_X1 U908 ( .A1(n816), .A2(n896), .ZN(n817) );
  XNOR2_X1 U909 ( .A(KEYINPUT106), .B(n817), .ZN(n962) );
  NOR2_X1 U910 ( .A1(G1996), .A2(n890), .ZN(n947) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n819) );
  AND2_X1 U912 ( .A1(n818), .A2(n880), .ZN(n954) );
  NOR2_X1 U913 ( .A1(n819), .A2(n954), .ZN(n820) );
  NOR2_X1 U914 ( .A1(n821), .A2(n820), .ZN(n822) );
  NOR2_X1 U915 ( .A1(n947), .A2(n822), .ZN(n823) );
  XNOR2_X1 U916 ( .A(n823), .B(KEYINPUT39), .ZN(n824) );
  XNOR2_X1 U917 ( .A(n824), .B(KEYINPUT105), .ZN(n825) );
  NOR2_X1 U918 ( .A1(n966), .A2(n825), .ZN(n826) );
  NOR2_X1 U919 ( .A1(n962), .A2(n826), .ZN(n827) );
  NOR2_X1 U920 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U921 ( .A(n829), .B(KEYINPUT107), .ZN(n830) );
  NAND2_X1 U922 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U923 ( .A(n833), .B(n832), .ZN(G329) );
  XOR2_X1 U924 ( .A(G2454), .B(G2430), .Z(n835) );
  XNOR2_X1 U925 ( .A(G2451), .B(G2446), .ZN(n834) );
  XNOR2_X1 U926 ( .A(n835), .B(n834), .ZN(n842) );
  XOR2_X1 U927 ( .A(G2443), .B(G2427), .Z(n837) );
  XNOR2_X1 U928 ( .A(G2438), .B(KEYINPUT109), .ZN(n836) );
  XNOR2_X1 U929 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U930 ( .A(n838), .B(G2435), .Z(n840) );
  XNOR2_X1 U931 ( .A(G1348), .B(G1341), .ZN(n839) );
  XNOR2_X1 U932 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U933 ( .A(n842), .B(n841), .ZN(n843) );
  NAND2_X1 U934 ( .A1(n843), .A2(G14), .ZN(n920) );
  XOR2_X1 U935 ( .A(KEYINPUT110), .B(n920), .Z(G401) );
  NAND2_X1 U936 ( .A1(G2106), .A2(n844), .ZN(G217) );
  AND2_X1 U937 ( .A1(G15), .A2(G2), .ZN(n845) );
  NAND2_X1 U938 ( .A1(G661), .A2(n845), .ZN(G259) );
  NAND2_X1 U939 ( .A1(G3), .A2(G1), .ZN(n846) );
  NAND2_X1 U940 ( .A1(n847), .A2(n846), .ZN(G188) );
  INV_X1 U942 ( .A(G120), .ZN(G236) );
  INV_X1 U943 ( .A(G96), .ZN(G221) );
  INV_X1 U944 ( .A(G69), .ZN(G235) );
  NOR2_X1 U945 ( .A1(n849), .A2(n848), .ZN(G325) );
  INV_X1 U946 ( .A(G325), .ZN(G261) );
  XOR2_X1 U947 ( .A(KEYINPUT113), .B(G1986), .Z(n851) );
  XNOR2_X1 U948 ( .A(G1961), .B(G1976), .ZN(n850) );
  XNOR2_X1 U949 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U950 ( .A(n852), .B(KEYINPUT41), .Z(n854) );
  XNOR2_X1 U951 ( .A(G1996), .B(G1991), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U953 ( .A(G1981), .B(G1971), .Z(n856) );
  XNOR2_X1 U954 ( .A(G1966), .B(G1956), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U956 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U957 ( .A(KEYINPUT114), .B(G2474), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n860), .B(n859), .ZN(G229) );
  XOR2_X1 U959 ( .A(KEYINPUT112), .B(G2096), .Z(n862) );
  XNOR2_X1 U960 ( .A(KEYINPUT43), .B(G2678), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U962 ( .A(G2100), .B(G2090), .Z(n864) );
  XNOR2_X1 U963 ( .A(G2072), .B(G2067), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U965 ( .A(n866), .B(n865), .Z(n868) );
  XNOR2_X1 U966 ( .A(KEYINPUT42), .B(KEYINPUT111), .ZN(n867) );
  XNOR2_X1 U967 ( .A(n868), .B(n867), .ZN(n870) );
  XOR2_X1 U968 ( .A(G2078), .B(G2084), .Z(n869) );
  XNOR2_X1 U969 ( .A(n870), .B(n869), .ZN(G227) );
  INV_X1 U970 ( .A(n871), .ZN(G319) );
  NAND2_X1 U971 ( .A1(G100), .A2(n901), .ZN(n873) );
  NAND2_X1 U972 ( .A1(G112), .A2(n897), .ZN(n872) );
  NAND2_X1 U973 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U974 ( .A(n874), .B(KEYINPUT115), .ZN(n876) );
  NAND2_X1 U975 ( .A1(G136), .A2(n902), .ZN(n875) );
  NAND2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n879) );
  NAND2_X1 U977 ( .A1(n898), .A2(G124), .ZN(n877) );
  XOR2_X1 U978 ( .A(KEYINPUT44), .B(n877), .Z(n878) );
  NOR2_X1 U979 ( .A1(n879), .A2(n878), .ZN(G162) );
  XOR2_X1 U980 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n882) );
  XNOR2_X1 U981 ( .A(n880), .B(n953), .ZN(n881) );
  XNOR2_X1 U982 ( .A(n882), .B(n881), .ZN(n894) );
  NAND2_X1 U983 ( .A1(G103), .A2(n901), .ZN(n884) );
  NAND2_X1 U984 ( .A1(G139), .A2(n902), .ZN(n883) );
  NAND2_X1 U985 ( .A1(n884), .A2(n883), .ZN(n889) );
  NAND2_X1 U986 ( .A1(G115), .A2(n897), .ZN(n886) );
  NAND2_X1 U987 ( .A1(G127), .A2(n898), .ZN(n885) );
  NAND2_X1 U988 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U989 ( .A(KEYINPUT47), .B(n887), .Z(n888) );
  NOR2_X1 U990 ( .A1(n889), .A2(n888), .ZN(n949) );
  XOR2_X1 U991 ( .A(n949), .B(G162), .Z(n892) );
  XOR2_X1 U992 ( .A(n890), .B(G164), .Z(n891) );
  XNOR2_X1 U993 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U994 ( .A(n894), .B(n893), .Z(n895) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n911) );
  NAND2_X1 U996 ( .A1(G118), .A2(n897), .ZN(n900) );
  NAND2_X1 U997 ( .A1(G130), .A2(n898), .ZN(n899) );
  NAND2_X1 U998 ( .A1(n900), .A2(n899), .ZN(n908) );
  NAND2_X1 U999 ( .A1(G106), .A2(n901), .ZN(n904) );
  NAND2_X1 U1000 ( .A1(G142), .A2(n902), .ZN(n903) );
  NAND2_X1 U1001 ( .A1(n904), .A2(n903), .ZN(n905) );
  XOR2_X1 U1002 ( .A(KEYINPUT45), .B(n905), .Z(n906) );
  XNOR2_X1 U1003 ( .A(KEYINPUT116), .B(n906), .ZN(n907) );
  NOR2_X1 U1004 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1005 ( .A(G160), .B(n909), .ZN(n910) );
  XNOR2_X1 U1006 ( .A(n911), .B(n910), .ZN(n912) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n912), .ZN(G395) );
  XNOR2_X1 U1008 ( .A(n913), .B(KEYINPUT117), .ZN(n915) );
  XNOR2_X1 U1009 ( .A(n982), .B(G171), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(n915), .B(n914), .ZN(n917) );
  XNOR2_X1 U1011 ( .A(G286), .B(n989), .ZN(n916) );
  XNOR2_X1 U1012 ( .A(n917), .B(n916), .ZN(n918) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n918), .ZN(G397) );
  NOR2_X1 U1014 ( .A1(G229), .A2(G227), .ZN(n919) );
  XOR2_X1 U1015 ( .A(KEYINPUT49), .B(n919), .Z(n923) );
  NAND2_X1 U1016 ( .A1(G319), .A2(n920), .ZN(n921) );
  XOR2_X1 U1017 ( .A(KEYINPUT118), .B(n921), .Z(n922) );
  NAND2_X1 U1018 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1019 ( .A(KEYINPUT119), .B(n924), .ZN(n926) );
  NOR2_X1 U1020 ( .A1(G395), .A2(G397), .ZN(n925) );
  NAND2_X1 U1021 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1022 ( .A(KEYINPUT120), .B(n927), .Z(G308) );
  INV_X1 U1023 ( .A(G308), .ZN(G225) );
  INV_X1 U1024 ( .A(G171), .ZN(G301) );
  INV_X1 U1025 ( .A(G108), .ZN(G238) );
  INV_X1 U1026 ( .A(KEYINPUT55), .ZN(n968) );
  XNOR2_X1 U1027 ( .A(G2090), .B(G35), .ZN(n942) );
  XNOR2_X1 U1028 ( .A(G27), .B(n928), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(G1996), .B(G32), .ZN(n930) );
  XNOR2_X1 U1030 ( .A(G26), .B(G2067), .ZN(n929) );
  NOR2_X1 U1031 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1032 ( .A1(n932), .A2(n931), .ZN(n934) );
  XNOR2_X1 U1033 ( .A(G33), .B(G2072), .ZN(n933) );
  NOR2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1035 ( .A(KEYINPUT122), .B(n935), .ZN(n936) );
  NAND2_X1 U1036 ( .A1(n936), .A2(G28), .ZN(n939) );
  XOR2_X1 U1037 ( .A(G25), .B(G1991), .Z(n937) );
  XNOR2_X1 U1038 ( .A(KEYINPUT121), .B(n937), .ZN(n938) );
  NOR2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1040 ( .A(KEYINPUT53), .B(n940), .ZN(n941) );
  NOR2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n945) );
  XOR2_X1 U1042 ( .A(G2084), .B(KEYINPUT54), .Z(n943) );
  XNOR2_X1 U1043 ( .A(G34), .B(n943), .ZN(n944) );
  NAND2_X1 U1044 ( .A1(n945), .A2(n944), .ZN(n1023) );
  OR2_X1 U1045 ( .A1(n968), .A2(n1023), .ZN(n972) );
  XOR2_X1 U1046 ( .A(G2090), .B(G162), .Z(n946) );
  NOR2_X1 U1047 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1048 ( .A(KEYINPUT51), .B(n948), .Z(n964) );
  XOR2_X1 U1049 ( .A(G2072), .B(n949), .Z(n951) );
  XOR2_X1 U1050 ( .A(G164), .B(G2078), .Z(n950) );
  NOR2_X1 U1051 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1052 ( .A(KEYINPUT50), .B(n952), .ZN(n956) );
  NOR2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1054 ( .A1(n956), .A2(n955), .ZN(n958) );
  XOR2_X1 U1055 ( .A(G160), .B(G2084), .Z(n957) );
  NOR2_X1 U1056 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  NOR2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(n967), .B(KEYINPUT52), .ZN(n969) );
  NAND2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1063 ( .A1(G29), .A2(n970), .ZN(n971) );
  NAND2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n1030) );
  XOR2_X1 U1065 ( .A(G16), .B(KEYINPUT56), .Z(n997) );
  XNOR2_X1 U1066 ( .A(G1966), .B(G168), .ZN(n974) );
  NAND2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(n975), .B(KEYINPUT123), .ZN(n976) );
  XOR2_X1 U1069 ( .A(KEYINPUT57), .B(n976), .Z(n979) );
  XOR2_X1 U1070 ( .A(G1971), .B(G303), .Z(n977) );
  XNOR2_X1 U1071 ( .A(KEYINPUT124), .B(n977), .ZN(n978) );
  NAND2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n995) );
  XOR2_X1 U1073 ( .A(G1961), .B(G171), .Z(n980) );
  NOR2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n986) );
  XNOR2_X1 U1075 ( .A(G299), .B(G1956), .ZN(n984) );
  XNOR2_X1 U1076 ( .A(n982), .B(G1341), .ZN(n983) );
  NOR2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  NOR2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n993) );
  XOR2_X1 U1080 ( .A(G1348), .B(n989), .Z(n990) );
  NOR2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1083 ( .A1(n995), .A2(n994), .ZN(n996) );
  NOR2_X1 U1084 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1085 ( .A(KEYINPUT125), .B(n998), .ZN(n1028) );
  XNOR2_X1 U1086 ( .A(G1961), .B(KEYINPUT126), .ZN(n999) );
  XNOR2_X1 U1087 ( .A(n999), .B(G5), .ZN(n1006) );
  XNOR2_X1 U1088 ( .A(G1971), .B(G22), .ZN(n1001) );
  XNOR2_X1 U1089 ( .A(G23), .B(G1976), .ZN(n1000) );
  NOR2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1003) );
  XOR2_X1 U1091 ( .A(G1986), .B(G24), .Z(n1002) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(KEYINPUT58), .B(n1004), .ZN(n1005) );
  NOR2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1017) );
  XNOR2_X1 U1095 ( .A(KEYINPUT59), .B(G1348), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(n1007), .B(G4), .ZN(n1014) );
  XNOR2_X1 U1097 ( .A(G1956), .B(G20), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(G1341), .B(G19), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(G1981), .B(G6), .ZN(n1008) );
  NOR2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1101 ( .A(KEYINPUT127), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1104 ( .A(KEYINPUT60), .B(n1015), .Z(n1016) );
  NAND2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(G21), .B(G1966), .ZN(n1018) );
  NOR2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1108 ( .A(KEYINPUT61), .B(n1020), .Z(n1021) );
  NOR2_X1 U1109 ( .A1(G16), .A2(n1021), .ZN(n1026) );
  NOR2_X1 U1110 ( .A1(G29), .A2(KEYINPUT55), .ZN(n1022) );
  NAND2_X1 U1111 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1112 ( .A1(G11), .A2(n1024), .ZN(n1025) );
  NOR2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1116 ( .A(n1031), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

