//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 0 0 1 1 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 1 0 0 0 0 1 0 1 1 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0 0 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n859, new_n860, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982;
  XNOR2_X1  g000(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n202));
  XNOR2_X1  g001(.A(G1gat), .B(G29gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G57gat), .B(G85gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT73), .ZN(new_n208));
  AND2_X1   g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G155gat), .ZN(new_n212));
  INV_X1    g011(.A(G162gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n214), .A2(KEYINPUT73), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G148gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G141gat), .ZN(new_n219));
  INV_X1    g018(.A(G141gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G148gat), .ZN(new_n221));
  AOI22_X1  g020(.A1(new_n219), .A2(new_n221), .B1(KEYINPUT2), .B2(new_n215), .ZN(new_n222));
  OR2_X1    g021(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT75), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n215), .B1(new_n214), .B2(KEYINPUT2), .ZN(new_n225));
  OR2_X1    g024(.A1(KEYINPUT74), .A2(G141gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(KEYINPUT74), .A2(G141gat), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n218), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n219), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n224), .B(new_n225), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  AND2_X1   g030(.A1(KEYINPUT74), .A2(G141gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(KEYINPUT74), .A2(G141gat), .ZN(new_n233));
  OAI21_X1  g032(.A(G148gat), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(new_n219), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n224), .B1(new_n235), .B2(new_n225), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n223), .B1(new_n231), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G120gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G113gat), .ZN(new_n239));
  INV_X1    g038(.A(G113gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G120gat), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT1), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G127gat), .B(G134gat), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT67), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G134gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(G127gat), .ZN(new_n246));
  INV_X1    g045(.A(G127gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(G134gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n250));
  XNOR2_X1  g049(.A(G113gat), .B(G120gat), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n249), .B(new_n250), .C1(new_n251), .C2(KEYINPUT1), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n244), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT68), .B(G113gat), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n239), .B1(new_n254), .B2(new_n238), .ZN(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT70), .B(KEYINPUT1), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n249), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n243), .A2(KEYINPUT69), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n255), .A2(new_n257), .A3(new_n259), .A4(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n253), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(KEYINPUT4), .B1(new_n237), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n217), .A2(new_n222), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT74), .B(G141gat), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n229), .B1(new_n265), .B2(G148gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT2), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n209), .B1(new_n267), .B2(new_n210), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT75), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n264), .B1(new_n269), .B2(new_n230), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n240), .A2(KEYINPUT68), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n240), .A2(KEYINPUT68), .ZN(new_n273));
  OAI21_X1  g072(.A(G120gat), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n256), .B1(new_n274), .B2(new_n239), .ZN(new_n275));
  AND3_X1   g074(.A1(new_n246), .A2(new_n248), .A3(KEYINPUT69), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT69), .B1(new_n246), .B2(new_n248), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n275), .A2(new_n278), .B1(new_n244), .B2(new_n252), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n270), .A2(new_n271), .A3(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n279), .B1(new_n270), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n237), .A2(KEYINPUT3), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n263), .A2(new_n280), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G225gat), .A2(G233gat), .ZN(new_n286));
  XOR2_X1   g085(.A(new_n286), .B(KEYINPUT77), .Z(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n237), .A2(new_n262), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n269), .A2(new_n230), .ZN(new_n290));
  AOI22_X1  g089(.A1(new_n290), .A2(new_n223), .B1(new_n253), .B2(new_n261), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n287), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  AOI22_X1  g091(.A1(new_n285), .A2(new_n288), .B1(KEYINPUT5), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n263), .A2(new_n280), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n223), .B(new_n282), .C1(new_n231), .C2(new_n236), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT3), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n295), .B(new_n262), .C1(new_n296), .C2(new_n270), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n294), .A2(KEYINPUT5), .A3(new_n288), .A4(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n207), .B1(new_n293), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT79), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT6), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n292), .A2(KEYINPUT5), .ZN(new_n304));
  NOR3_X1   g103(.A1(new_n237), .A2(new_n262), .A3(KEYINPUT4), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n271), .B1(new_n270), .B2(new_n279), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n297), .B(new_n288), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n206), .B1(new_n308), .B2(new_n298), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT79), .B1(new_n309), .B2(KEYINPUT6), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(new_n206), .A3(new_n298), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n303), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n302), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT65), .ZN(new_n317));
  OR2_X1    g116(.A1(new_n317), .A2(KEYINPUT25), .ZN(new_n318));
  OAI21_X1  g117(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NOR3_X1   g119(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n316), .B(new_n318), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(G183gat), .A2(G190gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT24), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT64), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT64), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n328), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n325), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT23), .ZN(new_n331));
  INV_X1    g130(.A(G169gat), .ZN(new_n332));
  INV_X1    g131(.A(G176gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n334), .A2(new_n319), .B1(G169gat), .B2(G176gat), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n322), .B(new_n330), .C1(new_n317), .C2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n316), .B1(new_n320), .B2(new_n321), .ZN(new_n337));
  AND3_X1   g136(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n338), .B1(new_n324), .B2(new_n323), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT25), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(G190gat), .ZN(new_n341));
  AND2_X1   g140(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  OR3_X1    g146(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(new_n316), .A3(new_n349), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n341), .B(new_n345), .C1(new_n342), .C2(new_n343), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n347), .A2(new_n350), .A3(new_n324), .A4(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n340), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(G226gat), .ZN(new_n354));
  INV_X1    g153(.A(G233gat), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G197gat), .B(G204gat), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT22), .ZN(new_n359));
  INV_X1    g158(.A(G211gat), .ZN(new_n360));
  INV_X1    g159(.A(G218gat), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AND2_X1   g161(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  XOR2_X1   g162(.A(G211gat), .B(G218gat), .Z(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT71), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n363), .B(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n356), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT72), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT72), .ZN(new_n372));
  AOI211_X1 g171(.A(new_n372), .B(new_n356), .C1(new_n353), .C2(new_n368), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n357), .B(new_n367), .C1(new_n371), .C2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n369), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n357), .B1(new_n375), .B2(new_n356), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n366), .ZN(new_n377));
  XOR2_X1   g176(.A(G8gat), .B(G36gat), .Z(new_n378));
  XNOR2_X1  g177(.A(new_n378), .B(G64gat), .ZN(new_n379));
  INV_X1    g178(.A(G92gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n379), .B(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n374), .A2(new_n377), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT30), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n381), .B1(new_n374), .B2(new_n377), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n374), .A2(new_n377), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT30), .ZN(new_n387));
  INV_X1    g186(.A(new_n381), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n385), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(G227gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n393), .A2(new_n355), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n262), .A2(new_n340), .A3(new_n352), .A4(new_n336), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n353), .A2(new_n279), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n395), .A2(new_n394), .A3(new_n396), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT34), .ZN(new_n399));
  AND3_X1   g198(.A1(new_n398), .A2(KEYINPUT32), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n399), .B1(new_n398), .B2(KEYINPUT32), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n397), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n398), .A2(KEYINPUT32), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT34), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n398), .A2(KEYINPUT32), .A3(new_n399), .ZN(new_n405));
  INV_X1    g204(.A(new_n397), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(G15gat), .B(G43gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n408), .B(G71gat), .ZN(new_n409));
  INV_X1    g208(.A(G99gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n398), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n411), .B1(new_n412), .B2(KEYINPUT33), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n402), .A2(new_n407), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n402), .A2(new_n407), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n413), .ZN(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(KEYINPUT81), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(G50gat), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n366), .B1(new_n295), .B2(new_n368), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(G228gat), .A2(G233gat), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n358), .A2(KEYINPUT82), .A3(new_n362), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n364), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT82), .B1(new_n358), .B2(new_n362), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n368), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NOR3_X1   g227(.A1(new_n363), .A2(KEYINPUT82), .A3(new_n364), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n282), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n430), .A2(KEYINPUT83), .A3(new_n237), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT83), .B1(new_n430), .B2(new_n237), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n423), .B(new_n424), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n366), .A2(new_n368), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n270), .B1(new_n434), .B2(new_n296), .ZN(new_n435));
  OAI211_X1 g234(.A(G228gat), .B(G233gat), .C1(new_n435), .C2(new_n422), .ZN(new_n436));
  XNOR2_X1  g235(.A(G78gat), .B(G106gat), .ZN(new_n437));
  INV_X1    g236(.A(G22gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n433), .A2(new_n436), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n440), .B1(new_n433), .B2(new_n436), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n421), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n433), .A2(new_n436), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n439), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n433), .A2(new_n436), .A3(new_n440), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n445), .A2(new_n420), .A3(new_n446), .ZN(new_n447));
  AND4_X1   g246(.A1(new_n415), .A2(new_n417), .A3(new_n443), .A4(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n315), .A2(new_n392), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT35), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n443), .A2(new_n447), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n206), .B(KEYINPUT85), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n308), .A2(new_n298), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n300), .A2(new_n302), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n314), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n415), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n414), .B1(new_n402), .B2(new_n407), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT35), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n451), .A2(new_n455), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n386), .A2(new_n388), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n461), .A2(KEYINPUT30), .A3(new_n382), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n462), .A2(KEYINPUT84), .A3(new_n389), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT84), .B1(new_n462), .B2(new_n389), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT88), .B1(new_n460), .B2(new_n465), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n417), .A2(new_n443), .A3(new_n447), .A4(new_n415), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n467), .A2(KEYINPUT35), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT88), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT84), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n470), .B1(new_n385), .B2(new_n390), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n462), .A2(KEYINPUT84), .A3(new_n389), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n468), .A2(new_n469), .A3(new_n473), .A4(new_n455), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n450), .A2(new_n466), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n453), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n288), .B1(new_n294), .B2(new_n297), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  OR2_X1    g277(.A1(new_n289), .A2(new_n291), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n478), .B(KEYINPUT39), .C1(new_n287), .C2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT86), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT39), .ZN(new_n482));
  AOI211_X1 g281(.A(new_n481), .B(new_n452), .C1(new_n477), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n294), .A2(new_n297), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n484), .A2(new_n482), .A3(new_n287), .ZN(new_n485));
  INV_X1    g284(.A(new_n452), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT86), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n480), .B1(new_n483), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT40), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n476), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI211_X1 g289(.A(KEYINPUT40), .B(new_n480), .C1(new_n483), .C2(new_n487), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n490), .A2(new_n472), .A3(new_n471), .A4(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n309), .A2(KEYINPUT6), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n313), .B1(new_n493), .B2(new_n453), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n356), .B1(new_n353), .B2(new_n368), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(KEYINPUT72), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n496), .A2(KEYINPUT87), .A3(new_n357), .A4(new_n366), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n357), .B(new_n366), .C1(new_n371), .C2(new_n373), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT87), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n376), .A2(new_n367), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n497), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT37), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT37), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n388), .B1(new_n386), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT38), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n374), .A2(KEYINPUT37), .A3(new_n377), .ZN(new_n507));
  AND3_X1   g306(.A1(new_n505), .A2(KEYINPUT38), .A3(new_n507), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n461), .B(new_n494), .C1(new_n506), .C2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n492), .A2(new_n509), .A3(new_n451), .ZN(new_n510));
  INV_X1    g309(.A(new_n451), .ZN(new_n511));
  INV_X1    g310(.A(new_n311), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n300), .A2(new_n302), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n512), .B1(new_n513), .B2(KEYINPUT79), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n313), .B1(new_n514), .B2(new_n303), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n511), .B1(new_n515), .B2(new_n391), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n458), .B(KEYINPUT36), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n510), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n475), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT15), .ZN(new_n520));
  XOR2_X1   g319(.A(KEYINPUT92), .B(G50gat), .Z(new_n521));
  NOR2_X1   g320(.A1(new_n521), .A2(G43gat), .ZN(new_n522));
  INV_X1    g321(.A(G50gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(G43gat), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT91), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n520), .B1(new_n522), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(G43gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(G50gat), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n529), .A2(new_n524), .A3(KEYINPUT15), .ZN(new_n530));
  NAND2_X1  g329(.A1(G29gat), .A2(G36gat), .ZN(new_n531));
  NOR2_X1   g330(.A1(G29gat), .A2(G36gat), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT14), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n527), .A2(new_n530), .A3(new_n531), .A4(new_n534), .ZN(new_n535));
  OAI211_X1 g334(.A(KEYINPUT89), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n531), .B(new_n536), .C1(new_n534), .C2(KEYINPUT89), .ZN(new_n537));
  INV_X1    g336(.A(new_n530), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n537), .A2(KEYINPUT90), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT90), .B1(new_n537), .B2(new_n538), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n535), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT17), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G15gat), .B(G22gat), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT16), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n544), .B1(new_n545), .B2(G1gat), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n546), .B1(G1gat), .B2(new_n544), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(G8gat), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  OAI211_X1 g348(.A(KEYINPUT17), .B(new_n535), .C1(new_n539), .C2(new_n540), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n543), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n541), .A2(new_n548), .ZN(new_n552));
  NAND2_X1  g351(.A1(G229gat), .A2(G233gat), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(KEYINPUT93), .A2(KEYINPUT18), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n541), .B(new_n548), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n553), .B(KEYINPUT13), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n555), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n551), .A2(new_n552), .A3(new_n553), .A4(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n556), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G113gat), .B(G141gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(G197gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT11), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(new_n332), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT12), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n563), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n556), .A2(new_n568), .A3(new_n560), .A4(new_n562), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G57gat), .B(G64gat), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  OR2_X1    g373(.A1(G71gat), .A2(G78gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(G71gat), .A2(G78gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT9), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n574), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n576), .B(new_n575), .C1(new_n573), .C2(new_n578), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT95), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(G106gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n410), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G99gat), .A2(G106gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G85gat), .A2(G92gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT7), .ZN(new_n590));
  INV_X1    g389(.A(G85gat), .ZN(new_n591));
  AOI22_X1  g390(.A1(KEYINPUT8), .A2(new_n587), .B1(new_n591), .B2(new_n380), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n588), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n590), .A2(new_n588), .A3(new_n592), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n594), .A2(KEYINPUT98), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT98), .ZN(new_n597));
  AND3_X1   g396(.A1(new_n590), .A2(new_n588), .A3(new_n592), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n597), .B1(new_n598), .B2(new_n593), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n584), .A2(KEYINPUT10), .A3(new_n596), .A4(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT100), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n581), .B(new_n580), .C1(new_n598), .C2(new_n593), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n594), .A2(new_n582), .A3(new_n595), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT10), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n601), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI211_X1 g405(.A(KEYINPUT100), .B(KEYINPUT10), .C1(new_n602), .C2(new_n603), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n600), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G230gat), .A2(G233gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n609), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n602), .A2(new_n603), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G120gat), .B(G148gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT101), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(new_n333), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(G204gat), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n613), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n572), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n548), .B1(new_n584), .B2(KEYINPUT21), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT96), .B(KEYINPUT20), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n625), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n623), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n628), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n630), .A2(new_n626), .A3(new_n622), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(KEYINPUT21), .B1(new_n580), .B2(new_n581), .ZN(new_n633));
  XOR2_X1   g432(.A(G127gat), .B(G155gat), .Z(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G183gat), .B(G211gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(G231gat), .A2(G233gat), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n637), .B(new_n638), .Z(new_n639));
  OR2_X1    g438(.A1(new_n632), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n632), .A2(new_n639), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G134gat), .B(G162gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT99), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(G218gat), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n596), .A2(new_n599), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n543), .A2(new_n646), .A3(new_n550), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n541), .A2(new_n596), .A3(new_n599), .ZN(new_n648));
  NAND3_X1  g447(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT97), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(G190gat), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n653), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n647), .A2(new_n648), .A3(new_n649), .A4(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n645), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n654), .A2(new_n645), .A3(new_n656), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n642), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n519), .A2(new_n621), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(new_n515), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g464(.A1(new_n662), .A2(new_n473), .ZN(new_n666));
  INV_X1    g465(.A(G8gat), .ZN(new_n667));
  OAI21_X1  g466(.A(KEYINPUT42), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n545), .A2(new_n667), .ZN(new_n669));
  NAND2_X1  g468(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n666), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT102), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT42), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  MUX2_X1   g474(.A(new_n673), .B(KEYINPUT102), .S(new_n675), .Z(G1325gat));
  INV_X1    g475(.A(new_n517), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n663), .A2(G15gat), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(G15gat), .B1(new_n663), .B2(new_n458), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(G1326gat));
  INV_X1    g479(.A(KEYINPUT43), .ZN(new_n681));
  OR3_X1    g480(.A1(new_n662), .A2(KEYINPUT103), .A3(new_n451), .ZN(new_n682));
  OAI21_X1  g481(.A(KEYINPUT103), .B1(new_n662), .B2(new_n451), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n682), .A2(new_n681), .A3(new_n683), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n685), .A2(G22gat), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(G22gat), .B1(new_n685), .B2(new_n686), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(G1327gat));
  NAND2_X1  g488(.A1(new_n519), .A2(new_n660), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n621), .A2(new_n642), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(G29gat), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n692), .A2(new_n693), .A3(new_n515), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n694), .A2(KEYINPUT104), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(KEYINPUT104), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT45), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT105), .ZN(new_n701));
  INV_X1    g500(.A(new_n659), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n701), .B1(new_n702), .B2(new_n657), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n658), .A2(KEYINPUT105), .A3(new_n659), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n519), .A2(new_n700), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n700), .B1(new_n519), .B2(new_n660), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n706), .B1(new_n707), .B2(KEYINPUT106), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n703), .A2(new_n704), .ZN(new_n709));
  AOI211_X1 g508(.A(KEYINPUT44), .B(new_n709), .C1(new_n475), .C2(new_n518), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n691), .B1(new_n708), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(G29gat), .B1(new_n714), .B2(new_n315), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n695), .A2(KEYINPUT45), .A3(new_n696), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n699), .A2(new_n715), .A3(new_n716), .ZN(G1328gat));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n718), .B1(new_n714), .B2(new_n473), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n713), .A2(KEYINPUT107), .A3(new_n465), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n719), .A2(G36gat), .A3(new_n720), .ZN(new_n721));
  NOR4_X1   g520(.A1(new_n690), .A2(G36gat), .A3(new_n473), .A4(new_n691), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT46), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(G1329gat));
  AOI21_X1  g523(.A(new_n528), .B1(new_n713), .B2(new_n677), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n456), .A2(new_n457), .A3(G43gat), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n692), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n726), .A2(KEYINPUT47), .A3(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT47), .ZN(new_n730));
  INV_X1    g529(.A(new_n728), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n730), .B1(new_n725), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n729), .A2(new_n732), .ZN(G1330gat));
  INV_X1    g532(.A(KEYINPUT48), .ZN(new_n734));
  INV_X1    g533(.A(new_n691), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n690), .A2(KEYINPUT44), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n710), .B1(new_n736), .B2(new_n711), .ZN(new_n737));
  INV_X1    g536(.A(new_n712), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n511), .B(new_n735), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n521), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n692), .A2(new_n521), .A3(new_n511), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n734), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n742), .ZN(new_n744));
  AOI211_X1 g543(.A(KEYINPUT48), .B(new_n744), .C1(new_n739), .C2(new_n740), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n743), .A2(new_n745), .ZN(G1331gat));
  NAND3_X1  g545(.A1(new_n661), .A2(new_n620), .A3(new_n572), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT108), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n748), .A2(new_n519), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n515), .B(KEYINPUT109), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g551(.A1(new_n749), .A2(new_n465), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n754));
  XOR2_X1   g553(.A(KEYINPUT49), .B(G64gat), .Z(new_n755));
  OAI21_X1  g554(.A(new_n754), .B1(new_n753), .B2(new_n755), .ZN(G1333gat));
  XOR2_X1   g555(.A(new_n458), .B(KEYINPUT110), .Z(new_n757));
  AOI21_X1  g556(.A(G71gat), .B1(new_n749), .B2(new_n757), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n677), .A2(G71gat), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n758), .B1(new_n749), .B2(new_n759), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n760), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g560(.A1(new_n749), .A2(new_n511), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g562(.A1(new_n642), .A2(new_n572), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n764), .B(KEYINPUT111), .Z(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n620), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(new_n737), .B2(new_n738), .ZN(new_n768));
  OAI21_X1  g567(.A(G85gat), .B1(new_n768), .B2(new_n315), .ZN(new_n769));
  INV_X1    g568(.A(new_n660), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n475), .B2(new_n518), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n765), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT112), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n771), .A2(KEYINPUT51), .A3(new_n765), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n776), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(KEYINPUT112), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n515), .A2(new_n591), .A3(new_n620), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n769), .B1(new_n780), .B2(new_n781), .ZN(G1336gat));
  OAI21_X1  g581(.A(G92gat), .B1(new_n768), .B2(new_n473), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784));
  INV_X1    g583(.A(new_n620), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n473), .A2(G92gat), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n777), .A2(new_n779), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT114), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n777), .A2(new_n779), .A3(new_n789), .A4(new_n786), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n783), .A2(new_n784), .A3(new_n788), .A4(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT51), .B1(new_n771), .B2(new_n765), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n786), .B1(new_n778), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT113), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI211_X1 g594(.A(KEYINPUT113), .B(new_n786), .C1(new_n778), .C2(new_n792), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n766), .B1(new_n708), .B2(new_n712), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n380), .B1(new_n798), .B2(new_n465), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT52), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n791), .A2(new_n800), .ZN(G1337gat));
  OAI21_X1  g600(.A(G99gat), .B1(new_n768), .B2(new_n517), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n458), .A2(new_n620), .A3(new_n410), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n802), .B1(new_n780), .B2(new_n803), .ZN(G1338gat));
  OAI21_X1  g603(.A(G106gat), .B1(new_n768), .B2(new_n451), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n785), .A2(G106gat), .A3(new_n451), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n777), .A2(new_n779), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(KEYINPUT116), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n777), .A2(new_n779), .A3(new_n810), .A4(new_n807), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n805), .A2(new_n806), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n807), .B1(new_n778), .B2(new_n792), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT115), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n815), .B(new_n807), .C1(new_n778), .C2(new_n792), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n585), .B1(new_n798), .B2(new_n511), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT53), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n812), .A2(new_n819), .ZN(G1339gat));
  NAND2_X1  g619(.A1(new_n570), .A2(new_n571), .ZN(new_n821));
  NOR4_X1   g620(.A1(new_n642), .A2(new_n821), .A3(new_n660), .A4(new_n620), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT10), .B1(new_n602), .B2(new_n603), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(new_n601), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n611), .B1(new_n825), .B2(new_n600), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n611), .B(new_n600), .C1(new_n606), .C2(new_n607), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT54), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n608), .A2(new_n830), .A3(new_n609), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n617), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n823), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n610), .A2(KEYINPUT54), .A3(new_n827), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n834), .A2(KEYINPUT55), .A3(new_n617), .A4(new_n831), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n833), .A2(new_n618), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n557), .A2(new_n559), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n553), .B1(new_n551), .B2(new_n552), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n567), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n571), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n836), .A2(new_n703), .A3(new_n704), .A4(new_n840), .ZN(new_n841));
  AOI22_X1  g640(.A1(new_n836), .A2(new_n821), .B1(new_n620), .B2(new_n840), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n841), .B1(new_n842), .B2(new_n705), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n822), .B1(new_n843), .B2(new_n642), .ZN(new_n844));
  INV_X1    g643(.A(new_n750), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n844), .A2(new_n465), .A3(new_n845), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n846), .A2(new_n448), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n847), .B(new_n821), .C1(new_n272), .C2(new_n273), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n843), .A2(new_n642), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n661), .A2(new_n785), .A3(new_n572), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n465), .A2(new_n315), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n851), .A2(new_n448), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(G113gat), .B1(new_n853), .B2(new_n572), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n848), .A2(new_n854), .ZN(G1340gat));
  NAND3_X1  g654(.A1(new_n847), .A2(new_n238), .A3(new_n620), .ZN(new_n856));
  OAI21_X1  g655(.A(G120gat), .B1(new_n853), .B2(new_n785), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(G1341gat));
  INV_X1    g657(.A(new_n642), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n847), .A2(new_n247), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(G127gat), .B1(new_n853), .B2(new_n642), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XOR2_X1   g661(.A(new_n862), .B(KEYINPUT117), .Z(G1342gat));
  NAND4_X1  g662(.A1(new_n846), .A2(new_n245), .A3(new_n660), .A4(new_n448), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(KEYINPUT56), .ZN(new_n865));
  XOR2_X1   g664(.A(new_n865), .B(KEYINPUT119), .Z(new_n866));
  NOR2_X1   g665(.A1(new_n864), .A2(KEYINPUT56), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(KEYINPUT118), .ZN(new_n868));
  OAI21_X1  g667(.A(G134gat), .B1(new_n853), .B2(new_n770), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n866), .A2(new_n868), .A3(new_n869), .ZN(G1343gat));
  OAI21_X1  g669(.A(new_n841), .B1(new_n842), .B2(new_n660), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n822), .B1(new_n871), .B2(new_n642), .ZN(new_n872));
  OAI21_X1  g671(.A(KEYINPUT57), .B1(new_n872), .B2(new_n451), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n852), .A2(new_n517), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n840), .A2(new_n620), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n833), .A2(new_n618), .A3(new_n835), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(new_n572), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n709), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n859), .B1(new_n879), .B2(new_n841), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n875), .B(new_n511), .C1(new_n880), .C2(new_n822), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n873), .A2(new_n821), .A3(new_n874), .A4(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(new_n265), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT120), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n517), .A2(new_n511), .ZN(new_n886));
  NOR4_X1   g685(.A1(new_n844), .A2(new_n465), .A3(new_n845), .A4(new_n886), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n572), .A2(G141gat), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n884), .A2(new_n885), .A3(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n885), .B1(new_n884), .B2(new_n889), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT58), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n884), .A2(new_n889), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(KEYINPUT120), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT58), .B1(new_n896), .B2(new_n890), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n894), .A2(new_n897), .ZN(G1344gat));
  NAND3_X1  g697(.A1(new_n887), .A2(new_n218), .A3(new_n620), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n822), .B(KEYINPUT121), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n836), .A2(new_n660), .A3(new_n840), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n902), .B1(new_n842), .B2(new_n660), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n642), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT57), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n511), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n851), .A2(new_n511), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT57), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n906), .A2(new_n908), .A3(new_n620), .A4(new_n874), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n218), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI22_X1  g710(.A1(new_n511), .A2(new_n905), .B1(new_n907), .B2(KEYINPUT57), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n912), .A2(KEYINPUT122), .A3(new_n620), .A4(new_n874), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n900), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n873), .A2(new_n874), .A3(new_n881), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n900), .B1(new_n915), .B2(new_n785), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n916), .A2(new_n218), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n899), .B1(new_n914), .B2(new_n917), .ZN(G1345gat));
  NOR3_X1   g717(.A1(new_n915), .A2(new_n212), .A3(new_n642), .ZN(new_n919));
  AOI21_X1  g718(.A(G155gat), .B1(new_n887), .B2(new_n859), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n919), .A2(new_n920), .ZN(G1346gat));
  NOR3_X1   g720(.A1(new_n915), .A2(new_n213), .A3(new_n709), .ZN(new_n922));
  AOI21_X1  g721(.A(G162gat), .B1(new_n887), .B2(new_n660), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n922), .A2(new_n923), .ZN(G1347gat));
  NOR2_X1   g723(.A1(new_n750), .A2(new_n473), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n451), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(new_n757), .A3(new_n851), .ZN(new_n928));
  OAI21_X1  g727(.A(G169gat), .B1(new_n928), .B2(new_n572), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT123), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n844), .A2(new_n515), .A3(new_n473), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(new_n448), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(new_n332), .A3(new_n821), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n930), .A2(new_n934), .ZN(G1348gat));
  NOR3_X1   g734(.A1(new_n928), .A2(new_n333), .A3(new_n785), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n933), .A2(new_n620), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n936), .B1(new_n937), .B2(new_n333), .ZN(G1349gat));
  OAI21_X1  g737(.A(KEYINPUT124), .B1(new_n928), .B2(new_n642), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n851), .A2(new_n757), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n940), .A2(new_n941), .A3(new_n859), .A4(new_n927), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n939), .A2(new_n942), .A3(G183gat), .ZN(new_n943));
  OAI211_X1 g742(.A(new_n933), .B(new_n859), .C1(new_n343), .C2(new_n342), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g745(.A(G190gat), .B1(new_n928), .B2(new_n770), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT61), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n933), .A2(new_n341), .A3(new_n705), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(G1351gat));
  INV_X1    g749(.A(new_n886), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n931), .A2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(G197gat), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n953), .A2(new_n954), .A3(new_n821), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n906), .A2(new_n908), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n925), .A2(new_n517), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT125), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n956), .A2(new_n958), .A3(new_n572), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n955), .B1(new_n959), .B2(new_n954), .ZN(G1352gat));
  NOR2_X1   g759(.A1(new_n956), .A2(new_n958), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n961), .A2(new_n962), .A3(new_n620), .ZN(new_n963));
  INV_X1    g762(.A(new_n958), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n964), .A2(new_n912), .A3(new_n620), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(KEYINPUT126), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n963), .A2(new_n966), .A3(G204gat), .ZN(new_n967));
  OR3_X1    g766(.A1(new_n952), .A2(G204gat), .A3(new_n785), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(KEYINPUT62), .ZN(new_n969));
  OR2_X1    g768(.A1(new_n968), .A2(KEYINPUT62), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n967), .A2(new_n969), .A3(new_n970), .ZN(G1353gat));
  NAND3_X1  g770(.A1(new_n953), .A2(new_n360), .A3(new_n859), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n912), .A2(new_n859), .A3(new_n517), .A4(new_n925), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n973), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT63), .B1(new_n973), .B2(G211gat), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(G1354gat));
  INV_X1    g775(.A(KEYINPUT127), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n961), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n964), .A2(new_n912), .A3(new_n977), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(new_n660), .ZN(new_n980));
  OAI21_X1  g779(.A(G218gat), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n953), .A2(new_n361), .A3(new_n705), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(G1355gat));
endmodule


