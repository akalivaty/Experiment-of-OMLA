

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753;

  NAND2_X1 U368 ( .A1(n546), .A2(n625), .ZN(n548) );
  XNOR2_X1 U369 ( .A(KEYINPUT69), .B(KEYINPUT34), .ZN(n523) );
  BUF_X1 U370 ( .A(G107), .Z(n383) );
  NOR2_X2 U371 ( .A1(n442), .A2(n556), .ZN(n443) );
  INV_X1 U372 ( .A(n611), .ZN(n345) );
  NOR2_X1 U373 ( .A1(n662), .A2(n520), .ZN(n424) );
  NAND2_X1 U374 ( .A1(n424), .A2(n558), .ZN(n566) );
  XNOR2_X1 U375 ( .A(n512), .B(n511), .ZN(n653) );
  INV_X1 U376 ( .A(G953), .ZN(n742) );
  NOR2_X1 U377 ( .A1(n576), .A2(n575), .ZN(n717) );
  BUF_X1 U378 ( .A(G143), .Z(n379) );
  NOR2_X1 U379 ( .A1(n653), .A2(G902), .ZN(n513) );
  XNOR2_X2 U380 ( .A(n586), .B(KEYINPUT19), .ZN(n574) );
  NAND2_X2 U381 ( .A1(n421), .A2(n420), .ZN(n586) );
  AND2_X2 U382 ( .A1(n423), .A2(n422), .ZN(n421) );
  OR2_X1 U383 ( .A1(n627), .A2(n626), .ZN(n549) );
  NAND2_X1 U384 ( .A1(n549), .A2(KEYINPUT44), .ZN(n357) );
  NOR2_X1 U385 ( .A1(n532), .A2(n583), .ZN(n376) );
  AND2_X1 U386 ( .A1(n356), .A2(n355), .ZN(n354) );
  XNOR2_X1 U387 ( .A(n357), .B(n550), .ZN(n353) );
  INV_X1 U388 ( .A(n621), .ZN(n364) );
  NOR2_X1 U389 ( .A1(n702), .A2(n539), .ZN(n363) );
  AND2_X1 U390 ( .A1(n515), .A2(n514), .ZN(n366) );
  XNOR2_X1 U391 ( .A(n661), .B(n489), .ZN(n583) );
  INV_X1 U392 ( .A(KEYINPUT96), .ZN(n539) );
  BUF_X1 U393 ( .A(KEYINPUT45), .Z(n551) );
  INV_X1 U394 ( .A(KEYINPUT48), .ZN(n350) );
  INV_X1 U395 ( .A(KEYINPUT41), .ZN(n561) );
  XNOR2_X1 U396 ( .A(n351), .B(n350), .ZN(n609) );
  NAND2_X1 U397 ( .A1(n354), .A2(n353), .ZN(n352) );
  NAND2_X1 U398 ( .A1(n364), .A2(n363), .ZN(n361) );
  NAND2_X1 U399 ( .A1(n360), .A2(n678), .ZN(n358) );
  AND2_X1 U400 ( .A1(n621), .A2(n539), .ZN(n359) );
  XNOR2_X1 U401 ( .A(n565), .B(n349), .ZN(n751) );
  AND2_X1 U402 ( .A1(n583), .A2(n544), .ZN(n545) );
  XNOR2_X1 U403 ( .A(n562), .B(n561), .ZN(n694) );
  NOR2_X1 U404 ( .A1(n679), .A2(n677), .ZN(n562) );
  INV_X1 U405 ( .A(n678), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n604), .B(KEYINPUT38), .ZN(n675) );
  XNOR2_X1 U407 ( .A(n630), .B(n632), .ZN(n633) );
  XNOR2_X1 U408 ( .A(n644), .B(KEYINPUT62), .ZN(n645) );
  XNOR2_X1 U409 ( .A(n638), .B(n637), .ZN(n639) );
  INV_X1 U410 ( .A(n476), .ZN(n348) );
  XNOR2_X1 U411 ( .A(n564), .B(KEYINPUT109), .ZN(n349) );
  XNOR2_X1 U412 ( .A(n475), .B(n474), .ZN(n476) );
  BUF_X1 U413 ( .A(KEYINPUT64), .Z(n550) );
  XNOR2_X2 U414 ( .A(n347), .B(n516), .ZN(n627) );
  NAND2_X1 U415 ( .A1(n519), .A2(n366), .ZN(n347) );
  NAND2_X1 U416 ( .A1(n519), .A2(n545), .ZN(n625) );
  XNOR2_X2 U417 ( .A(n477), .B(n348), .ZN(n519) );
  NAND2_X1 U418 ( .A1(n599), .A2(n598), .ZN(n351) );
  NOR2_X2 U419 ( .A1(n627), .A2(n626), .ZN(n398) );
  XNOR2_X2 U420 ( .A(n352), .B(n551), .ZN(n612) );
  XNOR2_X1 U421 ( .A(n375), .B(n374), .ZN(n355) );
  NAND2_X1 U422 ( .A1(n531), .A2(n530), .ZN(n356) );
  NOR2_X1 U423 ( .A1(n359), .A2(n358), .ZN(n362) );
  NAND2_X1 U424 ( .A1(n702), .A2(n539), .ZN(n360) );
  XNOR2_X2 U425 ( .A(n535), .B(KEYINPUT31), .ZN(n621) );
  NAND2_X1 U426 ( .A1(n362), .A2(n361), .ZN(n546) );
  OR2_X2 U427 ( .A1(n560), .A2(n367), .ZN(n420) );
  XNOR2_X2 U428 ( .A(n378), .B(KEYINPUT0), .ZN(n538) );
  NOR2_X2 U429 ( .A1(n574), .A2(n443), .ZN(n378) );
  INV_X1 U430 ( .A(KEYINPUT83), .ZN(n374) );
  XNOR2_X1 U431 ( .A(G119), .B(G116), .ZN(n419) );
  OR2_X1 U432 ( .A1(n674), .A2(KEYINPUT86), .ZN(n422) );
  INV_X1 U433 ( .A(n570), .ZN(n381) );
  OR2_X1 U434 ( .A1(n644), .A2(G902), .ZN(n488) );
  NAND2_X1 U435 ( .A1(n393), .A2(n345), .ZN(n392) );
  BUF_X1 U436 ( .A(n661), .Z(n382) );
  XNOR2_X1 U437 ( .A(n410), .B(n505), .ZN(n662) );
  NAND2_X1 U438 ( .A1(n606), .A2(n703), .ZN(n678) );
  NAND2_X1 U439 ( .A1(n552), .A2(n400), .ZN(n399) );
  INV_X1 U440 ( .A(KEYINPUT79), .ZN(n400) );
  AND2_X1 U441 ( .A1(n365), .A2(n408), .ZN(n401) );
  XNOR2_X1 U442 ( .A(G131), .B(G134), .ZN(n478) );
  XNOR2_X1 U443 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n426) );
  XNOR2_X1 U444 ( .A(G125), .B(G146), .ZN(n458) );
  NOR2_X1 U445 ( .A1(n520), .A2(n570), .ZN(n409) );
  XNOR2_X1 U446 ( .A(n434), .B(KEYINPUT90), .ZN(n435) );
  XNOR2_X1 U447 ( .A(n416), .B(G122), .ZN(n415) );
  XNOR2_X1 U448 ( .A(G119), .B(G128), .ZN(n490) );
  XNOR2_X1 U449 ( .A(KEYINPUT24), .B(KEYINPUT78), .ZN(n492) );
  XNOR2_X1 U450 ( .A(G134), .B(G122), .ZN(n445) );
  INV_X1 U451 ( .A(G128), .ZN(n429) );
  XNOR2_X1 U452 ( .A(n412), .B(n411), .ZN(n496) );
  INV_X1 U453 ( .A(KEYINPUT8), .ZN(n411) );
  NAND2_X1 U454 ( .A1(n742), .A2(G234), .ZN(n412) );
  XNOR2_X1 U455 ( .A(G113), .B(G131), .ZN(n460) );
  XOR2_X1 U456 ( .A(G122), .B(G104), .Z(n461) );
  BUF_X1 U457 ( .A(n673), .Z(n693) );
  AND2_X1 U458 ( .A1(n568), .A2(n380), .ZN(n580) );
  AND2_X1 U459 ( .A1(n569), .A2(n381), .ZN(n380) );
  BUF_X1 U460 ( .A(n521), .Z(n658) );
  XNOR2_X1 U461 ( .A(n389), .B(KEYINPUT80), .ZN(n699) );
  NAND2_X1 U462 ( .A1(n392), .A2(n391), .ZN(n390) );
  INV_X1 U463 ( .A(KEYINPUT2), .ZN(n391) );
  AND2_X1 U464 ( .A1(n519), .A2(n518), .ZN(n626) );
  AND2_X1 U465 ( .A1(n581), .A2(n715), .ZN(n365) );
  NAND2_X1 U466 ( .A1(n674), .A2(KEYINPUT86), .ZN(n367) );
  AND2_X1 U467 ( .A1(n399), .A2(KEYINPUT79), .ZN(n368) );
  XNOR2_X1 U468 ( .A(KEYINPUT15), .B(G902), .ZN(n552) );
  NAND2_X1 U469 ( .A1(n610), .A2(KEYINPUT2), .ZN(n369) );
  NAND2_X1 U470 ( .A1(n610), .A2(KEYINPUT79), .ZN(n370) );
  AND2_X1 U471 ( .A1(n370), .A2(n399), .ZN(n371) );
  NOR2_X1 U472 ( .A1(n742), .A2(G952), .ZN(n656) );
  INV_X1 U473 ( .A(n592), .ZN(n521) );
  XNOR2_X1 U474 ( .A(n376), .B(n377), .ZN(n673) );
  OR2_X2 U475 ( .A1(n628), .A2(KEYINPUT44), .ZN(n529) );
  XNOR2_X1 U476 ( .A(n417), .B(G104), .ZN(n506) );
  XNOR2_X1 U477 ( .A(n413), .B(n419), .ZN(n485) );
  XNOR2_X1 U478 ( .A(n418), .B(KEYINPUT3), .ZN(n413) );
  XNOR2_X1 U479 ( .A(n506), .B(n415), .ZN(n414) );
  BUF_X1 U480 ( .A(n506), .Z(n507) );
  BUF_X1 U481 ( .A(n485), .Z(n372) );
  BUF_X1 U482 ( .A(n731), .Z(n373) );
  XNOR2_X1 U483 ( .A(n414), .B(n485), .ZN(n731) );
  INV_X1 U484 ( .A(n724), .ZN(n393) );
  NAND2_X1 U485 ( .A1(n395), .A2(n390), .ZN(n389) );
  NAND2_X1 U486 ( .A1(n393), .A2(n394), .ZN(n395) );
  NAND2_X1 U487 ( .A1(n675), .A2(n674), .ZN(n679) );
  NOR2_X2 U488 ( .A1(n548), .A2(n547), .ZN(n375) );
  XNOR2_X1 U489 ( .A(n396), .B(KEYINPUT81), .ZN(n394) );
  XOR2_X1 U490 ( .A(n522), .B(KEYINPUT33), .Z(n377) );
  BUF_X1 U491 ( .A(n560), .Z(n604) );
  AND2_X2 U492 ( .A1(n397), .A2(n395), .ZN(n643) );
  NOR2_X1 U493 ( .A1(n753), .A2(n408), .ZN(n407) );
  NAND2_X1 U494 ( .A1(n388), .A2(n369), .ZN(n397) );
  NAND2_X1 U495 ( .A1(n387), .A2(n345), .ZN(n388) );
  AND2_X2 U496 ( .A1(n628), .A2(KEYINPUT44), .ZN(n547) );
  XNOR2_X2 U497 ( .A(n527), .B(KEYINPUT35), .ZN(n628) );
  NAND2_X1 U498 ( .A1(n385), .A2(n384), .ZN(n387) );
  NAND2_X1 U499 ( .A1(n612), .A2(n371), .ZN(n384) );
  NAND2_X1 U500 ( .A1(n386), .A2(n368), .ZN(n385) );
  INV_X1 U501 ( .A(n612), .ZN(n386) );
  NAND2_X1 U502 ( .A1(n345), .A2(KEYINPUT2), .ZN(n396) );
  XNOR2_X1 U503 ( .A(n398), .B(KEYINPUT84), .ZN(n531) );
  NOR2_X2 U504 ( .A1(n641), .A2(n656), .ZN(n642) );
  NOR2_X2 U505 ( .A1(n647), .A2(n656), .ZN(n649) );
  NOR2_X2 U506 ( .A1(n635), .A2(n656), .ZN(n636) );
  NAND2_X1 U507 ( .A1(n402), .A2(n401), .ZN(n406) );
  NAND2_X1 U508 ( .A1(n751), .A2(n403), .ZN(n402) );
  INV_X1 U509 ( .A(n753), .ZN(n403) );
  NAND2_X1 U510 ( .A1(n406), .A2(n404), .ZN(n599) );
  NAND2_X1 U511 ( .A1(n407), .A2(n405), .ZN(n404) );
  AND2_X1 U512 ( .A1(n365), .A2(n751), .ZN(n405) );
  INV_X1 U513 ( .A(KEYINPUT46), .ZN(n408) );
  NAND2_X1 U514 ( .A1(n613), .A2(n501), .ZN(n410) );
  AND2_X1 U515 ( .A1(n662), .A2(n409), .ZN(n582) );
  XNOR2_X2 U516 ( .A(KEYINPUT72), .B(KEYINPUT16), .ZN(n416) );
  XNOR2_X2 U517 ( .A(G110), .B(G107), .ZN(n417) );
  XNOR2_X2 U518 ( .A(G113), .B(KEYINPUT89), .ZN(n418) );
  NAND2_X1 U519 ( .A1(n560), .A2(n438), .ZN(n423) );
  BUF_X1 U520 ( .A(n621), .Z(n623) );
  XNOR2_X1 U521 ( .A(n618), .B(n617), .ZN(n619) );
  XNOR2_X1 U522 ( .A(n614), .B(n613), .ZN(n616) );
  BUF_X1 U523 ( .A(n643), .Z(n650) );
  NOR2_X1 U524 ( .A1(n703), .A2(n607), .ZN(n573) );
  INV_X1 U525 ( .A(n656), .ZN(n615) );
  INV_X1 U526 ( .A(n751), .ZN(n752) );
  NAND2_X1 U527 ( .A1(n742), .A2(G224), .ZN(n425) );
  XNOR2_X1 U528 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U529 ( .A(n427), .B(n458), .ZN(n428) );
  XNOR2_X1 U530 ( .A(n731), .B(n428), .ZN(n432) );
  XNOR2_X2 U531 ( .A(KEYINPUT77), .B(G143), .ZN(n430) );
  XNOR2_X2 U532 ( .A(n430), .B(n429), .ZN(n449) );
  XNOR2_X2 U533 ( .A(n449), .B(KEYINPUT4), .ZN(n739) );
  XNOR2_X1 U534 ( .A(KEYINPUT65), .B(G101), .ZN(n431) );
  XNOR2_X2 U535 ( .A(n739), .B(n431), .ZN(n480) );
  XNOR2_X1 U536 ( .A(n432), .B(n480), .ZN(n629) );
  INV_X1 U537 ( .A(n552), .ZN(n610) );
  OR2_X2 U538 ( .A1(n629), .A2(n610), .ZN(n436) );
  INV_X1 U539 ( .A(G902), .ZN(n501) );
  INV_X1 U540 ( .A(G237), .ZN(n433) );
  NAND2_X1 U541 ( .A1(n501), .A2(n433), .ZN(n437) );
  NAND2_X1 U542 ( .A1(n437), .A2(G210), .ZN(n434) );
  XNOR2_X2 U543 ( .A(n436), .B(n435), .ZN(n560) );
  NAND2_X1 U544 ( .A1(n437), .A2(G214), .ZN(n674) );
  INV_X1 U545 ( .A(KEYINPUT86), .ZN(n438) );
  XNOR2_X1 U546 ( .A(G898), .B(KEYINPUT91), .ZN(n727) );
  NAND2_X1 U547 ( .A1(n727), .A2(G953), .ZN(n439) );
  XNOR2_X1 U548 ( .A(n439), .B(KEYINPUT92), .ZN(n732) );
  NAND2_X1 U549 ( .A1(G234), .A2(G237), .ZN(n440) );
  XNOR2_X1 U550 ( .A(n440), .B(KEYINPUT14), .ZN(n441) );
  NAND2_X1 U551 ( .A1(G902), .A2(n441), .ZN(n553) );
  NOR2_X1 U552 ( .A1(n732), .A2(n553), .ZN(n442) );
  NAND2_X1 U553 ( .A1(G952), .A2(n441), .ZN(n691) );
  NOR2_X1 U554 ( .A1(n691), .A2(G953), .ZN(n556) );
  XNOR2_X1 U555 ( .A(G116), .B(n383), .ZN(n444) );
  XNOR2_X1 U556 ( .A(n444), .B(KEYINPUT7), .ZN(n448) );
  XOR2_X1 U557 ( .A(KEYINPUT9), .B(KEYINPUT101), .Z(n446) );
  XNOR2_X1 U558 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U559 ( .A(n448), .B(n447), .Z(n452) );
  NAND2_X1 U560 ( .A1(G217), .A2(n496), .ZN(n450) );
  XNOR2_X1 U561 ( .A(n449), .B(n450), .ZN(n451) );
  XNOR2_X1 U562 ( .A(n452), .B(n451), .ZN(n617) );
  NAND2_X1 U563 ( .A1(n617), .A2(n501), .ZN(n455) );
  INV_X1 U564 ( .A(KEYINPUT102), .ZN(n453) );
  XNOR2_X1 U565 ( .A(n453), .B(G478), .ZN(n454) );
  XNOR2_X1 U566 ( .A(n455), .B(n454), .ZN(n542) );
  INV_X1 U567 ( .A(n542), .ZN(n525) );
  XOR2_X1 U568 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n457) );
  NOR2_X1 U569 ( .A1(G953), .A2(G237), .ZN(n482) );
  NAND2_X1 U570 ( .A1(G214), .A2(n482), .ZN(n456) );
  XNOR2_X1 U571 ( .A(n457), .B(n456), .ZN(n459) );
  XNOR2_X1 U572 ( .A(n458), .B(KEYINPUT10), .ZN(n499) );
  XNOR2_X1 U573 ( .A(n459), .B(n499), .ZN(n467) );
  XNOR2_X1 U574 ( .A(n461), .B(n460), .ZN(n465) );
  XOR2_X1 U575 ( .A(KEYINPUT97), .B(KEYINPUT11), .Z(n463) );
  XNOR2_X1 U576 ( .A(n379), .B(G140), .ZN(n462) );
  XNOR2_X1 U577 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U578 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U579 ( .A(n467), .B(n466), .ZN(n638) );
  NAND2_X1 U580 ( .A1(n638), .A2(n501), .ZN(n470) );
  XOR2_X1 U581 ( .A(G475), .B(KEYINPUT99), .Z(n468) );
  XOR2_X1 U582 ( .A(KEYINPUT13), .B(n468), .Z(n469) );
  XNOR2_X1 U583 ( .A(n470), .B(n469), .ZN(n540) );
  OR2_X1 U584 ( .A1(n525), .A2(n540), .ZN(n677) );
  NAND2_X1 U585 ( .A1(n552), .A2(G234), .ZN(n471) );
  XNOR2_X1 U586 ( .A(n471), .B(KEYINPUT20), .ZN(n502) );
  AND2_X1 U587 ( .A1(n502), .A2(G221), .ZN(n472) );
  XNOR2_X1 U588 ( .A(n472), .B(KEYINPUT21), .ZN(n663) );
  INV_X1 U589 ( .A(n663), .ZN(n520) );
  NOR2_X1 U590 ( .A1(n677), .A2(n520), .ZN(n473) );
  NAND2_X1 U591 ( .A1(n538), .A2(n473), .ZN(n477) );
  XNOR2_X1 U592 ( .A(KEYINPUT71), .B(KEYINPUT22), .ZN(n475) );
  INV_X1 U593 ( .A(KEYINPUT70), .ZN(n474) );
  XNOR2_X1 U594 ( .A(n478), .B(KEYINPUT68), .ZN(n737) );
  XNOR2_X1 U595 ( .A(n737), .B(G146), .ZN(n479) );
  XNOR2_X2 U596 ( .A(n480), .B(n479), .ZN(n512) );
  XNOR2_X1 U597 ( .A(G137), .B(KEYINPUT5), .ZN(n481) );
  XNOR2_X1 U598 ( .A(n481), .B(KEYINPUT74), .ZN(n484) );
  NAND2_X1 U599 ( .A1(n482), .A2(G210), .ZN(n483) );
  XNOR2_X1 U600 ( .A(n484), .B(n483), .ZN(n486) );
  XNOR2_X1 U601 ( .A(n372), .B(n486), .ZN(n487) );
  XNOR2_X1 U602 ( .A(n512), .B(n487), .ZN(n644) );
  XNOR2_X2 U603 ( .A(n488), .B(G472), .ZN(n661) );
  XNOR2_X1 U604 ( .A(KEYINPUT104), .B(KEYINPUT6), .ZN(n489) );
  XNOR2_X1 U605 ( .A(n583), .B(KEYINPUT76), .ZN(n515) );
  XOR2_X1 U606 ( .A(KEYINPUT93), .B(G110), .Z(n491) );
  XNOR2_X1 U607 ( .A(n491), .B(n490), .ZN(n495) );
  XOR2_X1 U608 ( .A(KEYINPUT94), .B(KEYINPUT23), .Z(n493) );
  XNOR2_X1 U609 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U610 ( .A(n495), .B(n494), .Z(n498) );
  NAND2_X1 U611 ( .A1(G221), .A2(n496), .ZN(n497) );
  XNOR2_X1 U612 ( .A(n498), .B(n497), .ZN(n500) );
  XOR2_X1 U613 ( .A(G137), .B(G140), .Z(n509) );
  XNOR2_X1 U614 ( .A(n509), .B(n499), .ZN(n741) );
  XNOR2_X1 U615 ( .A(n500), .B(n741), .ZN(n613) );
  XOR2_X1 U616 ( .A(KEYINPUT95), .B(KEYINPUT25), .Z(n504) );
  NAND2_X1 U617 ( .A1(G217), .A2(n502), .ZN(n503) );
  XNOR2_X1 U618 ( .A(n504), .B(n503), .ZN(n505) );
  NAND2_X1 U619 ( .A1(G227), .A2(n742), .ZN(n508) );
  XOR2_X1 U620 ( .A(n508), .B(n507), .Z(n510) );
  XNOR2_X1 U621 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X2 U622 ( .A(n513), .B(G469), .ZN(n536) );
  XNOR2_X2 U623 ( .A(n536), .B(KEYINPUT1), .ZN(n592) );
  AND2_X1 U624 ( .A1(n662), .A2(n658), .ZN(n514) );
  XNOR2_X1 U625 ( .A(KEYINPUT75), .B(KEYINPUT32), .ZN(n516) );
  NAND2_X1 U626 ( .A1(n662), .A2(n592), .ZN(n517) );
  NOR2_X1 U627 ( .A1(n382), .A2(n517), .ZN(n518) );
  NAND2_X1 U628 ( .A1(n424), .A2(n521), .ZN(n532) );
  INV_X1 U629 ( .A(KEYINPUT105), .ZN(n522) );
  NAND2_X1 U630 ( .A1(n538), .A2(n673), .ZN(n524) );
  XNOR2_X1 U631 ( .A(n524), .B(n523), .ZN(n526) );
  AND2_X1 U632 ( .A1(n525), .A2(n540), .ZN(n577) );
  NAND2_X1 U633 ( .A1(n526), .A2(n577), .ZN(n527) );
  INV_X1 U634 ( .A(KEYINPUT66), .ZN(n528) );
  XNOR2_X1 U635 ( .A(n529), .B(n528), .ZN(n530) );
  INV_X1 U636 ( .A(n532), .ZN(n533) );
  NAND2_X1 U637 ( .A1(n382), .A2(n533), .ZN(n668) );
  INV_X1 U638 ( .A(n668), .ZN(n534) );
  NAND2_X1 U639 ( .A1(n538), .A2(n534), .ZN(n535) );
  INV_X1 U640 ( .A(n536), .ZN(n558) );
  NOR2_X1 U641 ( .A1(n382), .A2(n566), .ZN(n537) );
  AND2_X1 U642 ( .A1(n538), .A2(n537), .ZN(n702) );
  XNOR2_X1 U643 ( .A(n540), .B(KEYINPUT100), .ZN(n543) );
  OR2_X1 U644 ( .A1(n543), .A2(n542), .ZN(n705) );
  INV_X1 U645 ( .A(KEYINPUT103), .ZN(n541) );
  XNOR2_X1 U646 ( .A(n705), .B(n541), .ZN(n606) );
  NAND2_X1 U647 ( .A1(n543), .A2(n542), .ZN(n703) );
  NOR2_X1 U648 ( .A1(n662), .A2(n658), .ZN(n544) );
  OR2_X1 U649 ( .A1(n742), .A2(n553), .ZN(n554) );
  NOR2_X1 U650 ( .A1(G900), .A2(n554), .ZN(n555) );
  NOR2_X1 U651 ( .A1(n556), .A2(n555), .ZN(n570) );
  AND2_X1 U652 ( .A1(n661), .A2(n582), .ZN(n557) );
  XNOR2_X1 U653 ( .A(KEYINPUT28), .B(n557), .ZN(n559) );
  NAND2_X1 U654 ( .A1(n559), .A2(n558), .ZN(n576) );
  INV_X1 U655 ( .A(n576), .ZN(n563) );
  NAND2_X1 U656 ( .A1(n563), .A2(n694), .ZN(n565) );
  XOR2_X1 U657 ( .A(KEYINPUT42), .B(KEYINPUT108), .Z(n564) );
  INV_X1 U658 ( .A(n566), .ZN(n569) );
  NAND2_X1 U659 ( .A1(n661), .A2(n674), .ZN(n567) );
  XOR2_X1 U660 ( .A(KEYINPUT30), .B(n567), .Z(n568) );
  NAND2_X1 U661 ( .A1(n580), .A2(n675), .ZN(n572) );
  XOR2_X1 U662 ( .A(KEYINPUT82), .B(KEYINPUT39), .Z(n571) );
  XNOR2_X1 U663 ( .A(n572), .B(n571), .ZN(n607) );
  XNOR2_X1 U664 ( .A(n573), .B(KEYINPUT40), .ZN(n753) );
  BUF_X1 U665 ( .A(n574), .Z(n575) );
  NAND2_X1 U666 ( .A1(n717), .A2(n678), .ZN(n594) );
  NAND2_X1 U667 ( .A1(KEYINPUT47), .A2(n594), .ZN(n581) );
  INV_X1 U668 ( .A(n577), .ZN(n578) );
  NOR2_X1 U669 ( .A1(n604), .A2(n578), .ZN(n579) );
  NAND2_X1 U670 ( .A1(n580), .A2(n579), .ZN(n715) );
  NOR2_X1 U671 ( .A1(n703), .A2(n583), .ZN(n584) );
  NAND2_X1 U672 ( .A1(n582), .A2(n584), .ZN(n585) );
  XNOR2_X1 U673 ( .A(KEYINPUT106), .B(n585), .ZN(n600) );
  BUF_X1 U674 ( .A(n586), .Z(n587) );
  INV_X1 U675 ( .A(n587), .ZN(n588) );
  NOR2_X1 U676 ( .A1(n600), .A2(n588), .ZN(n590) );
  XNOR2_X1 U677 ( .A(KEYINPUT36), .B(KEYINPUT85), .ZN(n589) );
  XNOR2_X1 U678 ( .A(n590), .B(n589), .ZN(n591) );
  NOR2_X1 U679 ( .A1(n592), .A2(n591), .ZN(n720) );
  INV_X1 U680 ( .A(n720), .ZN(n597) );
  XOR2_X1 U681 ( .A(KEYINPUT47), .B(KEYINPUT67), .Z(n593) );
  NOR2_X1 U682 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U683 ( .A(KEYINPUT73), .B(n595), .ZN(n596) );
  AND2_X1 U684 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U685 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n603) );
  NOR2_X1 U686 ( .A1(n600), .A2(n658), .ZN(n601) );
  NAND2_X1 U687 ( .A1(n601), .A2(n674), .ZN(n602) );
  XNOR2_X1 U688 ( .A(n603), .B(n602), .ZN(n605) );
  AND2_X1 U689 ( .A1(n605), .A2(n604), .ZN(n620) );
  NOR2_X1 U690 ( .A1(n607), .A2(n606), .ZN(n723) );
  NOR2_X1 U691 ( .A1(n620), .A2(n723), .ZN(n608) );
  NAND2_X1 U692 ( .A1(n609), .A2(n608), .ZN(n611) );
  INV_X1 U693 ( .A(n612), .ZN(n724) );
  NAND2_X1 U694 ( .A1(n650), .A2(G217), .ZN(n614) );
  AND2_X1 U695 ( .A1(n616), .A2(n615), .ZN(G66) );
  NAND2_X1 U696 ( .A1(n650), .A2(G478), .ZN(n618) );
  AND2_X1 U697 ( .A1(n619), .A2(n615), .ZN(G63) );
  XOR2_X1 U698 ( .A(n620), .B(G140), .Z(G42) );
  INV_X1 U699 ( .A(n703), .ZN(n716) );
  NAND2_X1 U700 ( .A1(n623), .A2(n716), .ZN(n622) );
  XNOR2_X1 U701 ( .A(n622), .B(G113), .ZN(G15) );
  INV_X1 U702 ( .A(n705), .ZN(n710) );
  NAND2_X1 U703 ( .A1(n623), .A2(n710), .ZN(n624) );
  XNOR2_X1 U704 ( .A(n624), .B(G116), .ZN(G18) );
  XNOR2_X1 U705 ( .A(n625), .B(G101), .ZN(G3) );
  XOR2_X1 U706 ( .A(G110), .B(n626), .Z(G12) );
  XOR2_X1 U707 ( .A(n627), .B(G119), .Z(G21) );
  XOR2_X1 U708 ( .A(n628), .B(G122), .Z(G24) );
  NAND2_X1 U709 ( .A1(n643), .A2(G210), .ZN(n634) );
  BUF_X1 U710 ( .A(n629), .Z(n630) );
  XNOR2_X1 U711 ( .A(KEYINPUT87), .B(KEYINPUT54), .ZN(n631) );
  XNOR2_X1 U712 ( .A(n631), .B(KEYINPUT55), .ZN(n632) );
  XNOR2_X1 U713 ( .A(n634), .B(n633), .ZN(n635) );
  XNOR2_X1 U714 ( .A(n636), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U715 ( .A1(n643), .A2(G475), .ZN(n640) );
  XNOR2_X1 U716 ( .A(KEYINPUT88), .B(KEYINPUT59), .ZN(n637) );
  XNOR2_X1 U717 ( .A(n640), .B(n639), .ZN(n641) );
  XNOR2_X1 U718 ( .A(n642), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U719 ( .A1(n643), .A2(G472), .ZN(n646) );
  XNOR2_X1 U720 ( .A(n646), .B(n645), .ZN(n647) );
  INV_X1 U721 ( .A(KEYINPUT63), .ZN(n648) );
  XNOR2_X1 U722 ( .A(n649), .B(n648), .ZN(G57) );
  NAND2_X1 U723 ( .A1(n650), .A2(G469), .ZN(n655) );
  XNOR2_X1 U724 ( .A(KEYINPUT121), .B(KEYINPUT57), .ZN(n651) );
  XNOR2_X1 U725 ( .A(n651), .B(KEYINPUT58), .ZN(n652) );
  XNOR2_X1 U726 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U727 ( .A(n655), .B(n654), .ZN(n657) );
  NOR2_X1 U728 ( .A1(n657), .A2(n656), .ZN(G54) );
  XOR2_X1 U729 ( .A(KEYINPUT51), .B(KEYINPUT114), .Z(n671) );
  NOR2_X1 U730 ( .A1(n424), .A2(n658), .ZN(n659) );
  XNOR2_X1 U731 ( .A(n659), .B(KEYINPUT50), .ZN(n660) );
  NOR2_X1 U732 ( .A1(n382), .A2(n660), .ZN(n667) );
  INV_X1 U733 ( .A(n662), .ZN(n664) );
  NOR2_X1 U734 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U735 ( .A(n665), .B(KEYINPUT49), .ZN(n666) );
  NAND2_X1 U736 ( .A1(n667), .A2(n666), .ZN(n669) );
  NAND2_X1 U737 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U738 ( .A(n671), .B(n670), .ZN(n672) );
  NAND2_X1 U739 ( .A1(n672), .A2(n694), .ZN(n687) );
  NOR2_X1 U740 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U741 ( .A1(n677), .A2(n676), .ZN(n682) );
  NOR2_X1 U742 ( .A1(n346), .A2(n679), .ZN(n680) );
  XOR2_X1 U743 ( .A(KEYINPUT115), .B(n680), .Z(n681) );
  NOR2_X1 U744 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U745 ( .A(KEYINPUT116), .B(n683), .Z(n684) );
  NAND2_X1 U746 ( .A1(n693), .A2(n684), .ZN(n685) );
  XOR2_X1 U747 ( .A(KEYINPUT117), .B(n685), .Z(n686) );
  NAND2_X1 U748 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U749 ( .A(n688), .B(KEYINPUT52), .ZN(n689) );
  XOR2_X1 U750 ( .A(KEYINPUT118), .B(n689), .Z(n690) );
  NOR2_X1 U751 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U752 ( .A(KEYINPUT119), .B(n692), .Z(n697) );
  NAND2_X1 U753 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U754 ( .A1(n695), .A2(n742), .ZN(n696) );
  NOR2_X1 U755 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U756 ( .A1(n699), .A2(n698), .ZN(n701) );
  XOR2_X1 U757 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n700) );
  XNOR2_X1 U758 ( .A(n701), .B(n700), .ZN(G75) );
  INV_X1 U759 ( .A(n702), .ZN(n706) );
  NOR2_X1 U760 ( .A1(n706), .A2(n703), .ZN(n704) );
  XOR2_X1 U761 ( .A(G104), .B(n704), .Z(G6) );
  NOR2_X1 U762 ( .A1(n706), .A2(n705), .ZN(n708) );
  XNOR2_X1 U763 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n707) );
  XNOR2_X1 U764 ( .A(n708), .B(n707), .ZN(n709) );
  XNOR2_X1 U765 ( .A(n383), .B(n709), .ZN(G9) );
  XOR2_X1 U766 ( .A(KEYINPUT111), .B(KEYINPUT29), .Z(n712) );
  NAND2_X1 U767 ( .A1(n717), .A2(n710), .ZN(n711) );
  XNOR2_X1 U768 ( .A(n712), .B(n711), .ZN(n714) );
  XOR2_X1 U769 ( .A(G128), .B(KEYINPUT110), .Z(n713) );
  XNOR2_X1 U770 ( .A(n714), .B(n713), .ZN(G30) );
  XNOR2_X1 U771 ( .A(n379), .B(n715), .ZN(G45) );
  XNOR2_X1 U772 ( .A(G146), .B(KEYINPUT112), .ZN(n719) );
  NAND2_X1 U773 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U774 ( .A(n719), .B(n718), .ZN(G48) );
  XOR2_X1 U775 ( .A(KEYINPUT37), .B(KEYINPUT113), .Z(n722) );
  XNOR2_X1 U776 ( .A(G125), .B(n720), .ZN(n721) );
  XNOR2_X1 U777 ( .A(n722), .B(n721), .ZN(G27) );
  XOR2_X1 U778 ( .A(G134), .B(n723), .Z(G36) );
  NOR2_X1 U779 ( .A1(n724), .A2(G953), .ZN(n730) );
  XOR2_X1 U780 ( .A(KEYINPUT122), .B(KEYINPUT61), .Z(n726) );
  NAND2_X1 U781 ( .A1(G224), .A2(G953), .ZN(n725) );
  XNOR2_X1 U782 ( .A(n726), .B(n725), .ZN(n728) );
  NOR2_X1 U783 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X1 U784 ( .A1(n730), .A2(n729), .ZN(n736) );
  XNOR2_X1 U785 ( .A(n373), .B(G101), .ZN(n733) );
  NAND2_X1 U786 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U787 ( .A(n734), .B(KEYINPUT123), .ZN(n735) );
  XOR2_X1 U788 ( .A(n736), .B(n735), .Z(G69) );
  XNOR2_X1 U789 ( .A(n737), .B(KEYINPUT124), .ZN(n738) );
  XNOR2_X1 U790 ( .A(n739), .B(n738), .ZN(n740) );
  XOR2_X1 U791 ( .A(n741), .B(n740), .Z(n744) );
  XOR2_X1 U792 ( .A(n611), .B(n744), .Z(n743) );
  NAND2_X1 U793 ( .A1(n743), .A2(n742), .ZN(n750) );
  XNOR2_X1 U794 ( .A(n744), .B(G227), .ZN(n745) );
  XNOR2_X1 U795 ( .A(n745), .B(KEYINPUT125), .ZN(n746) );
  NAND2_X1 U796 ( .A1(n746), .A2(G900), .ZN(n747) );
  XNOR2_X1 U797 ( .A(KEYINPUT126), .B(n747), .ZN(n748) );
  NAND2_X1 U798 ( .A1(n748), .A2(G953), .ZN(n749) );
  NAND2_X1 U799 ( .A1(n750), .A2(n749), .ZN(G72) );
  XOR2_X1 U800 ( .A(G137), .B(n752), .Z(G39) );
  XOR2_X1 U801 ( .A(G131), .B(n753), .Z(G33) );
endmodule

