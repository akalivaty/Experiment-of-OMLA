//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 0 0 1 0 0 0 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 0 1 0 1 0 1 0 0 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 1 1 0 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n809, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1051, new_n1052;
  INV_X1    g000(.A(KEYINPUT96), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n204));
  INV_X1    g003(.A(G22gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G15gat), .ZN(new_n206));
  INV_X1    g005(.A(G15gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G22gat), .ZN(new_n208));
  AND3_X1   g007(.A1(new_n206), .A2(new_n208), .A3(KEYINPUT86), .ZN(new_n209));
  AOI21_X1  g008(.A(KEYINPUT86), .B1(new_n206), .B2(new_n208), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n204), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n206), .A2(new_n208), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT86), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n206), .A2(new_n208), .A3(KEYINPUT86), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n214), .A2(new_n203), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT87), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n211), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n219), .A3(G8gat), .ZN(new_n220));
  INV_X1    g019(.A(G8gat), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n211), .B(new_n216), .C1(new_n218), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G57gat), .B(G64gat), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT89), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G71gat), .B(G78gat), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  OAI211_X1 g028(.A(KEYINPUT89), .B(new_n227), .C1(new_n224), .C2(new_n225), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n223), .B1(KEYINPUT21), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT91), .B(KEYINPUT20), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n232), .B(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G127gat), .B(G155gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(G231gat), .A2(G233gat), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n238), .B1(new_n231), .B2(KEYINPUT21), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NOR3_X1   g039(.A1(new_n231), .A2(KEYINPUT21), .A3(new_n238), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NOR3_X1   g042(.A1(new_n240), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  OR3_X1    g043(.A1(new_n231), .A2(KEYINPUT21), .A3(new_n238), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n242), .B1(new_n245), .B2(new_n239), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n236), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(G183gat), .B(G211gat), .Z(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n243), .B1(new_n240), .B2(new_n241), .ZN(new_n250));
  INV_X1    g049(.A(new_n236), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n245), .A2(new_n239), .A3(new_n242), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n247), .A2(new_n249), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n249), .B1(new_n247), .B2(new_n253), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n235), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n247), .A2(new_n253), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(new_n248), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n247), .A2(new_n249), .A3(new_n253), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(new_n234), .A3(new_n259), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(KEYINPUT94), .B(KEYINPUT95), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT7), .ZN(new_n264));
  OAI211_X1 g063(.A(G85gat), .B(G92gat), .C1(new_n264), .C2(KEYINPUT92), .ZN(new_n265));
  NAND2_X1  g064(.A1(G85gat), .A2(G92gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT92), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(new_n267), .A3(KEYINPUT7), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(KEYINPUT93), .A2(G85gat), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(G92gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(KEYINPUT93), .A2(G85gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(G99gat), .A2(G106gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT8), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n269), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G99gat), .ZN(new_n278));
  INV_X1    g077(.A(G106gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n277), .A2(new_n275), .A3(new_n280), .ZN(new_n281));
  AND2_X1   g080(.A1(KEYINPUT93), .A2(G85gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n282), .A2(new_n270), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n283), .A2(new_n272), .B1(KEYINPUT8), .B2(new_n275), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n280), .A2(new_n275), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n284), .A2(new_n285), .A3(new_n269), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT85), .ZN(new_n288));
  INV_X1    g087(.A(G43gat), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n288), .B1(new_n289), .B2(G50gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT15), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT14), .ZN(new_n293));
  INV_X1    g092(.A(G29gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n296));
  AOI21_X1  g095(.A(G36gat), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n294), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n292), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(G43gat), .B(G50gat), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n297), .A2(new_n299), .ZN(new_n303));
  AOI22_X1  g102(.A1(new_n300), .A2(new_n302), .B1(new_n303), .B2(new_n291), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n292), .B(new_n301), .C1(new_n297), .C2(new_n299), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT17), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G36gat), .ZN(new_n307));
  AND2_X1   g106(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n310), .A2(new_n291), .A3(new_n298), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n310), .A2(new_n298), .B1(new_n291), .B2(new_n290), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n311), .B1(new_n312), .B2(new_n301), .ZN(new_n313));
  INV_X1    g112(.A(new_n305), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT17), .ZN(new_n315));
  NOR3_X1   g114(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n287), .B1(new_n306), .B2(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n313), .A2(new_n314), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n285), .B1(new_n284), .B2(new_n269), .ZN(new_n319));
  AND4_X1   g118(.A1(new_n285), .A2(new_n269), .A3(new_n274), .A4(new_n276), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AND2_X1   g120(.A1(G232gat), .A2(G233gat), .ZN(new_n322));
  AOI22_X1  g121(.A1(new_n318), .A2(new_n321), .B1(KEYINPUT41), .B2(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(KEYINPUT41), .ZN(new_n324));
  XNOR2_X1  g123(.A(G134gat), .B(G162gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n317), .A2(new_n323), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n326), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n304), .A2(KEYINPUT17), .A3(new_n305), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n315), .B1(new_n313), .B2(new_n314), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n321), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n322), .A2(KEYINPUT41), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n304), .A2(new_n305), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n332), .B1(new_n333), .B2(new_n287), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n328), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G190gat), .B(G218gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  AND3_X1   g136(.A1(new_n327), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n337), .B1(new_n327), .B2(new_n335), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n263), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n327), .A2(new_n335), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(new_n336), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n327), .A2(new_n335), .A3(new_n337), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n342), .A2(new_n262), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n202), .B1(new_n261), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n345), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n256), .A2(new_n260), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(new_n348), .A3(KEYINPUT96), .ZN(new_n349));
  AND2_X1   g148(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G230gat), .A2(G233gat), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n229), .B(new_n230), .C1(new_n319), .C2(new_n320), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n231), .A2(new_n281), .A3(new_n286), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT10), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n321), .A2(KEYINPUT10), .A3(new_n231), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n352), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n353), .A2(new_n354), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n358), .B1(new_n359), .B2(new_n352), .ZN(new_n360));
  XNOR2_X1  g159(.A(G120gat), .B(G148gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(G176gat), .B(G204gat), .ZN(new_n362));
  XOR2_X1   g161(.A(new_n361), .B(new_n362), .Z(new_n363));
  OR2_X1    g162(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n356), .A2(new_n357), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n351), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n359), .A2(new_n352), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(new_n367), .A3(new_n363), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n364), .A2(KEYINPUT97), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT97), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n360), .A2(new_n363), .ZN(new_n371));
  INV_X1    g170(.A(new_n368), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n350), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT78), .ZN(new_n376));
  NAND2_X1  g175(.A1(G228gat), .A2(G233gat), .ZN(new_n377));
  OR2_X1    g176(.A1(G155gat), .A2(G162gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(G155gat), .A2(G162gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(G141gat), .B(G148gat), .Z(new_n381));
  INV_X1    g180(.A(KEYINPUT2), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT75), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n378), .A2(new_n384), .A3(new_n379), .ZN(new_n385));
  AND2_X1   g184(.A1(G155gat), .A2(G162gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(G155gat), .A2(G162gat), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT75), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n381), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT76), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n390), .B1(new_n386), .B2(new_n382), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n379), .A2(KEYINPUT76), .A3(KEYINPUT2), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n383), .B1(new_n389), .B2(new_n393), .ZN(new_n394));
  XOR2_X1   g193(.A(G197gat), .B(G204gat), .Z(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(KEYINPUT72), .B(G211gat), .ZN(new_n397));
  INV_X1    g196(.A(G218gat), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n396), .B1(new_n399), .B2(KEYINPUT22), .ZN(new_n400));
  XNOR2_X1  g199(.A(G211gat), .B(G218gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT29), .ZN(new_n403));
  INV_X1    g202(.A(new_n401), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n396), .B(new_n404), .C1(new_n399), .C2(KEYINPUT22), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n402), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT3), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n394), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  XOR2_X1   g207(.A(KEYINPUT72), .B(G211gat), .Z(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(G218gat), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT22), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n395), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n404), .B1(new_n412), .B2(KEYINPUT73), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT73), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n400), .A2(new_n414), .A3(new_n401), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n393), .A2(new_n381), .A3(new_n385), .A4(new_n388), .ZN(new_n416));
  XNOR2_X1  g215(.A(G141gat), .B(G148gat), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n379), .B(new_n378), .C1(new_n417), .C2(KEYINPUT2), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n407), .A3(new_n418), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n413), .A2(new_n415), .B1(new_n419), .B2(new_n403), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n377), .B1(new_n408), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n413), .A2(new_n403), .A3(new_n415), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n394), .B1(new_n422), .B2(new_n407), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n400), .A2(new_n414), .A3(new_n401), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n401), .B1(new_n400), .B2(new_n414), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT29), .B1(new_n394), .B2(new_n407), .ZN(new_n427));
  OAI211_X1 g226(.A(G228gat), .B(G233gat), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n421), .B1(new_n423), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n376), .B1(new_n429), .B2(G22gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(G78gat), .B(G106gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(KEYINPUT31), .B(G50gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n421), .B(new_n205), .C1(new_n423), .C2(new_n428), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n420), .A2(new_n377), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT3), .B1(new_n426), .B2(new_n403), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n437), .B1(new_n438), .B2(new_n394), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n205), .B1(new_n439), .B2(new_n421), .ZN(new_n440));
  OAI22_X1  g239(.A1(new_n430), .A2(new_n434), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n429), .A2(G22gat), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n442), .A2(new_n376), .A3(new_n435), .A4(new_n433), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n381), .A2(new_n385), .A3(new_n388), .ZN(new_n445));
  INV_X1    g244(.A(new_n392), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT76), .B1(new_n379), .B2(KEYINPUT2), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n418), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT3), .ZN(new_n450));
  XOR2_X1   g249(.A(G127gat), .B(G134gat), .Z(new_n451));
  XNOR2_X1  g250(.A(G113gat), .B(G120gat), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n451), .B1(KEYINPUT1), .B2(new_n452), .ZN(new_n453));
  XOR2_X1   g252(.A(G113gat), .B(G120gat), .Z(new_n454));
  INV_X1    g253(.A(KEYINPUT1), .ZN(new_n455));
  XNOR2_X1  g254(.A(G127gat), .B(G134gat), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n450), .A2(new_n419), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT68), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n453), .A2(new_n457), .A3(KEYINPUT68), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n461), .A2(new_n394), .A3(KEYINPUT4), .A4(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(G225gat), .A2(G233gat), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT4), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n465), .B1(new_n449), .B2(new_n458), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n459), .A2(new_n463), .A3(new_n464), .A4(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT5), .ZN(new_n468));
  AND2_X1   g267(.A1(new_n453), .A2(new_n457), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n469), .A2(new_n418), .A3(new_n416), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n449), .A2(new_n458), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n464), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n468), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n467), .A2(new_n474), .ZN(new_n475));
  NOR3_X1   g274(.A1(new_n449), .A2(new_n458), .A3(new_n465), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n461), .A2(new_n394), .A3(new_n462), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n476), .B1(new_n477), .B2(new_n465), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n469), .B1(KEYINPUT3), .B2(new_n449), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n473), .B1(new_n479), .B2(new_n419), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(new_n480), .A3(new_n468), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n475), .A2(new_n481), .ZN(new_n482));
  XOR2_X1   g281(.A(G1gat), .B(G29gat), .Z(new_n483));
  XNOR2_X1  g282(.A(G57gat), .B(G85gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n483), .B(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n482), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT6), .ZN(new_n489));
  INV_X1    g288(.A(new_n487), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n475), .A2(new_n481), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n488), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n482), .A2(KEYINPUT6), .A3(new_n487), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(G226gat), .A2(G233gat), .ZN(new_n495));
  XOR2_X1   g294(.A(new_n495), .B(KEYINPUT74), .Z(new_n496));
  INV_X1    g295(.A(G183gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT27), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT27), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(G183gat), .ZN(new_n500));
  INV_X1    g299(.A(G190gat), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n498), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT67), .ZN(new_n503));
  XNOR2_X1  g302(.A(KEYINPUT27), .B(G183gat), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT67), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(new_n505), .A3(new_n501), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT66), .ZN(new_n508));
  OR2_X1    g307(.A1(new_n508), .A2(KEYINPUT28), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n508), .A2(KEYINPUT28), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n503), .A2(new_n506), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(G183gat), .A2(G190gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(G169gat), .A2(G176gat), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT26), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n513), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n517), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n510), .A2(new_n512), .A3(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT24), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n513), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n497), .A2(new_n501), .ZN(new_n523));
  NAND3_X1  g322(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT64), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n514), .A2(KEYINPUT23), .ZN(new_n527));
  NAND2_X1  g326(.A1(G169gat), .A2(G176gat), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT23), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n529), .B1(G169gat), .B2(G176gat), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT64), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n522), .A2(new_n523), .A3(new_n532), .A4(new_n524), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n526), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT25), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT65), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n513), .B1(new_n536), .B2(KEYINPUT24), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n521), .A2(KEYINPUT65), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n523), .B(new_n524), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  AND4_X1   g338(.A1(KEYINPUT25), .A2(new_n527), .A3(new_n528), .A4(new_n530), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n534), .A2(new_n535), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n496), .B1(new_n520), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n534), .A2(new_n535), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n540), .A2(new_n539), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n510), .A2(new_n512), .A3(new_n519), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT29), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n495), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n542), .B(new_n426), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n495), .B1(new_n545), .B2(new_n546), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n403), .B1(new_n520), .B2(new_n541), .ZN(new_n551));
  INV_X1    g350(.A(new_n496), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n549), .B1(new_n553), .B2(new_n426), .ZN(new_n554));
  XNOR2_X1  g353(.A(G8gat), .B(G36gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(G64gat), .B(G92gat), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n555), .B(new_n556), .Z(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n413), .A2(new_n415), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n546), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n496), .B1(new_n561), .B2(new_n403), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n560), .B1(new_n562), .B2(new_n550), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n563), .A2(new_n549), .A3(new_n557), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n559), .A2(KEYINPUT30), .A3(new_n564), .ZN(new_n565));
  OR3_X1    g364(.A1(new_n554), .A2(KEYINPUT30), .A3(new_n558), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n444), .B1(new_n494), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n477), .A2(new_n465), .ZN(new_n569));
  INV_X1    g368(.A(new_n476), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(new_n459), .A3(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(KEYINPUT79), .B(KEYINPUT39), .Z(new_n572));
  NAND3_X1  g371(.A1(new_n571), .A2(new_n473), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n464), .B1(new_n478), .B2(new_n459), .ZN(new_n574));
  OAI21_X1  g373(.A(KEYINPUT39), .B1(new_n472), .B2(new_n473), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n573), .B(new_n490), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT40), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n488), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n577), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT80), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n576), .A2(KEYINPUT80), .A3(new_n577), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n578), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n567), .ZN(new_n584));
  AOI22_X1  g383(.A1(new_n583), .A2(new_n584), .B1(new_n443), .B2(new_n441), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT37), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n548), .B1(new_n520), .B2(new_n541), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n587), .B(new_n426), .C1(new_n547), .C2(new_n496), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n586), .B1(new_n589), .B2(KEYINPUT81), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT81), .ZN(new_n591));
  AOI22_X1  g390(.A1(new_n551), .A2(new_n495), .B1(new_n561), .B2(new_n496), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n591), .B(new_n588), .C1(new_n592), .C2(new_n426), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT38), .B1(new_n590), .B2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT82), .B(KEYINPUT37), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n549), .B(new_n595), .C1(new_n553), .C2(new_n426), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT83), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT83), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n563), .A2(new_n598), .A3(new_n549), .A4(new_n595), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n594), .A2(new_n600), .A3(new_n558), .ZN(new_n601));
  AND3_X1   g400(.A1(new_n492), .A2(new_n493), .A3(new_n564), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n586), .B1(new_n563), .B2(new_n549), .ZN(new_n603));
  AOI211_X1 g402(.A(new_n557), .B(new_n603), .C1(new_n597), .C2(new_n599), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT38), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n601), .B(new_n602), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n568), .B1(new_n585), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT34), .ZN(new_n608));
  INV_X1    g407(.A(G227gat), .ZN(new_n609));
  INV_X1    g408(.A(G233gat), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n462), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT68), .B1(new_n453), .B2(new_n457), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n614), .B1(new_n520), .B2(new_n541), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n461), .A2(new_n462), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n616), .A2(new_n545), .A3(new_n546), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n611), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT69), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n608), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n611), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n616), .A2(new_n545), .A3(new_n546), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n616), .B1(new_n545), .B2(new_n546), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n619), .B(new_n621), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n624), .A2(KEYINPUT70), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT70), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n626), .B1(new_n618), .B2(new_n619), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n620), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n629));
  AOI21_X1  g428(.A(KEYINPUT34), .B1(new_n629), .B2(KEYINPUT69), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n618), .A2(new_n619), .A3(new_n626), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n624), .A2(KEYINPUT70), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n615), .A2(new_n611), .A3(new_n617), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(KEYINPUT32), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT33), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(G15gat), .B(G43gat), .Z(new_n639));
  XNOR2_X1  g438(.A(G71gat), .B(G99gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n636), .A2(new_n638), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n641), .ZN(new_n643));
  OAI211_X1 g442(.A(new_n635), .B(KEYINPUT32), .C1(new_n637), .C2(new_n643), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n634), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT36), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n642), .A2(new_n644), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n628), .A2(new_n648), .A3(new_n633), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n646), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(KEYINPUT71), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT71), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n628), .A2(new_n648), .A3(new_n633), .A4(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n651), .A2(new_n653), .A3(new_n646), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n650), .B1(KEYINPUT36), .B2(new_n654), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n651), .A2(new_n646), .A3(new_n444), .A4(new_n653), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n567), .A2(new_n494), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT35), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n657), .A2(KEYINPUT35), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n646), .A2(new_n649), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n659), .A2(new_n660), .A3(new_n444), .ZN(new_n661));
  AOI22_X1  g460(.A1(new_n607), .A2(new_n655), .B1(new_n658), .B2(new_n661), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n222), .B(new_n220), .C1(new_n306), .C2(new_n316), .ZN(new_n663));
  NAND2_X1  g462(.A1(G229gat), .A2(G233gat), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n223), .A2(new_n318), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT18), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n663), .A2(new_n665), .A3(KEYINPUT18), .A4(new_n664), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n664), .B(KEYINPUT13), .Z(new_n670));
  NOR2_X1   g469(.A1(new_n223), .A2(new_n318), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n333), .B1(new_n222), .B2(new_n220), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n668), .A2(new_n669), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT84), .ZN(new_n675));
  XNOR2_X1  g474(.A(G113gat), .B(G141gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(G197gat), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT11), .B(G169gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT12), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n674), .A2(new_n675), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n680), .B1(new_n674), .B2(new_n675), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(KEYINPUT88), .B1(new_n662), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n583), .A2(new_n584), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n606), .A2(new_n687), .A3(new_n444), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n654), .A2(KEYINPUT36), .ZN(new_n689));
  INV_X1    g488(.A(new_n650), .ZN(new_n690));
  INV_X1    g489(.A(new_n568), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n688), .A2(new_n689), .A3(new_n690), .A4(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n658), .A2(new_n661), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT88), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(new_n695), .A3(new_n684), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n375), .B1(new_n686), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n494), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(G1gat), .ZN(G1324gat));
  INV_X1    g499(.A(new_n375), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n695), .B1(new_n694), .B2(new_n684), .ZN(new_n702));
  AOI211_X1 g501(.A(KEYINPUT88), .B(new_n685), .C1(new_n692), .C2(new_n693), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n584), .B(new_n701), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT98), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT98), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n697), .A2(new_n706), .A3(new_n584), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n705), .A2(G8gat), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(KEYINPUT99), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT99), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n705), .A2(new_n707), .A3(new_n710), .A4(G8gat), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT42), .ZN(new_n713));
  XOR2_X1   g512(.A(KEYINPUT16), .B(G8gat), .Z(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n704), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n686), .A2(new_n696), .ZN(new_n717));
  AND4_X1   g516(.A1(new_n706), .A2(new_n717), .A3(new_n584), .A4(new_n701), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n706), .B1(new_n697), .B2(new_n584), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n714), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n716), .B1(new_n720), .B2(new_n713), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n712), .A2(new_n721), .ZN(G1325gat));
  NAND2_X1  g521(.A1(new_n717), .A2(new_n701), .ZN(new_n723));
  OAI21_X1  g522(.A(G15gat), .B1(new_n723), .B2(new_n655), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n697), .A2(new_n207), .A3(new_n660), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(G1326gat));
  OAI21_X1  g525(.A(KEYINPUT100), .B1(new_n723), .B2(new_n444), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT100), .ZN(new_n728));
  INV_X1    g527(.A(new_n444), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n697), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(KEYINPUT43), .B(G22gat), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n731), .B(new_n733), .ZN(G1327gat));
  INV_X1    g533(.A(new_n374), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n735), .A2(new_n348), .A3(new_n347), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n717), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n494), .A2(G29gat), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n737), .A2(KEYINPUT45), .A3(new_n738), .ZN(new_n739));
  XOR2_X1   g538(.A(new_n374), .B(KEYINPUT102), .Z(new_n740));
  XNOR2_X1  g539(.A(new_n348), .B(KEYINPUT101), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n740), .A2(new_n742), .A3(new_n685), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT103), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n345), .B(new_n744), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n662), .A2(KEYINPUT44), .A3(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n747), .B1(new_n694), .B2(new_n345), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n698), .B(new_n743), .C1(new_n746), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G29gat), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n717), .A2(new_n736), .ZN(new_n752));
  INV_X1    g551(.A(new_n738), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n750), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(KEYINPUT104), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT104), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n739), .A2(new_n757), .A3(new_n754), .A4(new_n750), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(G1328gat));
  NOR2_X1   g558(.A1(new_n746), .A2(new_n748), .ZN(new_n760));
  INV_X1    g559(.A(new_n743), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n584), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT105), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n762), .A2(KEYINPUT105), .A3(new_n584), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n765), .A2(G36gat), .A3(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n737), .A2(new_n307), .A3(new_n584), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(KEYINPUT46), .ZN(new_n769));
  OR2_X1    g568(.A1(new_n768), .A2(KEYINPUT46), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n767), .A2(new_n769), .A3(new_n770), .ZN(G1329gat));
  NAND3_X1  g570(.A1(new_n737), .A2(new_n289), .A3(new_n660), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n760), .A2(new_n655), .A3(new_n761), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n289), .B2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT47), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n772), .B(KEYINPUT47), .C1(new_n289), .C2(new_n773), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(G1330gat));
  INV_X1    g577(.A(G50gat), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n779), .B1(new_n762), .B2(new_n729), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT106), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT48), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n444), .A2(G50gat), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  OAI22_X1  g584(.A1(new_n752), .A2(new_n785), .B1(KEYINPUT106), .B2(KEYINPUT48), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n780), .A2(new_n783), .A3(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n783), .ZN(new_n788));
  OR2_X1    g587(.A1(new_n746), .A2(new_n748), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n789), .A2(new_n729), .A3(new_n743), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G50gat), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n737), .A2(new_n784), .B1(new_n781), .B2(new_n782), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n788), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n787), .A2(new_n793), .ZN(G1331gat));
  AND4_X1   g593(.A1(new_n694), .A2(new_n685), .A3(new_n350), .A4(new_n740), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n698), .ZN(new_n796));
  XNOR2_X1  g595(.A(KEYINPUT107), .B(G57gat), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n796), .B(new_n797), .ZN(G1332gat));
  NAND2_X1  g597(.A1(new_n795), .A2(new_n584), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n799), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n800));
  XOR2_X1   g599(.A(KEYINPUT49), .B(G64gat), .Z(new_n801));
  OAI21_X1  g600(.A(new_n800), .B1(new_n799), .B2(new_n801), .ZN(G1333gat));
  INV_X1    g601(.A(new_n655), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n795), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n660), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n805), .A2(G71gat), .ZN(new_n806));
  AOI22_X1  g605(.A1(new_n804), .A2(G71gat), .B1(new_n795), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g607(.A1(new_n795), .A2(new_n729), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g609(.A1(new_n662), .A2(new_n347), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n684), .A2(new_n348), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT51), .ZN(new_n814));
  OAI21_X1  g613(.A(KEYINPUT109), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT51), .B1(new_n811), .B2(new_n812), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  AND4_X1   g616(.A1(KEYINPUT51), .A2(new_n694), .A3(new_n345), .A4(new_n812), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT109), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n815), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n735), .A2(new_n698), .A3(new_n283), .ZN(new_n822));
  XOR2_X1   g621(.A(new_n822), .B(KEYINPUT110), .Z(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n812), .A2(new_n735), .ZN(new_n825));
  XOR2_X1   g624(.A(new_n825), .B(KEYINPUT108), .Z(new_n826));
  AND2_X1   g625(.A1(new_n789), .A2(new_n826), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n827), .A2(new_n698), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n824), .B1(new_n828), .B2(new_n283), .ZN(G1336gat));
  INV_X1    g628(.A(new_n740), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n830), .A2(G92gat), .A3(new_n567), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n821), .A2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n584), .B(new_n826), .C1(new_n746), .C2(new_n748), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(G92gat), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n832), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT111), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n831), .B1(new_n816), .B2(new_n818), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n837), .B1(new_n839), .B2(KEYINPUT52), .ZN(new_n840));
  AOI211_X1 g639(.A(KEYINPUT111), .B(new_n833), .C1(new_n835), .C2(new_n838), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n836), .B1(new_n840), .B2(new_n841), .ZN(G1337gat));
  NAND4_X1  g641(.A1(new_n821), .A2(new_n278), .A3(new_n660), .A4(new_n735), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n827), .A2(new_n803), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n843), .B1(new_n844), .B2(new_n278), .ZN(G1338gat));
  NAND3_X1  g644(.A1(new_n740), .A2(new_n279), .A3(new_n729), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(KEYINPUT112), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n821), .A2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n729), .B(new_n826), .C1(new_n746), .C2(new_n748), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(G106gat), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n848), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n847), .B1(new_n816), .B2(new_n818), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n853), .B1(new_n855), .B2(KEYINPUT53), .ZN(new_n856));
  AOI211_X1 g655(.A(KEYINPUT113), .B(new_n849), .C1(new_n851), .C2(new_n854), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n852), .B1(new_n856), .B2(new_n857), .ZN(G1339gat));
  AND4_X1   g657(.A1(new_n685), .A2(new_n346), .A3(new_n349), .A4(new_n374), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n356), .A2(new_n357), .A3(new_n352), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n366), .A2(KEYINPUT54), .A3(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n363), .B1(new_n358), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT55), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n861), .A2(KEYINPUT55), .A3(new_n863), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n368), .A3(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n668), .A2(new_n669), .A3(new_n673), .A4(new_n680), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n671), .A2(new_n672), .A3(new_n670), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n664), .B1(new_n663), .B2(new_n665), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n679), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n345), .B(KEYINPUT103), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n674), .A2(new_n675), .ZN(new_n879));
  INV_X1    g678(.A(new_n680), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n867), .A2(new_n368), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n881), .A2(new_n681), .A3(new_n866), .A4(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT114), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n874), .A2(new_n369), .A3(new_n373), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n745), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n884), .B1(new_n883), .B2(new_n885), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n878), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n859), .B1(new_n889), .B2(new_n741), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(new_n494), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n656), .A2(new_n584), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(new_n684), .A3(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(G113gat), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n584), .A2(new_n494), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  NOR4_X1   g695(.A1(new_n890), .A2(new_n805), .A3(new_n729), .A4(new_n896), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n685), .A2(new_n894), .ZN(new_n898));
  AOI22_X1  g697(.A1(new_n893), .A2(new_n894), .B1(new_n897), .B2(new_n898), .ZN(G1340gat));
  NAND3_X1  g698(.A1(new_n891), .A2(new_n735), .A3(new_n892), .ZN(new_n900));
  INV_X1    g699(.A(G120gat), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n830), .A2(new_n901), .ZN(new_n902));
  AOI22_X1  g701(.A1(new_n900), .A2(new_n901), .B1(new_n897), .B2(new_n902), .ZN(G1341gat));
  NAND2_X1  g702(.A1(new_n891), .A2(new_n892), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n904), .A2(G127gat), .A3(new_n261), .ZN(new_n905));
  INV_X1    g704(.A(G127gat), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n906), .B1(new_n897), .B2(new_n742), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n905), .A2(new_n907), .ZN(G1342gat));
  INV_X1    g707(.A(G134gat), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n909), .B1(new_n897), .B2(new_n345), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT56), .ZN(new_n911));
  AND4_X1   g710(.A1(new_n909), .A2(new_n891), .A3(new_n345), .A4(new_n892), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n912), .A2(new_n911), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT115), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n914), .A2(new_n915), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n913), .B1(new_n917), .B2(new_n918), .ZN(G1343gat));
  NOR2_X1   g718(.A1(new_n803), .A2(new_n444), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n891), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n584), .B1(new_n921), .B2(KEYINPUT118), .ZN(new_n922));
  INV_X1    g721(.A(G141gat), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT118), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n891), .A2(new_n924), .A3(new_n920), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n922), .A2(new_n923), .A3(new_n684), .A4(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT58), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT57), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n868), .A2(KEYINPUT116), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT116), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n882), .A2(new_n930), .A3(new_n866), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n684), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n345), .B1(new_n932), .B2(new_n885), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n745), .A2(new_n875), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n261), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT117), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n859), .ZN(new_n938));
  OAI211_X1 g737(.A(KEYINPUT117), .B(new_n261), .C1(new_n933), .C2(new_n934), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n928), .B1(new_n940), .B2(new_n729), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n883), .A2(new_n885), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(KEYINPUT114), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n943), .A2(new_n745), .A3(new_n886), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n742), .B1(new_n944), .B2(new_n878), .ZN(new_n945));
  OAI211_X1 g744(.A(new_n928), .B(new_n729), .C1(new_n945), .C2(new_n859), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n803), .A2(new_n896), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n941), .A2(new_n948), .A3(new_n685), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n926), .B(new_n927), .C1(new_n949), .C2(new_n923), .ZN(new_n950));
  NOR4_X1   g749(.A1(new_n921), .A2(G141gat), .A3(new_n584), .A4(new_n685), .ZN(new_n951));
  INV_X1    g750(.A(new_n949), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n951), .B1(new_n952), .B2(G141gat), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n950), .B1(new_n953), .B2(new_n927), .ZN(G1344gat));
  INV_X1    g753(.A(G148gat), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n922), .A2(new_n955), .A3(new_n735), .A4(new_n925), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT59), .ZN(new_n957));
  INV_X1    g756(.A(new_n890), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(new_n729), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n933), .B1(new_n345), .B2(new_n876), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n938), .B1(new_n960), .B2(new_n348), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n444), .A2(KEYINPUT57), .ZN(new_n962));
  AOI22_X1  g761(.A1(new_n959), .A2(KEYINPUT57), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n963), .A2(new_n735), .A3(new_n947), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n957), .B1(new_n964), .B2(G148gat), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n941), .A2(new_n948), .ZN(new_n966));
  AOI211_X1 g765(.A(KEYINPUT59), .B(new_n955), .C1(new_n966), .C2(new_n735), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n956), .B1(new_n965), .B2(new_n967), .ZN(G1345gat));
  INV_X1    g767(.A(KEYINPUT119), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n941), .A2(new_n948), .A3(new_n741), .ZN(new_n970));
  INV_X1    g769(.A(G155gat), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n921), .A2(KEYINPUT118), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n261), .A2(G155gat), .ZN(new_n974));
  AND4_X1   g773(.A1(new_n567), .A2(new_n973), .A3(new_n925), .A4(new_n974), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n969), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n922), .A2(new_n925), .A3(new_n974), .ZN(new_n977));
  OAI211_X1 g776(.A(new_n977), .B(KEYINPUT119), .C1(new_n971), .C2(new_n970), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n976), .A2(new_n978), .ZN(G1346gat));
  NAND2_X1  g778(.A1(new_n966), .A2(new_n877), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(G162gat), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n347), .A2(G162gat), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n922), .A2(new_n925), .A3(new_n982), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT120), .ZN(new_n984));
  AND2_X1   g783(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n983), .A2(new_n984), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n981), .B1(new_n985), .B2(new_n986), .ZN(G1347gat));
  NOR2_X1   g786(.A1(new_n698), .A2(new_n567), .ZN(new_n988));
  NAND4_X1  g787(.A1(new_n958), .A2(new_n660), .A3(new_n444), .A4(new_n988), .ZN(new_n989));
  OAI21_X1  g788(.A(G169gat), .B1(new_n989), .B2(new_n685), .ZN(new_n990));
  XNOR2_X1  g789(.A(new_n990), .B(KEYINPUT123), .ZN(new_n991));
  OR2_X1    g790(.A1(new_n656), .A2(new_n567), .ZN(new_n992));
  XNOR2_X1  g791(.A(new_n992), .B(KEYINPUT122), .ZN(new_n993));
  OAI21_X1  g792(.A(KEYINPUT121), .B1(new_n890), .B2(new_n698), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT121), .ZN(new_n995));
  OAI211_X1 g794(.A(new_n995), .B(new_n494), .C1(new_n945), .C2(new_n859), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n993), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  INV_X1    g796(.A(G169gat), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n997), .A2(new_n998), .A3(new_n684), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n991), .A2(new_n999), .ZN(G1348gat));
  INV_X1    g799(.A(G176gat), .ZN(new_n1001));
  NOR3_X1   g800(.A1(new_n989), .A2(new_n1001), .A3(new_n830), .ZN(new_n1002));
  AOI21_X1  g801(.A(G176gat), .B1(new_n997), .B2(new_n735), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT124), .ZN(new_n1004));
  OR2_X1    g803(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1006));
  AOI21_X1  g805(.A(new_n1002), .B1(new_n1005), .B2(new_n1006), .ZN(G1349gat));
  OAI21_X1  g806(.A(G183gat), .B1(new_n989), .B2(new_n741), .ZN(new_n1008));
  INV_X1    g807(.A(KEYINPUT125), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n996), .ZN(new_n1010));
  INV_X1    g809(.A(new_n993), .ZN(new_n1011));
  AND2_X1   g810(.A1(new_n348), .A2(new_n504), .ZN(new_n1012));
  AND4_X1   g811(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AOI21_X1  g812(.A(new_n1009), .B1(new_n997), .B2(new_n1012), .ZN(new_n1014));
  OAI21_X1  g813(.A(new_n1008), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1015), .A2(KEYINPUT60), .ZN(new_n1016));
  INV_X1    g815(.A(KEYINPUT60), .ZN(new_n1017));
  OAI211_X1 g816(.A(new_n1017), .B(new_n1008), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n1016), .A2(new_n1018), .ZN(G1350gat));
  OAI21_X1  g818(.A(G190gat), .B1(new_n989), .B2(new_n347), .ZN(new_n1020));
  INV_X1    g819(.A(KEYINPUT126), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g821(.A(KEYINPUT126), .B(G190gat), .C1(new_n989), .C2(new_n347), .ZN(new_n1023));
  NAND3_X1  g822(.A1(new_n1022), .A2(KEYINPUT61), .A3(new_n1023), .ZN(new_n1024));
  NAND3_X1  g823(.A1(new_n997), .A2(new_n501), .A3(new_n877), .ZN(new_n1025));
  OAI211_X1 g824(.A(new_n1024), .B(new_n1025), .C1(KEYINPUT61), .C2(new_n1022), .ZN(G1351gat));
  NAND2_X1  g825(.A1(new_n920), .A2(new_n584), .ZN(new_n1027));
  AOI21_X1  g826(.A(new_n1027), .B1(new_n994), .B2(new_n996), .ZN(new_n1028));
  AOI21_X1  g827(.A(G197gat), .B1(new_n1028), .B2(new_n684), .ZN(new_n1029));
  AND2_X1   g828(.A1(new_n655), .A2(new_n988), .ZN(new_n1030));
  AND2_X1   g829(.A1(new_n963), .A2(new_n1030), .ZN(new_n1031));
  AND2_X1   g830(.A1(new_n684), .A2(G197gat), .ZN(new_n1032));
  AOI21_X1  g831(.A(new_n1029), .B1(new_n1031), .B2(new_n1032), .ZN(G1352gat));
  INV_X1    g832(.A(KEYINPUT62), .ZN(new_n1034));
  INV_X1    g833(.A(KEYINPUT127), .ZN(new_n1035));
  NOR2_X1   g834(.A1(new_n374), .A2(G204gat), .ZN(new_n1036));
  NAND3_X1  g835(.A1(new_n1028), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g836(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g837(.A(new_n1035), .B1(new_n1028), .B2(new_n1036), .ZN(new_n1039));
  OAI21_X1  g838(.A(new_n1034), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g839(.A(new_n1039), .ZN(new_n1041));
  NAND3_X1  g840(.A1(new_n1041), .A2(KEYINPUT62), .A3(new_n1037), .ZN(new_n1042));
  NAND3_X1  g841(.A1(new_n963), .A2(new_n740), .A3(new_n1030), .ZN(new_n1043));
  NAND2_X1  g842(.A1(new_n1043), .A2(G204gat), .ZN(new_n1044));
  NAND3_X1  g843(.A1(new_n1040), .A2(new_n1042), .A3(new_n1044), .ZN(G1353gat));
  NAND3_X1  g844(.A1(new_n1028), .A2(new_n397), .A3(new_n348), .ZN(new_n1046));
  NAND3_X1  g845(.A1(new_n963), .A2(new_n348), .A3(new_n1030), .ZN(new_n1047));
  AND3_X1   g846(.A1(new_n1047), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1048));
  AOI21_X1  g847(.A(KEYINPUT63), .B1(new_n1047), .B2(G211gat), .ZN(new_n1049));
  OAI21_X1  g848(.A(new_n1046), .B1(new_n1048), .B2(new_n1049), .ZN(G1354gat));
  NAND3_X1  g849(.A1(new_n1028), .A2(new_n398), .A3(new_n877), .ZN(new_n1051));
  AND2_X1   g850(.A1(new_n1031), .A2(new_n345), .ZN(new_n1052));
  OAI21_X1  g851(.A(new_n1051), .B1(new_n1052), .B2(new_n398), .ZN(G1355gat));
endmodule


