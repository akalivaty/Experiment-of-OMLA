//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 0 1 0 0 0 0 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n986, new_n987, new_n988;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT15), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT14), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n206), .B(KEYINPUT92), .C1(G29gat), .C2(G36gat), .ZN(new_n207));
  INV_X1    g006(.A(G29gat), .ZN(new_n208));
  INV_X1    g007(.A(G36gat), .ZN(new_n209));
  OAI221_X1 g008(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n203), .C2(KEYINPUT15), .ZN(new_n210));
  OR3_X1    g009(.A1(KEYINPUT92), .A2(G29gat), .A3(G36gat), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT92), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(KEYINPUT14), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n205), .B1(new_n210), .B2(new_n214), .ZN(new_n215));
  XOR2_X1   g014(.A(G43gat), .B(G50gat), .Z(new_n216));
  INV_X1    g015(.A(KEYINPUT15), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n216), .A2(new_n217), .B1(G29gat), .B2(G36gat), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n218), .A2(new_n204), .A3(new_n213), .A4(new_n207), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT93), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G15gat), .B(G22gat), .ZN(new_n223));
  OR2_X1    g022(.A1(new_n223), .A2(G1gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT16), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n223), .B1(new_n225), .B2(G1gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G8gat), .ZN(new_n228));
  INV_X1    g027(.A(G8gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n224), .A2(new_n229), .A3(new_n226), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n219), .A3(KEYINPUT93), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n222), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  XOR2_X1   g032(.A(KEYINPUT94), .B(KEYINPUT17), .Z(new_n234));
  AND3_X1   g033(.A1(new_n222), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n231), .A2(KEYINPUT95), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n215), .A2(new_n219), .A3(KEYINPUT17), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT95), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n228), .A2(new_n238), .A3(new_n230), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n236), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n202), .B(new_n233), .C1(new_n235), .C2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT18), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n222), .A2(new_n232), .ZN(new_n244));
  INV_X1    g043(.A(new_n231), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(new_n233), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n202), .B(KEYINPUT13), .Z(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n222), .A2(new_n232), .A3(new_n234), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n250), .A2(new_n237), .A3(new_n239), .A4(new_n236), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n251), .A2(KEYINPUT18), .A3(new_n202), .A4(new_n233), .ZN(new_n252));
  XNOR2_X1  g051(.A(G113gat), .B(G141gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G169gat), .B(G197gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(KEYINPUT12), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n243), .A2(new_n249), .A3(new_n252), .A4(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n241), .A2(new_n242), .B1(new_n247), .B2(new_n248), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n258), .B1(new_n261), .B2(new_n252), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT64), .ZN(new_n264));
  NOR2_X1   g063(.A1(G169gat), .A2(G176gat), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n264), .B1(new_n265), .B2(KEYINPUT23), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT23), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n267), .B(KEYINPUT64), .C1(G169gat), .C2(G176gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G183gat), .A2(G190gat), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT24), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(G183gat), .ZN(new_n273));
  INV_X1    g072(.A(G190gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n272), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  AND2_X1   g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n278), .B1(KEYINPUT23), .B2(new_n265), .ZN(new_n279));
  AND3_X1   g078(.A1(new_n269), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT65), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n270), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(new_n271), .A3(new_n283), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n284), .A2(new_n275), .A3(new_n276), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n269), .A2(KEYINPUT25), .A3(new_n279), .ZN(new_n286));
  OAI22_X1  g085(.A1(new_n280), .A2(KEYINPUT25), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT67), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI211_X1 g089(.A(KEYINPUT67), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT26), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n278), .B1(new_n293), .B2(new_n265), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT68), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(new_n296), .A3(new_n270), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT28), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT66), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT27), .B(G183gat), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n299), .B1(new_n300), .B2(new_n274), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n273), .A2(KEYINPUT27), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT27), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G183gat), .ZN(new_n304));
  AND4_X1   g103(.A1(new_n299), .A2(new_n302), .A3(new_n304), .A4(new_n274), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n298), .B1(new_n301), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n302), .A2(new_n304), .A3(new_n274), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT66), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n300), .A2(new_n299), .A3(new_n274), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n308), .A2(new_n309), .A3(KEYINPUT28), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n297), .A2(new_n306), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n296), .B1(new_n295), .B2(new_n270), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n287), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(KEYINPUT71), .B(G120gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G113gat), .ZN(new_n315));
  INV_X1    g114(.A(G113gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(G120gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n315), .A2(KEYINPUT72), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT72), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n314), .A2(new_n319), .A3(G113gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT73), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT1), .ZN(new_n322));
  INV_X1    g121(.A(G134gat), .ZN(new_n323));
  OAI22_X1  g122(.A1(new_n321), .A2(new_n322), .B1(new_n323), .B2(G127gat), .ZN(new_n324));
  INV_X1    g123(.A(G127gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n325), .A2(G134gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(KEYINPUT73), .A2(KEYINPUT1), .ZN(new_n327));
  NOR3_X1   g126(.A1(new_n324), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n318), .A2(new_n320), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT69), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n330), .A2(new_n325), .A3(G134gat), .ZN(new_n331));
  OAI21_X1  g130(.A(KEYINPUT69), .B1(new_n323), .B2(G127gat), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n331), .B1(new_n332), .B2(new_n326), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT70), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT70), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n335), .B(new_n331), .C1(new_n332), .C2(new_n326), .ZN(new_n336));
  XOR2_X1   g135(.A(G113gat), .B(G120gat), .Z(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(new_n322), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n334), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n329), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n313), .A2(new_n341), .ZN(new_n342));
  AND2_X1   g141(.A1(G227gat), .A2(G233gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n295), .A2(new_n270), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT68), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n345), .A2(new_n297), .A3(new_n306), .A4(new_n310), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n346), .A2(new_n340), .A3(new_n287), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n342), .A2(new_n343), .A3(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G15gat), .B(G43gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(G71gat), .B(G99gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  XOR2_X1   g150(.A(KEYINPUT74), .B(KEYINPUT33), .Z(new_n352));
  OR2_X1    g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n348), .A2(KEYINPUT32), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT75), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT75), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n348), .A2(new_n356), .A3(KEYINPUT32), .A4(new_n353), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n351), .B1(new_n348), .B2(KEYINPUT32), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n348), .A2(new_n352), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  AND2_X1   g161(.A1(new_n342), .A2(new_n347), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n363), .A2(new_n343), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  XOR2_X1   g164(.A(KEYINPUT76), .B(KEYINPUT34), .Z(new_n366));
  INV_X1    g165(.A(new_n364), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n358), .A2(new_n367), .A3(new_n361), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n365), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n366), .ZN(new_n370));
  AOI221_X4 g169(.A(new_n364), .B1(new_n359), .B2(new_n360), .C1(new_n355), .C2(new_n357), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n367), .B1(new_n358), .B2(new_n361), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT77), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n369), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT36), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G78gat), .B(G106gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(KEYINPUT31), .B(G50gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(G211gat), .B(G218gat), .Z(new_n381));
  INV_X1    g180(.A(KEYINPUT79), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT22), .ZN(new_n383));
  INV_X1    g182(.A(G211gat), .ZN(new_n384));
  INV_X1    g183(.A(G218gat), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AOI22_X1  g185(.A1(new_n381), .A2(new_n382), .B1(KEYINPUT78), .B2(new_n386), .ZN(new_n387));
  OR2_X1    g186(.A1(new_n386), .A2(KEYINPUT78), .ZN(new_n388));
  INV_X1    g187(.A(G204gat), .ZN(new_n389));
  OR2_X1    g188(.A1(new_n389), .A2(G197gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(G197gat), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n387), .A2(new_n388), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n381), .A2(new_n382), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT84), .ZN(new_n395));
  AND2_X1   g194(.A1(KEYINPUT83), .A2(G141gat), .ZN(new_n396));
  NOR2_X1   g195(.A1(KEYINPUT83), .A2(G141gat), .ZN(new_n397));
  INV_X1    g196(.A(G148gat), .ZN(new_n398));
  NOR3_X1   g197(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(G141gat), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n400), .A2(G148gat), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n395), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n401), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT83), .B(G141gat), .ZN(new_n404));
  OAI211_X1 g203(.A(KEYINPUT84), .B(new_n403), .C1(new_n404), .C2(new_n398), .ZN(new_n405));
  NAND2_X1  g204(.A1(G155gat), .A2(G162gat), .ZN(new_n406));
  INV_X1    g205(.A(G155gat), .ZN(new_n407));
  INV_X1    g206(.A(G162gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n406), .B1(new_n409), .B2(KEYINPUT2), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n402), .A2(new_n405), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT3), .ZN(new_n412));
  XNOR2_X1  g211(.A(G141gat), .B(G148gat), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n406), .B(new_n409), .C1(new_n413), .C2(KEYINPUT2), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n411), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n394), .B1(KEYINPUT29), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT86), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n419), .A2(G228gat), .A3(G233gat), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n412), .B1(new_n394), .B2(KEYINPUT29), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n411), .A2(new_n414), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(G22gat), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(new_n425), .A3(new_n417), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n425), .B1(new_n424), .B2(new_n417), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n421), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n424), .A2(new_n417), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(G22gat), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n431), .A2(new_n426), .A3(new_n420), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n380), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n429), .A2(new_n380), .A3(new_n432), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G1gat), .B(G29gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n437), .B(KEYINPUT0), .ZN(new_n438));
  XNOR2_X1  g237(.A(G57gat), .B(G85gat), .ZN(new_n439));
  XOR2_X1   g238(.A(new_n438), .B(new_n439), .Z(new_n440));
  NAND2_X1  g239(.A1(new_n423), .A2(KEYINPUT3), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n441), .A2(new_n415), .A3(new_n340), .ZN(new_n442));
  INV_X1    g241(.A(new_n423), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n341), .A2(new_n443), .A3(KEYINPUT4), .ZN(new_n444));
  NAND2_X1  g243(.A1(G225gat), .A2(G233gat), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n329), .A2(new_n411), .A3(new_n414), .A4(new_n339), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT4), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n442), .A2(new_n444), .A3(new_n445), .A4(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT5), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n340), .A2(new_n423), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n446), .ZN(new_n452));
  INV_X1    g251(.A(new_n445), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n450), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT85), .B1(new_n449), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n449), .A2(new_n454), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n446), .B(KEYINPUT4), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n458), .A2(new_n450), .A3(new_n445), .A4(new_n442), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT85), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n440), .B(new_n456), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT6), .ZN(new_n463));
  INV_X1    g262(.A(new_n440), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n461), .B1(new_n457), .B2(new_n459), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n464), .B1(new_n465), .B2(new_n455), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n462), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  OAI211_X1 g266(.A(KEYINPUT6), .B(new_n464), .C1(new_n465), .C2(new_n455), .ZN(new_n468));
  AND2_X1   g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  XOR2_X1   g268(.A(G8gat), .B(G36gat), .Z(new_n470));
  XNOR2_X1  g269(.A(new_n470), .B(KEYINPUT80), .ZN(new_n471));
  XNOR2_X1  g270(.A(G64gat), .B(G92gat), .ZN(new_n472));
  XOR2_X1   g271(.A(new_n471), .B(new_n472), .Z(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  AND2_X1   g273(.A1(G226gat), .A2(G233gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n313), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT29), .B1(new_n346), .B2(new_n287), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n476), .B1(new_n477), .B2(new_n475), .ZN(new_n478));
  INV_X1    g277(.A(new_n394), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n476), .B(new_n394), .C1(new_n477), .C2(new_n475), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n474), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT30), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT82), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n482), .A2(KEYINPUT82), .A3(KEYINPUT30), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n480), .A2(new_n481), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT81), .B1(new_n488), .B2(new_n473), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT81), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n480), .A2(new_n490), .A3(new_n474), .A4(new_n481), .ZN(new_n491));
  INV_X1    g290(.A(new_n482), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT30), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n489), .A2(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n487), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n436), .B1(new_n469), .B2(new_n495), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n369), .A2(new_n373), .A3(new_n374), .A4(KEYINPUT36), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n377), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT87), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n377), .A2(new_n496), .A3(KEYINPUT87), .A4(new_n497), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT37), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n488), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT38), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n474), .B1(new_n488), .B2(new_n502), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n492), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT90), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g308(.A(KEYINPUT90), .B(new_n474), .C1(new_n488), .C2(new_n502), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(new_n510), .A3(new_n503), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n507), .B1(new_n511), .B2(KEYINPUT38), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n468), .A2(KEYINPUT89), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n512), .B(new_n513), .C1(new_n469), .C2(KEYINPUT89), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n458), .A2(new_n442), .ZN(new_n515));
  XOR2_X1   g314(.A(KEYINPUT88), .B(KEYINPUT39), .Z(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n453), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n440), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT39), .B1(new_n452), .B2(new_n453), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n519), .B1(new_n515), .B2(new_n453), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT40), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT40), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n523), .B1(new_n518), .B2(new_n520), .ZN(new_n524));
  AND3_X1   g323(.A1(new_n522), .A2(new_n466), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n436), .B1(new_n495), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n514), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n500), .A2(new_n501), .A3(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n495), .A2(KEYINPUT35), .ZN(new_n529));
  INV_X1    g328(.A(new_n435), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n530), .A2(new_n433), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n369), .A2(new_n373), .ZN(new_n532));
  AND3_X1   g331(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n513), .B1(new_n469), .B2(KEYINPUT89), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n467), .A2(new_n468), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n487), .A2(new_n494), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n532), .A2(new_n536), .A3(new_n537), .A4(new_n531), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT35), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n263), .B1(new_n528), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT21), .ZN(new_n542));
  INV_X1    g341(.A(G57gat), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n543), .A2(G64gat), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n543), .A2(G64gat), .ZN(new_n545));
  AND2_X1   g344(.A1(G71gat), .A2(G78gat), .ZN(new_n546));
  OAI22_X1  g345(.A1(new_n544), .A2(new_n545), .B1(new_n546), .B2(KEYINPUT9), .ZN(new_n547));
  XNOR2_X1  g346(.A(G71gat), .B(G78gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n245), .B1(new_n542), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n542), .ZN(new_n552));
  NAND2_X1  g351(.A1(G231gat), .A2(G233gat), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n552), .B(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(G127gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n552), .B(new_n553), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n325), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n551), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n556), .A2(new_n558), .A3(new_n551), .ZN(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(new_n407), .ZN(new_n563));
  XNOR2_X1  g362(.A(G183gat), .B(G211gat), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n563), .B(new_n564), .Z(new_n565));
  NAND3_X1  g364(.A1(new_n560), .A2(new_n561), .A3(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n565), .ZN(new_n567));
  INV_X1    g366(.A(new_n561), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n567), .B1(new_n568), .B2(new_n559), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(G134gat), .B(G162gat), .Z(new_n572));
  AND2_X1   g371(.A1(G232gat), .A2(G233gat), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n573), .A2(KEYINPUT41), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n572), .B(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(KEYINPUT96), .B(KEYINPUT97), .Z(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G99gat), .B(G106gat), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(G85gat), .ZN(new_n581));
  INV_X1    g380(.A(G92gat), .ZN(new_n582));
  OAI21_X1  g381(.A(KEYINPUT98), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT98), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n584), .A2(G85gat), .A3(G92gat), .ZN(new_n585));
  AND3_X1   g384(.A1(new_n583), .A2(KEYINPUT7), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G99gat), .A2(G106gat), .ZN(new_n587));
  AOI22_X1  g386(.A1(KEYINPUT8), .A2(new_n587), .B1(new_n581), .B2(new_n582), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT7), .ZN(new_n589));
  OAI211_X1 g388(.A(KEYINPUT98), .B(new_n589), .C1(new_n581), .C2(new_n582), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n580), .B1(new_n586), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n583), .A2(KEYINPUT7), .A3(new_n585), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n593), .A2(new_n579), .A3(new_n590), .A4(new_n588), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n592), .A2(KEYINPUT99), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT99), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n596), .B(new_n580), .C1(new_n586), .C2(new_n591), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n250), .A2(new_n237), .A3(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G190gat), .B(G218gat), .Z(new_n601));
  NAND3_X1  g400(.A1(new_n222), .A2(new_n232), .A3(new_n598), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n573), .A2(KEYINPUT41), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR3_X1   g403(.A1(new_n600), .A2(new_n601), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n601), .ZN(new_n606));
  INV_X1    g405(.A(new_n604), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n250), .A2(new_n237), .A3(new_n599), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n578), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n601), .B1(new_n600), .B2(new_n604), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n607), .A2(new_n606), .A3(new_n608), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(new_n577), .A3(new_n612), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(KEYINPUT100), .B1(new_n571), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT100), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n610), .A2(new_n613), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n570), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G230gat), .A2(G233gat), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n550), .A2(new_n595), .A3(new_n597), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT10), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n549), .A2(new_n592), .A3(new_n594), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n598), .A2(KEYINPUT10), .A3(new_n549), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n621), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n620), .B1(new_n622), .B2(new_n624), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G120gat), .B(G148gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(G176gat), .B(G204gat), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n630), .B(new_n631), .Z(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT101), .ZN(new_n635));
  OR3_X1    g434(.A1(new_n627), .A2(new_n628), .A3(new_n633), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n629), .A2(KEYINPUT101), .A3(new_n633), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n619), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n541), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n469), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g444(.A(KEYINPUT16), .B(G8gat), .Z(new_n646));
  NAND3_X1  g445(.A1(new_n643), .A2(new_n495), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(G8gat), .B1(new_n642), .B2(new_n537), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  MUX2_X1   g448(.A(new_n647), .B(new_n649), .S(KEYINPUT42), .Z(G1325gat));
  AOI21_X1  g449(.A(G15gat), .B1(new_n643), .B2(new_n532), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n377), .A2(new_n497), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(KEYINPUT102), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n377), .A2(new_n654), .A3(new_n497), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(G15gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT103), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n651), .B1(new_n643), .B2(new_n658), .ZN(G1326gat));
  NAND3_X1  g458(.A1(new_n541), .A2(new_n436), .A3(new_n641), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT104), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT43), .B(G22gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(G1327gat));
  NOR2_X1   g462(.A1(new_n640), .A2(new_n570), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n614), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n541), .A2(new_n208), .A3(new_n469), .A4(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT45), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OR2_X1    g468(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n617), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n673), .B1(new_n528), .B2(new_n540), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n531), .B1(new_n536), .B2(new_n537), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n675), .B1(new_n514), .B2(new_n526), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n653), .A2(new_n676), .A3(new_n655), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n540), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n614), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n674), .B1(new_n679), .B2(new_n671), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n263), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n664), .A2(new_n682), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n681), .A2(new_n536), .A3(new_n683), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n669), .B(new_n670), .C1(new_n684), .C2(new_n208), .ZN(G1328gat));
  NAND4_X1  g484(.A1(new_n541), .A2(new_n209), .A3(new_n495), .A4(new_n666), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(KEYINPUT46), .Z(new_n687));
  NOR3_X1   g486(.A1(new_n681), .A2(new_n537), .A3(new_n683), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n687), .B1(new_n209), .B2(new_n688), .ZN(G1329gat));
  INV_X1    g488(.A(new_n532), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n690), .A2(G43gat), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n541), .A2(new_n666), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(KEYINPUT106), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n541), .A2(new_n694), .A3(new_n666), .A4(new_n691), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n697));
  AOI21_X1  g496(.A(KEYINPUT47), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(KEYINPUT44), .B1(new_n678), .B2(new_n614), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n377), .A2(new_n654), .A3(new_n497), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n654), .B1(new_n377), .B2(new_n497), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR4_X1   g501(.A1(new_n699), .A2(new_n674), .A3(new_n702), .A4(new_n683), .ZN(new_n703));
  INV_X1    g502(.A(G43gat), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n696), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n698), .A2(new_n705), .ZN(new_n706));
  OAI221_X1 g505(.A(new_n696), .B1(new_n697), .B2(KEYINPUT47), .C1(new_n703), .C2(new_n704), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(G1330gat));
  INV_X1    g507(.A(G50gat), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n541), .A2(new_n709), .A3(new_n436), .A4(new_n666), .ZN(new_n710));
  NOR4_X1   g509(.A1(new_n699), .A2(new_n674), .A3(new_n531), .A4(new_n683), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n710), .B1(new_n711), .B2(new_n709), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT48), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OAI211_X1 g513(.A(KEYINPUT48), .B(new_n710), .C1(new_n711), .C2(new_n709), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(G1331gat));
  AOI22_X1  g515(.A1(new_n533), .A2(new_n534), .B1(KEYINPUT35), .B2(new_n538), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n717), .B1(new_n702), .B2(new_n676), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n615), .A2(new_n263), .A3(new_n618), .A4(new_n640), .ZN(new_n719));
  XOR2_X1   g518(.A(new_n719), .B(KEYINPUT107), .Z(new_n720));
  NOR2_X1   g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n469), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g522(.A(new_n537), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n725), .B(new_n726), .Z(G1333gat));
  NAND2_X1  g526(.A1(new_n721), .A2(new_n656), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n690), .A2(G71gat), .ZN(new_n729));
  AOI22_X1  g528(.A1(new_n728), .A2(G71gat), .B1(new_n721), .B2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g530(.A1(new_n721), .A2(new_n436), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g532(.A1(new_n536), .A2(G85gat), .A3(new_n639), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT108), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n617), .B1(new_n677), .B2(new_n540), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n682), .A2(new_n570), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n736), .A2(KEYINPUT51), .A3(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(KEYINPUT51), .B1(new_n736), .B2(new_n737), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n735), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n737), .A2(new_n640), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n699), .A2(new_n674), .A3(new_n742), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n743), .A2(new_n469), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n741), .B1(new_n744), .B2(new_n581), .ZN(G1336gat));
  NOR3_X1   g544(.A1(new_n537), .A2(G92gat), .A3(new_n639), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n746), .B1(new_n739), .B2(new_n740), .ZN(new_n747));
  NOR4_X1   g546(.A1(new_n699), .A2(new_n674), .A3(new_n537), .A4(new_n742), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n748), .B2(new_n582), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT52), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n747), .B(new_n751), .C1(new_n748), .C2(new_n582), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(G1337gat));
  INV_X1    g552(.A(G99gat), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n754), .B1(new_n743), .B2(new_n656), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n690), .A2(G99gat), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n678), .A2(new_n614), .A3(new_n737), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI211_X1 g559(.A(new_n639), .B(new_n757), .C1(new_n760), .C2(new_n738), .ZN(new_n761));
  OAI21_X1  g560(.A(KEYINPUT109), .B1(new_n755), .B2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n742), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n680), .A2(new_n656), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(G99gat), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n639), .B1(new_n760), .B2(new_n738), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n756), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n765), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n762), .A2(new_n769), .ZN(G1338gat));
  OAI21_X1  g569(.A(new_n671), .B1(new_n718), .B2(new_n617), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n528), .A2(new_n540), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n672), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n771), .A2(new_n436), .A3(new_n773), .A4(new_n763), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n680), .A2(KEYINPUT110), .A3(new_n436), .A4(new_n763), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n776), .A2(G106gat), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n531), .A2(G106gat), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT53), .B1(new_n766), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n774), .A2(G106gat), .ZN(new_n782));
  INV_X1    g581(.A(new_n779), .ZN(new_n783));
  AOI211_X1 g582(.A(new_n639), .B(new_n783), .C1(new_n760), .C2(new_n738), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT53), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n781), .A2(new_n785), .ZN(G1339gat));
  AND4_X1   g585(.A1(new_n263), .A2(new_n615), .A3(new_n618), .A4(new_n639), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n202), .B1(new_n251), .B2(new_n233), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n247), .A2(new_n248), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n257), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n259), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n627), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n625), .A2(new_n626), .A3(KEYINPUT111), .A4(new_n621), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n625), .A2(new_n626), .A3(new_n621), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n793), .A2(new_n794), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n632), .B1(new_n627), .B2(new_n792), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT55), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n614), .A2(new_n791), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n798), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n799), .A2(KEYINPUT55), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT112), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n798), .A2(new_n806), .A3(KEYINPUT55), .A4(new_n799), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n805), .A2(new_n636), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(KEYINPUT113), .B1(new_n802), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n259), .A2(new_n790), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n617), .A2(new_n810), .A3(new_n800), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n807), .A2(new_n636), .ZN(new_n812));
  INV_X1    g611(.A(new_n804), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n806), .B1(new_n813), .B2(new_n798), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT113), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n811), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n261), .A2(new_n252), .ZN(new_n818));
  INV_X1    g617(.A(new_n258), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n800), .B1(new_n820), .B2(new_n259), .ZN(new_n821));
  AOI22_X1  g620(.A1(new_n815), .A2(new_n821), .B1(new_n640), .B2(new_n791), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n809), .B(new_n817), .C1(new_n822), .C2(new_n614), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n570), .B1(new_n823), .B2(KEYINPUT114), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n801), .B1(new_n260), .B2(new_n262), .ZN(new_n825));
  OAI22_X1  g624(.A1(new_n825), .A2(new_n808), .B1(new_n639), .B2(new_n810), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n617), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n827), .A2(new_n828), .A3(new_n809), .A4(new_n817), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n787), .B1(new_n824), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(new_n536), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n690), .A2(new_n436), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(new_n495), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(G113gat), .B1(new_n835), .B2(new_n682), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n830), .A2(new_n436), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n537), .A2(new_n469), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n690), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n840), .A2(new_n316), .A3(new_n263), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n836), .A2(new_n841), .ZN(G1340gat));
  NAND3_X1  g641(.A1(new_n835), .A2(new_n314), .A3(new_n640), .ZN(new_n843));
  OAI21_X1  g642(.A(G120gat), .B1(new_n840), .B2(new_n639), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(G1341gat));
  INV_X1    g644(.A(new_n840), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(G127gat), .A3(new_n570), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n847), .A2(new_n848), .ZN(new_n850));
  AOI21_X1  g649(.A(G127gat), .B1(new_n835), .B2(new_n570), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(G1342gat));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n809), .A2(new_n817), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n815), .A2(new_n821), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n640), .A2(new_n791), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n614), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT114), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n829), .A3(new_n571), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n615), .A2(new_n263), .A3(new_n618), .A4(new_n639), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n617), .A2(G134gat), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n861), .A2(new_n469), .A3(new_n834), .A4(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT116), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n863), .B(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n853), .B1(new_n865), .B2(KEYINPUT56), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n863), .A2(new_n864), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT56), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n863), .A2(new_n864), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n867), .A2(KEYINPUT117), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n323), .B1(new_n846), .B2(new_n614), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n872), .B1(KEYINPUT56), .B2(new_n865), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(G1343gat));
  NOR2_X1   g673(.A1(new_n656), .A2(new_n838), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT57), .B1(new_n861), .B2(new_n436), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n531), .A2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n823), .A2(new_n571), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n879), .B1(new_n880), .B2(new_n860), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n682), .B(new_n875), .C1(new_n876), .C2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n404), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT118), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n656), .A2(new_n531), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n831), .A2(new_n537), .A3(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n263), .A2(G141gat), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n883), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n884), .A2(new_n890), .A3(KEYINPUT58), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT58), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n883), .B(new_n889), .C1(KEYINPUT118), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n893), .ZN(G1344gat));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895));
  AOI211_X1 g694(.A(new_n895), .B(G148gat), .C1(new_n887), .C2(new_n640), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n875), .B1(new_n876), .B2(new_n881), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n895), .B1(new_n897), .B2(new_n639), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n879), .B1(new_n859), .B2(new_n860), .ZN(new_n899));
  OAI22_X1  g698(.A1(new_n822), .A2(new_n614), .B1(new_n808), .B2(new_n802), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n571), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n860), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT57), .B1(new_n902), .B2(new_n436), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n875), .A2(KEYINPUT119), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n875), .A2(KEYINPUT119), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n905), .A2(KEYINPUT59), .A3(new_n640), .A4(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n898), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n896), .B1(new_n908), .B2(G148gat), .ZN(G1345gat));
  OAI21_X1  g708(.A(new_n407), .B1(new_n886), .B2(new_n571), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n570), .A2(G155gat), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT120), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n875), .B(new_n912), .C1(new_n876), .C2(new_n881), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT121), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n914), .B(new_n915), .ZN(G1346gat));
  OAI21_X1  g715(.A(G162gat), .B1(new_n897), .B2(new_n617), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n887), .A2(new_n408), .A3(new_n614), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT122), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n917), .A2(new_n918), .A3(KEYINPUT122), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1347gat));
  NAND2_X1  g722(.A1(new_n861), .A2(new_n536), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n924), .A2(new_n537), .A3(new_n833), .ZN(new_n925));
  AOI21_X1  g724(.A(G169gat), .B1(new_n925), .B2(new_n682), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n495), .A2(new_n536), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n690), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n837), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(G169gat), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n929), .A2(new_n930), .A3(new_n263), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n926), .A2(new_n931), .ZN(G1348gat));
  NOR2_X1   g731(.A1(new_n537), .A2(new_n639), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  OR4_X1    g733(.A1(G176gat), .A2(new_n924), .A3(new_n833), .A4(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(G176gat), .B1(new_n929), .B2(new_n639), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1349gat));
  NAND4_X1  g736(.A1(new_n861), .A2(new_n531), .A3(new_n570), .A4(new_n928), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n273), .B1(new_n938), .B2(KEYINPUT123), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n939), .B1(KEYINPUT123), .B2(new_n938), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n570), .A2(new_n300), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT124), .B1(new_n925), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(KEYINPUT60), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT60), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n940), .A2(new_n942), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n944), .A2(new_n946), .ZN(G1350gat));
  NAND3_X1  g746(.A1(new_n837), .A2(new_n614), .A3(new_n928), .ZN(new_n948));
  AOI21_X1  g747(.A(KEYINPUT125), .B1(new_n948), .B2(G190gat), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT61), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n617), .A2(G190gat), .ZN(new_n951));
  AOI22_X1  g750(.A1(new_n949), .A2(new_n950), .B1(new_n925), .B2(new_n951), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n949), .A2(new_n950), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n948), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(G1351gat));
  NOR2_X1   g754(.A1(new_n656), .A2(new_n927), .ZN(new_n956));
  OAI211_X1 g755(.A(new_n956), .B(new_n682), .C1(new_n899), .C2(new_n903), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT126), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n787), .B1(new_n571), .B2(new_n900), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n877), .B1(new_n960), .B2(new_n531), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n961), .B1(new_n830), .B2(new_n879), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n962), .A2(KEYINPUT126), .A3(new_n682), .A4(new_n956), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n959), .A2(new_n963), .A3(G197gat), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n924), .A2(new_n531), .A3(new_n656), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n263), .A2(G197gat), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n965), .A2(new_n495), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n964), .A2(KEYINPUT127), .A3(new_n967), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(G1352gat));
  NAND3_X1  g771(.A1(new_n965), .A2(new_n389), .A3(new_n933), .ZN(new_n973));
  OR2_X1    g772(.A1(new_n973), .A2(KEYINPUT62), .ZN(new_n974));
  AND2_X1   g773(.A1(new_n962), .A2(new_n956), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(new_n640), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(G204gat), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n973), .A2(KEYINPUT62), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n974), .A2(new_n977), .A3(new_n978), .ZN(G1353gat));
  AND2_X1   g778(.A1(new_n965), .A2(new_n495), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n980), .A2(new_n384), .A3(new_n570), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n975), .A2(new_n570), .ZN(new_n982));
  AND3_X1   g781(.A1(new_n982), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n983));
  AOI21_X1  g782(.A(KEYINPUT63), .B1(new_n982), .B2(G211gat), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n981), .B1(new_n983), .B2(new_n984), .ZN(G1354gat));
  NAND3_X1  g784(.A1(new_n980), .A2(new_n385), .A3(new_n614), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n975), .A2(new_n614), .ZN(new_n987));
  INV_X1    g786(.A(new_n987), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n986), .B1(new_n988), .B2(new_n385), .ZN(G1355gat));
endmodule


