//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0 1 1 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1017, new_n1018;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT34), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT72), .ZN(new_n204));
  INV_X1    g003(.A(G183gat), .ZN(new_n205));
  AOI21_X1  g004(.A(G190gat), .B1(new_n205), .B2(KEYINPUT27), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT27), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G183gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n206), .A2(KEYINPUT28), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT69), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(new_n205), .B2(KEYINPUT27), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n207), .A2(KEYINPUT69), .A3(G183gat), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n212), .A2(new_n206), .A3(KEYINPUT70), .A4(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT28), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n212), .A2(new_n206), .A3(new_n213), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT70), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n210), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  OR3_X1    g021(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT71), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT26), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT71), .B1(new_n221), .B2(new_n222), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n223), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n204), .B1(new_n220), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n219), .A2(new_n215), .A3(new_n214), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(new_n209), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n230), .A2(new_n231), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n235), .A2(new_n236), .A3(KEYINPUT72), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n233), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND4_X1  g040(.A1(KEYINPUT66), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT24), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n231), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G190gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n205), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n241), .A2(new_n242), .A3(new_n244), .A4(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n225), .A2(KEYINPUT23), .A3(new_n227), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT25), .ZN(new_n249));
  NAND2_X1  g048(.A1(G169gat), .A2(G176gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(KEYINPUT23), .ZN(new_n251));
  INV_X1    g050(.A(G169gat), .ZN(new_n252));
  INV_X1    g051(.A(G176gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n249), .B1(new_n251), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n247), .A2(new_n248), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n247), .A2(new_n248), .A3(new_n255), .A4(KEYINPUT67), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n222), .A2(KEYINPUT23), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n261), .B1(new_n254), .B2(new_n251), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n246), .A2(KEYINPUT64), .ZN(new_n263));
  OR3_X1    g062(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n263), .A2(new_n264), .A3(new_n239), .A4(new_n244), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(new_n249), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT68), .ZN(new_n269));
  AOI22_X1  g068(.A1(new_n258), .A2(new_n259), .B1(new_n266), .B2(new_n249), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT68), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n238), .A2(new_n269), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT73), .ZN(new_n274));
  XOR2_X1   g073(.A(G127gat), .B(G134gat), .Z(new_n275));
  XNOR2_X1  g074(.A(G113gat), .B(G120gat), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n275), .B1(KEYINPUT1), .B2(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(G113gat), .B(G120gat), .Z(new_n278));
  INV_X1    g077(.A(KEYINPUT1), .ZN(new_n279));
  XNOR2_X1  g078(.A(G127gat), .B(G134gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n238), .A2(new_n269), .A3(new_n283), .A4(new_n272), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n274), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  AND2_X1   g084(.A1(new_n277), .A2(new_n281), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n273), .A2(KEYINPUT73), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G227gat), .ZN(new_n289));
  INV_X1    g088(.A(G233gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n203), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  AOI211_X1 g092(.A(KEYINPUT34), .B(new_n291), .C1(new_n285), .C2(new_n287), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n285), .A2(new_n291), .A3(new_n287), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT32), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT33), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT74), .B(G71gat), .ZN(new_n300));
  INV_X1    g099(.A(G99gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  XOR2_X1   g101(.A(G15gat), .B(G43gat), .Z(new_n303));
  XOR2_X1   g102(.A(new_n302), .B(new_n303), .Z(new_n304));
  AND3_X1   g103(.A1(new_n297), .A2(new_n299), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n304), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n296), .B(KEYINPUT32), .C1(new_n298), .C2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n202), .B(new_n295), .C1(new_n305), .C2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n288), .A2(new_n292), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT34), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n288), .A2(new_n203), .A3(new_n292), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n311), .A2(new_n202), .A3(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT75), .B1(new_n293), .B2(new_n294), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n297), .A2(new_n299), .A3(new_n304), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n313), .A2(new_n314), .A3(new_n307), .A4(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n309), .A2(new_n316), .A3(KEYINPUT88), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT88), .B1(new_n309), .B2(new_n316), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT87), .ZN(new_n320));
  NAND2_X1  g119(.A1(G226gat), .A2(G233gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n322), .A2(KEYINPUT29), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n273), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G197gat), .B(G204gat), .ZN(new_n325));
  INV_X1    g124(.A(G218gat), .ZN(new_n326));
  OR2_X1    g125(.A1(KEYINPUT76), .A2(G211gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(KEYINPUT76), .A2(G211gat), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n325), .B1(new_n329), .B2(KEYINPUT22), .ZN(new_n330));
  XNOR2_X1  g129(.A(G211gat), .B(G218gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n325), .B(new_n331), .C1(new_n329), .C2(KEYINPUT22), .ZN(new_n334));
  AND2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n220), .A2(new_n232), .ZN(new_n336));
  NOR3_X1   g135(.A1(new_n336), .A2(new_n270), .A3(new_n321), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n324), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n238), .A2(new_n269), .A3(new_n272), .A4(new_n322), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n323), .B1(new_n336), .B2(new_n270), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n335), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n339), .A2(new_n344), .A3(KEYINPUT77), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n337), .B1(new_n273), .B2(new_n323), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT77), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n346), .A2(new_n347), .A3(new_n335), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G8gat), .B(G36gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(G64gat), .B(G92gat), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n350), .B(new_n351), .Z(new_n352));
  NAND3_X1  g151(.A1(new_n349), .A2(KEYINPUT30), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n352), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n345), .A2(new_n348), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n354), .B1(new_n345), .B2(new_n348), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n357), .A2(KEYINPUT30), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n320), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  XOR2_X1   g158(.A(G78gat), .B(G106gat), .Z(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT83), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT31), .B(G50gat), .ZN(new_n362));
  XOR2_X1   g161(.A(new_n361), .B(new_n362), .Z(new_n363));
  INV_X1    g162(.A(KEYINPUT29), .ZN(new_n364));
  NAND2_X1  g163(.A1(G155gat), .A2(G162gat), .ZN(new_n365));
  NOR2_X1   g164(.A1(G155gat), .A2(G162gat), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  OR2_X1    g166(.A1(G141gat), .A2(G148gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(G141gat), .A2(G148gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n365), .B(new_n367), .C1(new_n370), .C2(KEYINPUT2), .ZN(new_n371));
  XOR2_X1   g170(.A(G141gat), .B(G148gat), .Z(new_n372));
  INV_X1    g171(.A(KEYINPUT79), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT2), .ZN(new_n374));
  AND2_X1   g173(.A1(G155gat), .A2(G162gat), .ZN(new_n375));
  OAI22_X1  g174(.A1(new_n372), .A2(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n367), .A2(KEYINPUT80), .A3(new_n365), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT80), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n378), .B1(new_n375), .B2(new_n366), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n368), .A2(new_n373), .A3(new_n369), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n377), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n371), .B1(new_n376), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n364), .B1(new_n382), .B2(KEYINPUT3), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n335), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT29), .B1(new_n333), .B2(new_n334), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n382), .B1(new_n385), .B2(KEYINPUT3), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT84), .ZN(new_n388));
  INV_X1    g187(.A(G228gat), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n389), .A2(new_n290), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(G22gat), .ZN(new_n392));
  INV_X1    g191(.A(new_n390), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n387), .A2(KEYINPUT84), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n391), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n393), .B1(new_n387), .B2(KEYINPUT84), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT84), .ZN(new_n397));
  AOI211_X1 g196(.A(new_n397), .B(new_n390), .C1(new_n384), .C2(new_n386), .ZN(new_n398));
  OAI21_X1  g197(.A(G22gat), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n363), .B1(new_n395), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT85), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n391), .A2(new_n401), .A3(new_n394), .A4(new_n392), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(new_n399), .A3(new_n363), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n396), .A2(new_n398), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n401), .B1(new_n404), .B2(new_n392), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT86), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n363), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n394), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n407), .B1(new_n408), .B2(G22gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n395), .A2(KEYINPUT85), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT86), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n409), .A2(new_n410), .A3(new_n411), .A4(new_n402), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n400), .B1(new_n406), .B2(new_n412), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n370), .A2(KEYINPUT79), .B1(KEYINPUT2), .B2(new_n365), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n414), .A2(new_n377), .A3(new_n380), .A4(new_n379), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n286), .A2(new_n415), .A3(new_n416), .A4(new_n371), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT81), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n367), .A2(new_n365), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n420), .B1(new_n372), .B2(new_n374), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n377), .A2(new_n379), .A3(new_n380), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n421), .B1(new_n422), .B2(new_n414), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n423), .A2(KEYINPUT81), .A3(new_n416), .A4(new_n286), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT4), .B1(new_n382), .B2(new_n282), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n419), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(G225gat), .A2(G233gat), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT3), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n286), .B1(new_n423), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n382), .A2(KEYINPUT3), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n428), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n426), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT5), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n382), .B(new_n282), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n434), .B1(new_n435), .B2(new_n428), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT5), .B1(new_n425), .B2(new_n417), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n432), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G1gat), .B(G29gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n441), .B(KEYINPUT0), .ZN(new_n442));
  XNOR2_X1  g241(.A(G57gat), .B(G85gat), .ZN(new_n443));
  XOR2_X1   g242(.A(new_n442), .B(new_n443), .Z(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT6), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n433), .A2(new_n436), .B1(new_n432), .B2(new_n438), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n444), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n446), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT82), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n444), .B1(new_n437), .B2(new_n439), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n451), .B1(new_n452), .B2(KEYINPUT6), .ZN(new_n453));
  NOR4_X1   g252(.A1(new_n448), .A2(KEYINPUT82), .A3(new_n447), .A4(new_n444), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n450), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT35), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n413), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n349), .A2(new_n352), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT30), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n461), .A2(KEYINPUT87), .A3(new_n355), .A4(new_n353), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n359), .A2(new_n458), .A3(new_n462), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n318), .A2(new_n319), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n413), .B1(new_n309), .B2(new_n316), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n455), .B1(KEYINPUT30), .B2(new_n357), .ZN(new_n466));
  AOI211_X1 g265(.A(new_n460), .B(new_n354), .C1(new_n345), .C2(new_n348), .ZN(new_n467));
  INV_X1    g266(.A(new_n355), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT78), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT78), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n353), .A2(new_n470), .A3(new_n355), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n466), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n456), .B1(new_n465), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n466), .ZN(new_n474));
  NOR3_X1   g273(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT78), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n470), .B1(new_n353), .B2(new_n355), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n413), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n309), .A2(new_n316), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT36), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n309), .A2(new_n316), .A3(KEYINPUT36), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n478), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n413), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n455), .A2(new_n357), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n354), .A2(KEYINPUT37), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n355), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT37), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n488), .B1(new_n346), .B2(new_n343), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n342), .A2(new_n335), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT38), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n485), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT38), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n345), .A2(KEYINPUT37), .A3(new_n348), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n494), .B1(new_n487), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n484), .B1(new_n493), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n359), .A2(new_n462), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n430), .A2(new_n431), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n425), .A2(new_n417), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n427), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n502), .B(KEYINPUT39), .C1(new_n428), .C2(new_n435), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n503), .B(new_n444), .C1(KEYINPUT39), .C2(new_n502), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n446), .B1(new_n505), .B2(KEYINPUT40), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n506), .B1(KEYINPUT40), .B2(new_n505), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n497), .B1(new_n498), .B2(new_n507), .ZN(new_n508));
  OAI22_X1  g307(.A1(new_n464), .A2(new_n473), .B1(new_n483), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G43gat), .B(G50gat), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  XOR2_X1   g310(.A(KEYINPUT91), .B(KEYINPUT15), .Z(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(G29gat), .A2(G36gat), .ZN(new_n514));
  XOR2_X1   g313(.A(new_n514), .B(KEYINPUT90), .Z(new_n515));
  NAND2_X1  g314(.A1(new_n510), .A2(KEYINPUT15), .ZN(new_n516));
  OR3_X1    g315(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n513), .A2(new_n515), .A3(new_n516), .A4(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n514), .B(KEYINPUT90), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n518), .A2(KEYINPUT89), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n522), .A2(new_n517), .ZN(new_n523));
  OR2_X1    g322(.A1(new_n518), .A2(KEYINPUT89), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n520), .B1(new_n525), .B2(new_n516), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT17), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n524), .A2(new_n517), .A3(new_n522), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(new_n515), .ZN(new_n530));
  INV_X1    g329(.A(new_n516), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n532), .A2(KEYINPUT17), .A3(new_n520), .ZN(new_n533));
  XNOR2_X1  g332(.A(G15gat), .B(G22gat), .ZN(new_n534));
  INV_X1    g333(.A(G1gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT16), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n534), .A2(G1gat), .ZN(new_n539));
  OAI21_X1  g338(.A(G8gat), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n539), .ZN(new_n541));
  INV_X1    g340(.A(G8gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(new_n542), .A3(new_n537), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n528), .A2(new_n533), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G229gat), .A2(G233gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n540), .A2(new_n543), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n526), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT18), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n550), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n544), .A2(new_n532), .A3(new_n520), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(new_n548), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n546), .B(KEYINPUT13), .Z(new_n555));
  AOI21_X1  g354(.A(KEYINPUT92), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n555), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT92), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n551), .B(new_n552), .C1(new_n556), .C2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G113gat), .B(G141gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(G197gat), .ZN(new_n562));
  XOR2_X1   g361(.A(KEYINPUT11), .B(G169gat), .Z(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT12), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n560), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n557), .B(new_n558), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n568), .A2(new_n565), .A3(new_n551), .A4(new_n552), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  AND2_X1   g369(.A1(G232gat), .A2(G233gat), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n571), .A2(KEYINPUT41), .ZN(new_n572));
  XNOR2_X1  g371(.A(G134gat), .B(G162gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G190gat), .B(G218gat), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n576), .A2(KEYINPUT98), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G99gat), .A2(G106gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT8), .ZN(new_n580));
  NAND2_X1  g379(.A1(G85gat), .A2(G92gat), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT7), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(G85gat), .ZN(new_n584));
  INV_X1    g383(.A(G92gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n580), .A2(new_n583), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G99gat), .B(G106gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  AND3_X1   g390(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI22_X1  g393(.A1(KEYINPUT8), .A2(new_n579), .B1(new_n584), .B2(new_n585), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n589), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n528), .A2(new_n533), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT97), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n597), .B1(new_n526), .B2(new_n527), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT97), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n601), .A2(new_n602), .A3(new_n533), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n526), .A2(new_n597), .ZN(new_n605));
  AOI22_X1  g404(.A1(new_n576), .A2(KEYINPUT98), .B1(KEYINPUT41), .B2(new_n571), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n578), .B1(new_n604), .B2(new_n608), .ZN(new_n609));
  AOI211_X1 g408(.A(new_n577), .B(new_n607), .C1(new_n600), .C2(new_n603), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n575), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n603), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n602), .B1(new_n601), .B2(new_n533), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n608), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n577), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n604), .A2(new_n578), .A3(new_n608), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(new_n574), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G71gat), .B(G78gat), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n622));
  AND2_X1   g421(.A1(G57gat), .A2(G64gat), .ZN(new_n623));
  NOR2_X1   g422(.A1(G57gat), .A2(G64gat), .ZN(new_n624));
  NOR3_X1   g423(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G71gat), .A2(G78gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT93), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n621), .B1(new_n625), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT9), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  OR2_X1    g430(.A1(G57gat), .A2(G64gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(G57gat), .A2(G64gat), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n634), .A2(new_n620), .A3(new_n627), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n629), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n636), .A2(KEYINPUT21), .ZN(new_n637));
  XOR2_X1   g436(.A(G127gat), .B(G155gat), .Z(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT96), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n637), .B(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n547), .B1(KEYINPUT21), .B2(new_n636), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n640), .B(new_n641), .Z(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT20), .ZN(new_n644));
  NAND2_X1  g443(.A1(G231gat), .A2(G233gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT94), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n644), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G183gat), .B(G211gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n642), .B(new_n649), .Z(new_n650));
  NOR2_X1   g449(.A1(new_n619), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n594), .A2(new_n589), .A3(new_n595), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n588), .A2(new_n590), .ZN(new_n654));
  AND3_X1   g453(.A1(new_n634), .A2(new_n620), .A3(new_n627), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n620), .B1(new_n634), .B2(new_n627), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n653), .B(new_n654), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n629), .B(new_n635), .C1(new_n591), .C2(new_n596), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT10), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT99), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n597), .A2(new_n636), .A3(KEYINPUT10), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n657), .A2(new_n658), .A3(KEYINPUT99), .A4(new_n659), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(G230gat), .A2(G233gat), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n652), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n666), .B1(new_n657), .B2(new_n658), .ZN(new_n669));
  XNOR2_X1  g468(.A(G120gat), .B(G148gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT101), .ZN(new_n671));
  XNOR2_X1  g470(.A(G176gat), .B(G204gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n665), .A2(new_n652), .A3(new_n666), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n668), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n665), .A2(new_n666), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n673), .B1(new_n678), .B2(new_n669), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  AND4_X1   g480(.A1(new_n509), .A2(new_n570), .A3(new_n651), .A4(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n455), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g484(.A1(new_n682), .A2(new_n498), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT16), .B(G8gat), .Z(new_n687));
  AND2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n686), .A2(new_n542), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT42), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(KEYINPUT42), .B2(new_n688), .ZN(G1325gat));
  INV_X1    g490(.A(G15gat), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n318), .A2(new_n319), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n682), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n481), .A2(new_n482), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n682), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n694), .B1(new_n697), .B2(new_n692), .ZN(G1326gat));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n413), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT43), .B(G22gat), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1327gat));
  NAND2_X1  g500(.A1(new_n509), .A2(new_n619), .ZN(new_n702));
  INV_X1    g501(.A(new_n650), .ZN(new_n703));
  INV_X1    g502(.A(new_n570), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n703), .A2(new_n704), .A3(new_n680), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n708), .A2(G29gat), .A3(new_n455), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(KEYINPUT45), .Z(new_n710));
  INV_X1    g509(.A(KEYINPUT103), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n483), .A2(new_n508), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n359), .A2(new_n458), .A3(new_n462), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT88), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n479), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n714), .A2(new_n716), .A3(new_n317), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n479), .A2(new_n472), .A3(new_n484), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT35), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT102), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n717), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n720), .B1(new_n717), .B2(new_n719), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n713), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n618), .A2(KEYINPUT44), .ZN(new_n724));
  AOI22_X1  g523(.A1(new_n723), .A2(new_n724), .B1(new_n702), .B2(KEYINPUT44), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n711), .B1(new_n725), .B2(new_n706), .ZN(new_n726));
  INV_X1    g525(.A(new_n724), .ZN(new_n727));
  OAI21_X1  g526(.A(KEYINPUT102), .B1(new_n464), .B2(new_n473), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n717), .A2(new_n719), .A3(new_n720), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n727), .B1(new_n730), .B2(new_n713), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n732), .B1(new_n509), .B2(new_n619), .ZN(new_n733));
  OAI211_X1 g532(.A(KEYINPUT103), .B(new_n705), .C1(new_n731), .C2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n726), .A2(new_n683), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(G29gat), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n710), .A2(new_n736), .ZN(G1328gat));
  NAND3_X1  g536(.A1(new_n726), .A2(new_n498), .A3(new_n734), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(G36gat), .ZN(new_n739));
  INV_X1    g538(.A(G36gat), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n707), .A2(new_n740), .A3(new_n498), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n741), .B(KEYINPUT46), .Z(new_n742));
  NAND2_X1  g541(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT104), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n739), .A2(new_n742), .A3(KEYINPUT104), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(G1329gat));
  INV_X1    g546(.A(new_n725), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n705), .ZN(new_n749));
  OAI21_X1  g548(.A(G43gat), .B1(new_n749), .B2(new_n695), .ZN(new_n750));
  INV_X1    g549(.A(new_n693), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n708), .A2(G43gat), .A3(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n750), .A2(KEYINPUT47), .A3(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n726), .A2(new_n696), .A3(new_n734), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n752), .B1(new_n755), .B2(G43gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n756), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g556(.A(G50gat), .B1(new_n749), .B2(new_n484), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n708), .A2(G50gat), .A3(new_n484), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n758), .A2(KEYINPUT48), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n726), .A2(new_n413), .A3(new_n734), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n759), .B1(new_n762), .B2(G50gat), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n763), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR4_X1   g563(.A1(new_n650), .A2(new_n619), .A3(new_n570), .A4(new_n681), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n723), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n455), .B(KEYINPUT105), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G57gat), .ZN(G1332gat));
  INV_X1    g568(.A(KEYINPUT49), .ZN(new_n770));
  INV_X1    g569(.A(G64gat), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n498), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT106), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n766), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n770), .A2(new_n771), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n774), .B(new_n775), .ZN(G1333gat));
  NAND3_X1  g575(.A1(new_n766), .A2(KEYINPUT107), .A3(new_n693), .ZN(new_n777));
  INV_X1    g576(.A(G71gat), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT107), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n723), .A2(new_n765), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n780), .B2(new_n751), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n777), .A2(new_n778), .A3(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n766), .A2(G71gat), .A3(new_n696), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n785));
  XOR2_X1   g584(.A(new_n784), .B(new_n785), .Z(G1334gat));
  NAND2_X1  g585(.A1(new_n766), .A2(new_n413), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g587(.A1(new_n703), .A2(new_n570), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n790), .A2(new_n681), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n725), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(G85gat), .B1(new_n794), .B2(new_n455), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n790), .A2(new_n618), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n723), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n723), .A2(KEYINPUT51), .A3(new_n796), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT109), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n681), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n803), .B1(new_n802), .B2(new_n801), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n683), .A2(new_n584), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n795), .B1(new_n804), .B2(new_n805), .ZN(G1336gat));
  INV_X1    g605(.A(new_n498), .ZN(new_n807));
  OAI21_X1  g606(.A(G92gat), .B1(new_n794), .B2(new_n807), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n801), .A2(new_n585), .A3(new_n498), .A4(new_n680), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT52), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n808), .A2(new_n812), .A3(new_n809), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(G1337gat));
  OAI21_X1  g613(.A(G99gat), .B1(new_n794), .B2(new_n695), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n693), .A2(new_n301), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n815), .B1(new_n804), .B2(new_n816), .ZN(G1338gat));
  INV_X1    g616(.A(G106gat), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n818), .B1(new_n793), .B2(new_n413), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n484), .A2(G106gat), .A3(new_n681), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n821), .B1(new_n799), .B2(new_n800), .ZN(new_n822));
  OAI21_X1  g621(.A(KEYINPUT53), .B1(new_n819), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT110), .ZN(new_n824));
  INV_X1    g623(.A(new_n819), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT53), .B1(new_n822), .B2(KEYINPUT111), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n825), .B(new_n826), .C1(KEYINPUT111), .C2(new_n822), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT110), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n828), .B(KEYINPUT53), .C1(new_n819), .C2(new_n822), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n824), .A2(new_n827), .A3(new_n829), .ZN(G1339gat));
  AND3_X1   g629(.A1(new_n665), .A2(new_n652), .A3(new_n666), .ZN(new_n831));
  INV_X1    g630(.A(new_n666), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n662), .A2(new_n832), .A3(new_n663), .A4(new_n664), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT54), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n831), .A2(new_n667), .A3(new_n834), .ZN(new_n835));
  OAI211_X1 g634(.A(KEYINPUT55), .B(new_n673), .C1(new_n677), .C2(KEYINPUT54), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n676), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT112), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI211_X1 g638(.A(KEYINPUT112), .B(new_n676), .C1(new_n835), .C2(new_n836), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n673), .B1(new_n677), .B2(KEYINPUT54), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n841), .B1(new_n835), .B2(new_n842), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n839), .A2(new_n570), .A3(new_n840), .A4(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT114), .B1(new_n554), .B2(new_n555), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT114), .ZN(new_n846));
  INV_X1    g645(.A(new_n555), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n553), .A2(new_n548), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n546), .B1(new_n545), .B2(new_n548), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n845), .B(new_n848), .C1(new_n849), .C2(KEYINPUT113), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n849), .A2(KEYINPUT113), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n564), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n680), .A2(new_n569), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n844), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n618), .ZN(new_n855));
  AND4_X1   g654(.A1(new_n569), .A2(new_n611), .A3(new_n617), .A4(new_n852), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n856), .A2(new_n839), .A3(new_n840), .A4(new_n843), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(KEYINPUT115), .A3(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT115), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n619), .B1(new_n844), .B2(new_n853), .ZN(new_n860));
  INV_X1    g659(.A(new_n857), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n858), .A2(new_n650), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n651), .A2(new_n704), .A3(new_n681), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n863), .A2(KEYINPUT116), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT116), .B1(new_n863), .B2(new_n864), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n867), .A2(new_n767), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(new_n465), .A3(new_n807), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(G113gat), .B1(new_n870), .B2(new_n570), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n863), .A2(new_n864), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT116), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n863), .A2(KEYINPUT116), .A3(new_n864), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(new_n484), .A3(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT117), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n874), .A2(KEYINPUT117), .A3(new_n484), .A4(new_n875), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n498), .A2(new_n455), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n880), .A2(new_n693), .A3(new_n881), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n570), .A2(G113gat), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n871), .B1(new_n882), .B2(new_n883), .ZN(G1340gat));
  AND2_X1   g683(.A1(new_n882), .A2(new_n680), .ZN(new_n885));
  INV_X1    g684(.A(G120gat), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n680), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT118), .ZN(new_n888));
  OAI22_X1  g687(.A1(new_n885), .A2(new_n886), .B1(new_n869), .B2(new_n888), .ZN(G1341gat));
  NOR2_X1   g688(.A1(new_n869), .A2(new_n650), .ZN(new_n890));
  OR2_X1    g689(.A1(new_n890), .A2(KEYINPUT119), .ZN(new_n891));
  AOI21_X1  g690(.A(G127gat), .B1(new_n890), .B2(KEYINPUT119), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n703), .A2(G127gat), .ZN(new_n893));
  AOI22_X1  g692(.A1(new_n891), .A2(new_n892), .B1(new_n882), .B2(new_n893), .ZN(G1342gat));
  NOR3_X1   g693(.A1(new_n869), .A2(G134gat), .A3(new_n618), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT56), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n882), .A2(new_n619), .ZN(new_n897));
  INV_X1    g696(.A(G134gat), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(G1343gat));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n835), .A2(new_n836), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n570), .A2(new_n676), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n835), .A2(new_n842), .ZN(new_n903));
  XNOR2_X1  g702(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n853), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI211_X1 g707(.A(KEYINPUT121), .B(new_n853), .C1(new_n902), .C2(new_n905), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n618), .A3(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n861), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n908), .A2(KEYINPUT122), .A3(new_n618), .A4(new_n909), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n864), .B1(new_n914), .B2(new_n703), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT57), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n484), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n874), .A2(new_n413), .A3(new_n875), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n915), .A2(new_n917), .B1(new_n918), .B2(new_n916), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n695), .A2(new_n881), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n900), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n915), .A2(new_n917), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n918), .A2(new_n916), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(new_n920), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n924), .A2(KEYINPUT123), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n921), .A2(new_n926), .A3(new_n570), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n696), .A2(new_n484), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n867), .A2(new_n807), .A3(new_n767), .A4(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n704), .A2(G141gat), .ZN(new_n931));
  AOI22_X1  g730(.A1(new_n927), .A2(G141gat), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT58), .ZN(new_n933));
  INV_X1    g732(.A(new_n931), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n933), .B1(new_n929), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n924), .A2(new_n570), .A3(new_n925), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n935), .B1(new_n936), .B2(G141gat), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n937), .A2(KEYINPUT124), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT124), .ZN(new_n939));
  AOI211_X1 g738(.A(new_n939), .B(new_n935), .C1(new_n936), .C2(G141gat), .ZN(new_n940));
  OAI22_X1  g739(.A1(new_n932), .A2(new_n933), .B1(new_n938), .B2(new_n940), .ZN(G1344gat));
  INV_X1    g740(.A(KEYINPUT59), .ZN(new_n942));
  AOI211_X1 g741(.A(new_n942), .B(G148gat), .C1(new_n930), .C2(new_n680), .ZN(new_n943));
  INV_X1    g742(.A(G148gat), .ZN(new_n944));
  INV_X1    g743(.A(new_n864), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n910), .A2(new_n857), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n945), .B1(new_n946), .B2(new_n650), .ZN(new_n947));
  OR2_X1    g746(.A1(new_n947), .A2(new_n484), .ZN(new_n948));
  AOI22_X1  g747(.A1(new_n867), .A2(new_n917), .B1(new_n948), .B2(new_n916), .ZN(new_n949));
  OR3_X1    g748(.A1(new_n949), .A2(new_n681), .A3(new_n920), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n944), .B1(new_n950), .B2(KEYINPUT59), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n921), .A2(new_n926), .A3(new_n942), .A4(new_n680), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n943), .B1(new_n951), .B2(new_n952), .ZN(G1345gat));
  INV_X1    g752(.A(G155gat), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n930), .A2(new_n954), .A3(new_n703), .ZN(new_n955));
  AND3_X1   g754(.A1(new_n921), .A2(new_n926), .A3(new_n703), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n955), .B1(new_n956), .B2(new_n954), .ZN(G1346gat));
  INV_X1    g756(.A(G162gat), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n930), .A2(new_n958), .A3(new_n619), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n921), .A2(new_n926), .A3(new_n619), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n959), .B1(new_n960), .B2(new_n958), .ZN(G1347gat));
  NOR4_X1   g760(.A1(new_n865), .A2(new_n866), .A3(new_n683), .A4(new_n807), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n962), .A2(new_n465), .ZN(new_n963));
  AOI21_X1  g762(.A(G169gat), .B1(new_n963), .B2(new_n570), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n807), .A2(new_n767), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n693), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n966), .B1(new_n878), .B2(new_n879), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n704), .A2(new_n252), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(G1348gat));
  INV_X1    g768(.A(new_n967), .ZN(new_n970));
  OAI21_X1  g769(.A(G176gat), .B1(new_n970), .B2(new_n681), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n963), .A2(new_n253), .A3(new_n680), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(G1349gat));
  INV_X1    g772(.A(new_n966), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT117), .B1(new_n867), .B2(new_n484), .ZN(new_n975));
  INV_X1    g774(.A(new_n879), .ZN(new_n976));
  OAI211_X1 g775(.A(new_n703), .B(new_n974), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(KEYINPUT125), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT125), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n967), .A2(new_n979), .A3(new_n703), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n978), .A2(G183gat), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n205), .A2(KEYINPUT27), .ZN(new_n982));
  NAND4_X1  g781(.A1(new_n963), .A2(new_n208), .A3(new_n982), .A4(new_n703), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(KEYINPUT60), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT60), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n981), .A2(new_n986), .A3(new_n983), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n985), .A2(new_n987), .ZN(G1350gat));
  NAND3_X1  g787(.A1(new_n963), .A2(new_n245), .A3(new_n619), .ZN(new_n989));
  AOI211_X1 g788(.A(new_n618), .B(new_n966), .C1(new_n878), .C2(new_n879), .ZN(new_n990));
  OAI21_X1  g789(.A(KEYINPUT126), .B1(new_n990), .B2(new_n245), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n967), .A2(new_n619), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT126), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n992), .A2(new_n993), .A3(G190gat), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT61), .ZN(new_n995));
  AND3_X1   g794(.A1(new_n991), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n995), .B1(new_n991), .B2(new_n994), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n989), .B1(new_n996), .B2(new_n997), .ZN(G1351gat));
  NAND2_X1  g797(.A1(new_n962), .A2(new_n928), .ZN(new_n999));
  XNOR2_X1  g798(.A(new_n999), .B(KEYINPUT127), .ZN(new_n1000));
  AOI21_X1  g799(.A(G197gat), .B1(new_n1000), .B2(new_n570), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n695), .A2(new_n965), .ZN(new_n1002));
  NOR2_X1   g801(.A1(new_n949), .A2(new_n1002), .ZN(new_n1003));
  AND2_X1   g802(.A1(new_n570), .A2(G197gat), .ZN(new_n1004));
  AOI21_X1  g803(.A(new_n1001), .B1(new_n1003), .B2(new_n1004), .ZN(G1352gat));
  NOR3_X1   g804(.A1(new_n999), .A2(G204gat), .A3(new_n681), .ZN(new_n1006));
  XNOR2_X1  g805(.A(new_n1006), .B(KEYINPUT62), .ZN(new_n1007));
  INV_X1    g806(.A(G204gat), .ZN(new_n1008));
  NOR3_X1   g807(.A1(new_n949), .A2(new_n681), .A3(new_n1002), .ZN(new_n1009));
  OAI21_X1  g808(.A(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(G1353gat));
  NAND4_X1  g809(.A1(new_n1000), .A2(new_n327), .A3(new_n328), .A4(new_n703), .ZN(new_n1011));
  INV_X1    g810(.A(G211gat), .ZN(new_n1012));
  AOI21_X1  g811(.A(new_n1012), .B1(new_n1003), .B2(new_n703), .ZN(new_n1013));
  AND2_X1   g812(.A1(new_n1013), .A2(KEYINPUT63), .ZN(new_n1014));
  NOR2_X1   g813(.A1(new_n1013), .A2(KEYINPUT63), .ZN(new_n1015));
  OAI21_X1  g814(.A(new_n1011), .B1(new_n1014), .B2(new_n1015), .ZN(G1354gat));
  NAND3_X1  g815(.A1(new_n1000), .A2(new_n326), .A3(new_n619), .ZN(new_n1017));
  NOR3_X1   g816(.A1(new_n949), .A2(new_n618), .A3(new_n1002), .ZN(new_n1018));
  OAI21_X1  g817(.A(new_n1017), .B1(new_n326), .B2(new_n1018), .ZN(G1355gat));
endmodule


