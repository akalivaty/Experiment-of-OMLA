//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 1 1 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 1 1 1 1 0 0 0 1 1 1 0 1 0 1 0 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT9), .B(G234), .Z(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT77), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G469), .ZN(new_n193));
  XNOR2_X1  g007(.A(G110), .B(G140), .ZN(new_n194));
  INV_X1    g008(.A(G953), .ZN(new_n195));
  AND2_X1   g009(.A1(new_n195), .A2(G227), .ZN(new_n196));
  XNOR2_X1  g010(.A(new_n194), .B(new_n196), .ZN(new_n197));
  XOR2_X1   g011(.A(KEYINPUT81), .B(KEYINPUT10), .Z(new_n198));
  INV_X1    g012(.A(G104), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT3), .B1(new_n199), .B2(G107), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G104), .ZN(new_n203));
  INV_X1    g017(.A(G101), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n199), .A2(G107), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n200), .A2(new_n203), .A3(new_n204), .A4(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n202), .A2(G104), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n199), .A2(G107), .ZN(new_n208));
  OAI21_X1  g022(.A(G101), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AND2_X1   g023(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(G143), .B(G146), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT1), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(G128), .ZN(new_n213));
  INV_X1    g027(.A(G143), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT1), .B1(new_n214), .B2(G146), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G143), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n214), .A2(G146), .ZN(new_n218));
  AOI22_X1  g032(.A1(new_n215), .A2(G128), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT79), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n213), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G128), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n222), .B1(new_n217), .B2(KEYINPUT1), .ZN(new_n223));
  NOR3_X1   g037(.A1(new_n223), .A2(new_n211), .A3(KEYINPUT79), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n210), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT80), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT79), .B1(new_n223), .B2(new_n211), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n215), .A2(G128), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n217), .A2(new_n218), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(new_n220), .A3(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n227), .A2(new_n230), .A3(new_n213), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT80), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n232), .A3(new_n210), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n198), .B1(new_n226), .B2(new_n233), .ZN(new_n234));
  OAI211_X1 g048(.A(KEYINPUT66), .B(KEYINPUT1), .C1(new_n214), .C2(G146), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G128), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT66), .B1(new_n217), .B2(KEYINPUT1), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n229), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n213), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n210), .A2(KEYINPUT10), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n238), .A2(KEYINPUT68), .A3(new_n213), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n200), .A2(new_n203), .A3(new_n205), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G101), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n246), .A2(KEYINPUT4), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n211), .A2(KEYINPUT0), .A3(G128), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT0), .B(G128), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n248), .B1(new_n211), .B2(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n246), .A2(KEYINPUT78), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n206), .A2(KEYINPUT4), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT78), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n245), .A2(new_n254), .A3(G101), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n252), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n251), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n244), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT11), .ZN(new_n259));
  INV_X1    g073(.A(G134), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n259), .B1(new_n260), .B2(G137), .ZN(new_n261));
  INV_X1    g075(.A(G137), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n262), .A2(KEYINPUT11), .A3(G134), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n260), .A2(G137), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n261), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  AND2_X1   g079(.A1(KEYINPUT65), .A2(G131), .ZN(new_n266));
  OR2_X1    g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n266), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NOR3_X1   g083(.A1(new_n234), .A2(new_n258), .A3(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n269), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n238), .A2(KEYINPUT68), .A3(new_n213), .ZN(new_n272));
  AOI21_X1  g086(.A(KEYINPUT68), .B1(new_n238), .B2(new_n213), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n274), .A2(new_n242), .B1(new_n256), .B2(new_n251), .ZN(new_n275));
  INV_X1    g089(.A(new_n198), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n231), .A2(new_n232), .A3(new_n210), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n232), .B1(new_n231), .B2(new_n210), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n271), .B1(new_n275), .B2(new_n279), .ZN(new_n280));
  OAI211_X1 g094(.A(KEYINPUT83), .B(new_n197), .C1(new_n270), .C2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n197), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n275), .A2(new_n271), .A3(new_n279), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n239), .A2(new_n210), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n284), .B1(new_n226), .B2(new_n233), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT12), .ZN(new_n286));
  NOR3_X1   g100(.A1(new_n285), .A2(new_n286), .A3(new_n271), .ZN(new_n287));
  INV_X1    g101(.A(new_n284), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n288), .B1(new_n277), .B2(new_n278), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT12), .B1(new_n289), .B2(new_n269), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n282), .B(new_n283), .C1(new_n287), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n281), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n269), .B1(new_n234), .B2(new_n258), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n283), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT83), .B1(new_n294), .B2(new_n197), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n193), .B(new_n190), .C1(new_n292), .C2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(G469), .A2(G902), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n283), .B1(new_n287), .B2(new_n290), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT82), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT82), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n301), .B(new_n283), .C1(new_n287), .C2(new_n290), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n282), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  NOR3_X1   g117(.A1(new_n270), .A2(new_n280), .A3(new_n197), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n303), .A2(new_n193), .A3(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n192), .B1(new_n298), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT84), .ZN(new_n307));
  INV_X1    g121(.A(new_n302), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n286), .B1(new_n285), .B2(new_n271), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n289), .A2(KEYINPUT12), .A3(new_n269), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n301), .B1(new_n311), .B2(new_n283), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n197), .B1(new_n308), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n304), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(G469), .A3(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(new_n296), .A3(new_n297), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT84), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n317), .A3(new_n192), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT20), .ZN(new_n319));
  NOR2_X1   g133(.A1(G475), .A2(G902), .ZN(new_n320));
  XNOR2_X1  g134(.A(G125), .B(G140), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT16), .ZN(new_n322));
  INV_X1    g136(.A(G125), .ZN(new_n323));
  OR3_X1    g137(.A1(new_n323), .A2(KEYINPUT16), .A3(G140), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n216), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n322), .A2(G146), .A3(new_n324), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G237), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(new_n195), .A3(G214), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n330), .B(new_n214), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(KEYINPUT17), .A3(G131), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT88), .B1(new_n331), .B2(G131), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(G131), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n330), .B(G143), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT88), .ZN(new_n336));
  INV_X1    g150(.A(G131), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n333), .A2(new_n334), .A3(new_n338), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n328), .B(new_n332), .C1(new_n339), .C2(KEYINPUT17), .ZN(new_n340));
  XNOR2_X1  g154(.A(G113), .B(G122), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(G104), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT18), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n335), .B1(new_n344), .B2(new_n337), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n331), .A2(KEYINPUT18), .A3(G131), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n321), .B(new_n216), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n340), .A2(new_n343), .A3(new_n348), .ZN(new_n349));
  XOR2_X1   g163(.A(new_n321), .B(KEYINPUT19), .Z(new_n350));
  OR2_X1    g164(.A1(new_n350), .A2(G146), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(new_n339), .A3(new_n327), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n343), .B1(new_n352), .B2(new_n348), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n319), .B(new_n320), .C1(new_n349), .C2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT89), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n352), .A2(new_n348), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n342), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n340), .A2(new_n343), .A3(new_n348), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n360), .A2(KEYINPUT89), .A3(new_n319), .A4(new_n320), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n320), .B1(new_n349), .B2(new_n353), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(KEYINPUT20), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n356), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n343), .B1(new_n340), .B2(new_n348), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n190), .B1(new_n349), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G475), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n189), .A2(G217), .A3(new_n195), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n214), .A2(G128), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n222), .A2(G143), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n371), .A2(new_n372), .A3(new_n260), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n260), .B1(new_n371), .B2(new_n372), .ZN(new_n374));
  OR2_X1    g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(G116), .B(G122), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT14), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G116), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(KEYINPUT14), .A3(G122), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(G107), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n376), .A2(new_n202), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n375), .A2(KEYINPUT90), .A3(new_n381), .A4(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n376), .B(new_n202), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT13), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n371), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n372), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n371), .A2(new_n385), .ZN(new_n388));
  OAI21_X1  g202(.A(G134), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n373), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n384), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT90), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n378), .A2(G107), .A3(new_n380), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n382), .B1(new_n373), .B2(new_n374), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n370), .A2(new_n383), .A3(new_n391), .A4(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(new_n383), .A3(new_n391), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n369), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n396), .A2(new_n398), .A3(KEYINPUT91), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT91), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n397), .A2(new_n400), .A3(new_n369), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n190), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G478), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(KEYINPUT15), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n402), .B(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n368), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(G214), .B1(G237), .B2(G902), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(G116), .B(G119), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(KEYINPUT2), .B(G113), .ZN(new_n411));
  NOR3_X1   g225(.A1(new_n410), .A2(KEYINPUT67), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT67), .ZN(new_n413));
  XOR2_X1   g227(.A(KEYINPUT2), .B(G113), .Z(new_n414));
  AOI21_X1  g228(.A(new_n413), .B1(new_n414), .B2(new_n409), .ZN(new_n415));
  OAI22_X1  g229(.A1(new_n412), .A2(new_n415), .B1(new_n409), .B2(new_n414), .ZN(new_n416));
  INV_X1    g230(.A(new_n247), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n416), .A2(new_n256), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n415), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n414), .A2(new_n413), .A3(new_n409), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT5), .ZN(new_n422));
  INV_X1    g236(.A(G119), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n423), .A3(G116), .ZN(new_n424));
  OAI211_X1 g238(.A(G113), .B(new_n424), .C1(new_n410), .C2(new_n422), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n421), .A2(new_n210), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n418), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT6), .ZN(new_n428));
  XNOR2_X1  g242(.A(G110), .B(G122), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n427), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n418), .A2(new_n429), .A3(new_n426), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT6), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n429), .B1(new_n418), .B2(new_n426), .ZN(new_n434));
  OAI211_X1 g248(.A(KEYINPUT85), .B(new_n431), .C1(new_n433), .C2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n434), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT85), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n436), .A2(new_n437), .A3(KEYINPUT6), .A4(new_n432), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n239), .A2(new_n323), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n440), .B1(new_n323), .B2(new_n250), .ZN(new_n441));
  INV_X1    g255(.A(G224), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(G953), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n441), .B(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n439), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G210), .B1(G237), .B2(G902), .ZN(new_n447));
  OAI21_X1  g261(.A(KEYINPUT7), .B1(new_n442), .B2(G953), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  OR2_X1    g263(.A1(new_n441), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n421), .A2(new_n425), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT86), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n452), .A3(new_n210), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n210), .A2(new_n452), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n421), .A2(new_n454), .A3(new_n425), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n429), .B(KEYINPUT8), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n453), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n450), .A2(new_n457), .A3(new_n432), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n441), .A2(new_n449), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(KEYINPUT87), .ZN(new_n461));
  AOI21_X1  g275(.A(G902), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n446), .A2(new_n447), .A3(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n447), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n444), .B1(new_n435), .B2(new_n438), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT87), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n460), .B(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n190), .B1(new_n467), .B2(new_n458), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n464), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n408), .B1(new_n463), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n195), .A2(G952), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n472), .B1(G234), .B2(G237), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(G234), .ZN(new_n475));
  OAI211_X1 g289(.A(G902), .B(G953), .C1(new_n475), .C2(new_n329), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n476), .B(KEYINPUT92), .ZN(new_n477));
  XOR2_X1   g291(.A(KEYINPUT21), .B(G898), .Z(new_n478));
  OAI21_X1  g292(.A(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n479), .B(KEYINPUT93), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n406), .A2(new_n470), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n307), .A2(new_n318), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT94), .ZN(new_n483));
  INV_X1    g297(.A(G217), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n484), .B1(G234), .B2(new_n190), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n321), .A2(new_n216), .ZN(new_n486));
  AOI21_X1  g300(.A(KEYINPUT73), .B1(new_n222), .B2(G119), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT23), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n488), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n423), .A2(G128), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT74), .B(G110), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n222), .A2(G119), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n491), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT24), .B(G110), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  XOR2_X1   g312(.A(new_n498), .B(KEYINPUT75), .Z(new_n499));
  OAI211_X1 g313(.A(new_n327), .B(new_n486), .C1(new_n494), .C2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n326), .A2(new_n327), .ZN(new_n501));
  INV_X1    g315(.A(G110), .ZN(new_n502));
  OAI221_X1 g316(.A(new_n501), .B1(new_n502), .B2(new_n492), .C1(new_n496), .C2(new_n497), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT22), .B(G137), .ZN(new_n505));
  NOR3_X1   g319(.A1(new_n187), .A2(new_n475), .A3(G953), .ZN(new_n506));
  XOR2_X1   g320(.A(new_n505), .B(new_n506), .Z(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n507), .B1(new_n500), .B2(new_n503), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(KEYINPUT25), .B1(new_n511), .B2(new_n190), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT25), .ZN(new_n513));
  NOR4_X1   g327(.A1(new_n509), .A2(new_n510), .A3(new_n513), .A4(G902), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n485), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n485), .A2(G902), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(KEYINPUT76), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n511), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n265), .A2(new_n337), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n262), .A2(G134), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n522), .A2(new_n264), .A3(G131), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n241), .A2(new_n524), .A3(new_n243), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n250), .B1(new_n268), .B2(new_n267), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n525), .A2(KEYINPUT30), .A3(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n529));
  AND2_X1   g343(.A1(new_n238), .A2(new_n213), .ZN(new_n530));
  INV_X1    g344(.A(new_n524), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n529), .B1(new_n532), .B2(new_n526), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n528), .A2(new_n533), .A3(new_n416), .ZN(new_n534));
  INV_X1    g348(.A(new_n416), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n525), .A2(new_n535), .A3(new_n527), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT26), .B(G101), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n329), .A2(new_n195), .A3(G210), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n540), .B(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT29), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n416), .B1(new_n532), .B2(new_n526), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n536), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT28), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT28), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n536), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT70), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT70), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n536), .A2(new_n550), .A3(new_n547), .ZN(new_n551));
  INV_X1    g365(.A(new_n542), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n546), .A2(new_n549), .A3(new_n551), .A4(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n543), .A2(new_n553), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n536), .A2(KEYINPUT71), .ZN(new_n555));
  NOR3_X1   g369(.A1(new_n272), .A2(new_n273), .A3(new_n531), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n416), .B1(new_n556), .B2(new_n526), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT71), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n525), .A2(new_n558), .A3(new_n527), .A4(new_n535), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT28), .B1(new_n555), .B2(new_n560), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n536), .A2(new_n550), .A3(new_n547), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n550), .B1(new_n536), .B2(new_n547), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n552), .A2(KEYINPUT29), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n561), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n554), .A2(new_n190), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G472), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT32), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n534), .A2(new_n536), .A3(new_n552), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT31), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n534), .A2(KEYINPUT31), .A3(new_n536), .A4(new_n552), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n546), .A2(new_n549), .A3(new_n551), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n572), .A2(new_n573), .B1(new_n574), .B2(new_n542), .ZN(new_n575));
  NOR2_X1   g389(.A1(G472), .A2(G902), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n569), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n572), .A2(new_n573), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n574), .A2(new_n542), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n581), .A2(KEYINPUT32), .A3(new_n576), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n568), .A2(new_n578), .A3(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT72), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n568), .A2(new_n578), .A3(new_n582), .A4(KEYINPUT72), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n520), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT94), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n307), .A2(new_n588), .A3(new_n318), .A4(new_n481), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n483), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(G101), .ZN(G3));
  AND3_X1   g405(.A1(new_n316), .A2(new_n317), .A3(new_n192), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n317), .B1(new_n316), .B2(new_n192), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT96), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n463), .A2(new_n469), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n596), .A2(new_n407), .A3(new_n480), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n402), .A2(new_n403), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT95), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n402), .A2(KEYINPUT95), .A3(new_n403), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT33), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n399), .A2(new_n602), .A3(new_n401), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n396), .A2(new_n398), .A3(KEYINPUT33), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n403), .A2(G902), .ZN(new_n606));
  AOI22_X1  g420(.A1(new_n600), .A2(new_n601), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n368), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n595), .B1(new_n597), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n607), .B1(new_n367), .B2(new_n364), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n611), .A2(new_n470), .A3(KEYINPUT96), .A4(new_n480), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(G472), .B1(new_n575), .B2(G902), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n614), .B1(new_n575), .B2(new_n577), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n615), .A2(new_n520), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n594), .A2(new_n613), .A3(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT34), .B(G104), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G6));
  AOI21_X1  g433(.A(new_n319), .B1(new_n360), .B2(new_n320), .ZN(new_n620));
  INV_X1    g434(.A(new_n320), .ZN(new_n621));
  AOI211_X1 g435(.A(KEYINPUT20), .B(new_n621), .C1(new_n358), .C2(new_n359), .ZN(new_n622));
  OAI21_X1  g436(.A(KEYINPUT97), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT97), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n363), .A2(new_n624), .A3(new_n354), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n626), .A2(new_n367), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n405), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n628), .A2(new_n597), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n594), .A2(new_n616), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT35), .B(G107), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G9));
  NOR2_X1   g446(.A1(new_n508), .A2(KEYINPUT36), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n504), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n517), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n615), .B1(new_n515), .B2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n483), .A2(new_n589), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT37), .B(G110), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G12));
  NAND2_X1  g453(.A1(new_n515), .A2(new_n635), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n470), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n585), .B2(new_n586), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n477), .A2(G900), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n473), .ZN(new_n644));
  XOR2_X1   g458(.A(new_n644), .B(KEYINPUT98), .Z(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n626), .A2(new_n405), .A3(new_n367), .A4(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n594), .A2(new_n642), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G128), .ZN(G30));
  XOR2_X1   g464(.A(new_n645), .B(KEYINPUT39), .Z(new_n651));
  NAND2_X1  g465(.A1(new_n594), .A2(new_n651), .ZN(new_n652));
  OR2_X1    g466(.A1(new_n652), .A2(KEYINPUT40), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(KEYINPUT40), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n655));
  XOR2_X1   g469(.A(new_n596), .B(new_n655), .Z(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n555), .A2(new_n560), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n570), .B1(new_n658), .B2(new_n552), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n190), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(G472), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n578), .A2(new_n582), .A3(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n663), .A2(new_n640), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n368), .A2(new_n405), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  AND4_X1   g480(.A1(new_n407), .A2(new_n657), .A3(new_n664), .A4(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n653), .A2(new_n654), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G143), .ZN(G45));
  NAND3_X1  g483(.A1(new_n608), .A2(new_n368), .A3(new_n646), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n642), .A2(new_n307), .A3(new_n318), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G146), .ZN(G48));
  OAI21_X1  g487(.A(new_n190), .B1(new_n292), .B2(new_n295), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(G469), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n675), .A2(new_n192), .A3(new_n296), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(KEYINPUT100), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT100), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n675), .A2(new_n678), .A3(new_n192), .A4(new_n296), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n613), .A2(new_n587), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT41), .B(G113), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G15));
  NAND3_X1  g497(.A1(new_n680), .A2(new_n587), .A3(new_n629), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G116), .ZN(G18));
  NAND2_X1  g499(.A1(new_n585), .A2(new_n586), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n470), .A2(new_n675), .A3(new_n192), .A4(new_n296), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n406), .A2(new_n480), .A3(new_n640), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n686), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G119), .ZN(G21));
  NAND2_X1  g505(.A1(new_n561), .A2(new_n564), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT101), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n552), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n561), .A2(new_n564), .A3(KEYINPUT101), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n579), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n576), .ZN(new_n698));
  INV_X1    g512(.A(new_n520), .ZN(new_n699));
  AND3_X1   g513(.A1(new_n698), .A2(new_n699), .A3(new_n614), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n597), .A2(new_n665), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n680), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G122), .ZN(G24));
  INV_X1    g517(.A(KEYINPUT102), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n698), .A2(new_n704), .A3(new_n614), .A4(new_n640), .ZN(new_n705));
  AOI22_X1  g519(.A1(new_n694), .A2(new_n695), .B1(new_n572), .B2(new_n573), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n614), .B(new_n640), .C1(new_n706), .C2(new_n577), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT102), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n687), .A2(new_n670), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(KEYINPUT103), .B(G125), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G27));
  NOR2_X1   g527(.A1(new_n596), .A2(new_n408), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n306), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n587), .A2(new_n671), .A3(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT42), .ZN(new_n718));
  NOR4_X1   g532(.A1(new_n306), .A2(new_n715), .A3(new_n718), .A4(new_n670), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n568), .A2(new_n578), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n720), .B1(KEYINPUT104), .B2(new_n582), .ZN(new_n721));
  OR2_X1    g535(.A1(new_n582), .A2(KEYINPUT104), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n520), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n717), .A2(new_n718), .B1(new_n719), .B2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n337), .ZN(G33));
  INV_X1    g539(.A(KEYINPUT105), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n647), .B(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n587), .A2(new_n716), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(KEYINPUT106), .B(G134), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(G36));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n731), .B1(new_n303), .B2(new_n304), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n313), .A2(KEYINPUT45), .A3(new_n314), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n732), .A2(new_n733), .A3(G469), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n297), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT46), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n734), .A2(KEYINPUT46), .A3(new_n297), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n296), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n192), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n368), .A2(new_n607), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT107), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(KEYINPUT43), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n746), .B1(new_n742), .B2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(new_n615), .A3(new_n640), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n750));
  OR2_X1    g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n715), .B1(new_n749), .B2(new_n750), .ZN(new_n752));
  AND4_X1   g566(.A1(new_n651), .A2(new_n741), .A3(new_n751), .A4(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n262), .ZN(G39));
  INV_X1    g568(.A(new_n686), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n715), .A2(new_n699), .A3(new_n670), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n741), .A2(KEYINPUT47), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT47), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n740), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n757), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  XOR2_X1   g575(.A(new_n761), .B(G140), .Z(G42));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n666), .A2(new_n470), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n764), .A2(new_n306), .A3(new_n645), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n664), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n649), .A2(new_n672), .A3(new_n711), .A4(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n592), .A2(new_n593), .A3(new_n647), .ZN(new_n770));
  AOI22_X1  g584(.A1(new_n770), .A2(new_n642), .B1(new_n709), .B2(new_n710), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n771), .A2(KEYINPUT52), .A3(new_n672), .A4(new_n766), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n681), .A2(new_n684), .A3(new_n702), .A4(new_n690), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n306), .A2(new_n715), .A3(new_n670), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n709), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n405), .A2(new_n645), .ZN(new_n777));
  AND4_X1   g591(.A1(new_n627), .A2(new_n714), .A3(new_n640), .A4(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n778), .A2(new_n686), .A3(new_n307), .A4(new_n318), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n776), .A2(new_n728), .A3(new_n779), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n774), .A2(new_n724), .A3(new_n780), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n773), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n597), .A2(new_n609), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n594), .A2(new_n783), .A3(new_n616), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n590), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(KEYINPUT108), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT108), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n590), .A2(new_n787), .A3(new_n784), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n364), .A2(new_n405), .A3(new_n367), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n597), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT109), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(new_n594), .A3(new_n616), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n637), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n786), .A2(new_n788), .A3(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n782), .A2(new_n797), .A3(KEYINPUT53), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n771), .A2(new_n768), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n782), .A2(new_n797), .A3(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n763), .A2(new_n798), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n794), .B1(KEYINPUT108), .B2(new_n785), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n804), .A2(new_n773), .A3(new_n788), .A4(new_n781), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n763), .B(new_n802), .C1(new_n805), .C2(new_n799), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(KEYINPUT54), .B1(new_n803), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n782), .A2(new_n797), .A3(KEYINPUT53), .A4(new_n800), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n773), .A2(new_n781), .ZN(new_n811));
  OAI211_X1 g625(.A(KEYINPUT111), .B(new_n802), .C1(new_n811), .C2(new_n796), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT111), .B1(new_n805), .B2(new_n802), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n809), .B(new_n810), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n808), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n748), .A2(new_n473), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT112), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n748), .A2(KEYINPUT112), .A3(new_n473), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n821), .A2(new_n700), .A3(new_n714), .ZN(new_n822));
  XOR2_X1   g636(.A(new_n822), .B(KEYINPUT113), .Z(new_n823));
  AND2_X1   g637(.A1(new_n675), .A2(new_n296), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n192), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n826), .B1(new_n825), .B2(new_n824), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n758), .A2(new_n760), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n823), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n676), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n656), .A2(new_n408), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n821), .A2(new_n700), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT50), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n830), .A2(new_n714), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT115), .ZN(new_n837));
  AND4_X1   g651(.A1(new_n699), .A2(new_n837), .A3(new_n473), .A4(new_n663), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n608), .A2(new_n368), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n821), .A2(new_n837), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n838), .A2(new_n839), .B1(new_n840), .B2(new_n709), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n829), .A2(KEYINPUT51), .A3(new_n835), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n840), .A2(new_n723), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n843), .B(KEYINPUT48), .Z(new_n844));
  AOI21_X1  g658(.A(new_n472), .B1(new_n838), .B2(new_n611), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n821), .A2(new_n688), .A3(new_n700), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n845), .A2(KEYINPUT117), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT117), .B1(new_n845), .B2(new_n846), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n844), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n835), .A2(new_n841), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n850), .A2(KEYINPUT116), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(KEYINPUT116), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n851), .A2(new_n829), .A3(new_n852), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n842), .B(new_n849), .C1(new_n853), .C2(KEYINPUT51), .ZN(new_n854));
  OAI22_X1  g668(.A1(new_n816), .A2(new_n854), .B1(G952), .B2(G953), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n699), .A2(new_n742), .A3(new_n192), .A4(new_n407), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n657), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT49), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n824), .A2(new_n858), .ZN(new_n859));
  OR2_X1    g673(.A1(new_n824), .A2(new_n858), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n857), .A2(new_n663), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n855), .A2(new_n861), .ZN(G75));
  OAI21_X1  g676(.A(new_n810), .B1(new_n813), .B2(new_n814), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n863), .A2(G210), .A3(G902), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT56), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n439), .A2(new_n445), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n866), .A2(new_n465), .ZN(new_n867));
  XNOR2_X1  g681(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n867), .B(new_n868), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n864), .A2(new_n865), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n869), .B1(new_n864), .B2(new_n865), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n195), .A2(G952), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(G51));
  XOR2_X1   g687(.A(new_n297), .B(KEYINPUT57), .Z(new_n874));
  INV_X1    g688(.A(new_n815), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n802), .B1(new_n811), .B2(new_n796), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT111), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(new_n812), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n809), .B1(new_n879), .B2(new_n810), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n874), .B1(new_n875), .B2(new_n880), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n292), .A2(new_n295), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n805), .A2(new_n799), .ZN(new_n884));
  AOI22_X1  g698(.A1(new_n878), .A2(new_n812), .B1(new_n884), .B2(KEYINPUT53), .ZN(new_n885));
  OR3_X1    g699(.A1(new_n885), .A2(new_n190), .A3(new_n734), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n872), .B1(new_n883), .B2(new_n886), .ZN(G54));
  NAND2_X1  g701(.A1(KEYINPUT58), .A2(G475), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT119), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n863), .A2(G902), .A3(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n360), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n890), .A2(KEYINPUT120), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n872), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n893), .B1(new_n890), .B2(new_n891), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT120), .B1(new_n890), .B2(new_n891), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n892), .A2(new_n894), .A3(new_n895), .ZN(G60));
  NAND2_X1  g710(.A1(G478), .A2(G902), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT59), .Z(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n605), .B1(new_n816), .B2(new_n899), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n605), .A2(new_n899), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n901), .B1(new_n875), .B2(new_n880), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n893), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n900), .A2(new_n903), .ZN(G63));
  NAND2_X1  g718(.A1(G217), .A2(G902), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT121), .Z(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT60), .Z(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n519), .B1(new_n885), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n863), .A2(new_n634), .A3(new_n907), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n909), .A2(new_n893), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT61), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n909), .A2(KEYINPUT61), .A3(new_n910), .A4(new_n893), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(G66));
  AOI21_X1  g729(.A(new_n195), .B1(new_n478), .B2(G224), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n796), .A2(new_n774), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n916), .B1(new_n917), .B2(new_n195), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n435), .B(new_n438), .C1(G898), .C2(new_n195), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n918), .B(new_n919), .Z(G69));
  INV_X1    g734(.A(KEYINPUT123), .ZN(new_n921));
  INV_X1    g735(.A(new_n728), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n771), .A2(new_n672), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n753), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AOI211_X1 g738(.A(new_n520), .B(new_n764), .C1(new_n721), .C2(new_n722), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n741), .A2(new_n651), .A3(new_n925), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT124), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n761), .A2(new_n724), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n924), .A2(new_n927), .A3(new_n928), .A4(new_n195), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n528), .A2(new_n533), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(new_n350), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(G900), .B2(G953), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n921), .B1(new_n929), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT125), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n195), .B1(G227), .B2(G900), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n935), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(KEYINPUT125), .B1(new_n934), .B2(new_n937), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n929), .A2(new_n933), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n715), .B1(new_n609), .B2(new_n789), .ZN(new_n943));
  AND4_X1   g757(.A1(new_n587), .A2(new_n594), .A3(new_n651), .A4(new_n943), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n761), .A2(new_n753), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n668), .A2(new_n672), .A3(new_n771), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(KEYINPUT62), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT62), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n668), .A2(new_n948), .A3(new_n672), .A4(new_n771), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n945), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(KEYINPUT122), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT122), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n945), .A2(new_n947), .A3(new_n952), .A4(new_n949), .ZN(new_n953));
  AOI21_X1  g767(.A(G953), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n942), .B1(new_n954), .B2(new_n931), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n941), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n941), .A2(new_n955), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n956), .A2(new_n957), .ZN(G72));
  NAND2_X1  g772(.A1(G472), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT63), .Z(new_n960));
  NAND2_X1  g774(.A1(new_n951), .A2(new_n953), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n960), .B1(new_n961), .B2(new_n917), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n537), .B(KEYINPUT126), .Z(new_n963));
  AND2_X1   g777(.A1(new_n963), .A2(new_n552), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n924), .A2(new_n927), .A3(new_n928), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n960), .B1(new_n966), .B2(new_n917), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n963), .A2(new_n552), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n872), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n965), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n537), .A2(new_n542), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n570), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n960), .B(new_n972), .C1(new_n803), .C2(new_n807), .ZN(new_n973));
  OR2_X1    g787(.A1(new_n973), .A2(KEYINPUT127), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(KEYINPUT127), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n970), .B1(new_n974), .B2(new_n975), .ZN(G57));
endmodule


