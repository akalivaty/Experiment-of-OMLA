//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1 1 0 0 1 1 1 1 1 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n579,
    new_n580, new_n581, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n631, new_n634, new_n636, new_n637, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT65), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OR2_X1    g036(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G137), .ZN(new_n470));
  NAND2_X1  g045(.A1(G101), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  OAI21_X1  g049(.A(G125), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n475), .A2(new_n476), .B1(G113), .B2(G2104), .ZN(new_n477));
  OAI211_X1 g052(.A(KEYINPUT66), .B(G125), .C1(new_n473), .C2(new_n474), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n472), .B1(new_n479), .B2(G2105), .ZN(G160));
  INV_X1    g055(.A(G2105), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n481), .B1(new_n467), .B2(new_n468), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(new_n481), .B2(G112), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n473), .A2(new_n474), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT67), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT67), .B1(new_n487), .B2(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n486), .B1(new_n492), .B2(G136), .ZN(G162));
  OAI21_X1  g068(.A(G2104), .B1(new_n481), .B2(G114), .ZN(new_n494));
  NOR2_X1   g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT68), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT68), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n497), .A2(new_n499), .A3(new_n500), .A4(G2104), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n482), .A2(G126), .ZN(new_n503));
  OAI211_X1 g078(.A(G138), .B(new_n481), .C1(new_n473), .C2(new_n474), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n469), .A2(KEYINPUT4), .A3(G138), .A4(new_n481), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n502), .A2(new_n503), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  NAND2_X1  g084(.A1(G75), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT69), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n512), .B2(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(KEYINPUT69), .A3(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G62), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n510), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G651), .ZN(new_n521));
  INV_X1    g096(.A(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT6), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT6), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G651), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT70), .B(G88), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n526), .A2(new_n516), .A3(new_n517), .A4(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT71), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n526), .A2(G50), .A3(G543), .ZN(new_n530));
  AND3_X1   g105(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n529), .B1(new_n528), .B2(new_n530), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n521), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT72), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT72), .ZN(new_n535));
  OAI211_X1 g110(.A(new_n521), .B(new_n535), .C1(new_n531), .C2(new_n532), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(new_n536), .ZN(G166));
  AND2_X1   g112(.A1(new_n526), .A2(G543), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n516), .A2(new_n517), .ZN(new_n539));
  AND2_X1   g114(.A1(G63), .A2(G651), .ZN(new_n540));
  AOI22_X1  g115(.A1(G51), .A2(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT73), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT7), .ZN(new_n544));
  INV_X1    g119(.A(G89), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n539), .A2(new_n526), .ZN(new_n546));
  OAI211_X1 g121(.A(new_n541), .B(new_n544), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT74), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AND2_X1   g124(.A1(new_n539), .A2(new_n526), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G89), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n551), .A2(KEYINPUT74), .A3(new_n544), .A4(new_n541), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(G168));
  NAND2_X1  g128(.A1(G77), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G64), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n518), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G651), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n557), .A2(KEYINPUT75), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(KEYINPUT75), .ZN(new_n559));
  XNOR2_X1  g134(.A(KEYINPUT76), .B(G90), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n550), .A2(new_n560), .B1(G52), .B2(new_n538), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n558), .A2(new_n559), .A3(new_n561), .ZN(G301));
  INV_X1    g137(.A(G301), .ZN(G171));
  NAND2_X1  g138(.A1(new_n538), .A2(G43), .ZN(new_n564));
  INV_X1    g139(.A(G81), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n546), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(G68), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G56), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n518), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G651), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n567), .A2(KEYINPUT77), .A3(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n573));
  INV_X1    g148(.A(new_n571), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n574), .B2(new_n566), .ZN(new_n575));
  AND2_X1   g150(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G860), .ZN(G153));
  NAND4_X1  g152(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g153(.A1(G1), .A2(G3), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT8), .ZN(new_n580));
  NAND4_X1  g155(.A1(G319), .A2(G483), .A3(G661), .A4(new_n580), .ZN(new_n581));
  XOR2_X1   g156(.A(new_n581), .B(KEYINPUT78), .Z(G188));
  NAND3_X1  g157(.A1(new_n516), .A2(G65), .A3(new_n517), .ZN(new_n583));
  NAND2_X1  g158(.A1(G78), .A2(G543), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT79), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G651), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n539), .A2(G91), .A3(new_n526), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n523), .A2(new_n525), .A3(G53), .A4(G543), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT9), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n587), .A2(new_n588), .A3(new_n590), .ZN(G299));
  INV_X1    g166(.A(G168), .ZN(G286));
  INV_X1    g167(.A(G166), .ZN(G303));
  OAI21_X1  g168(.A(G651), .B1(new_n539), .B2(G74), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n538), .A2(G49), .ZN(new_n595));
  INV_X1    g170(.A(G87), .ZN(new_n596));
  OAI211_X1 g171(.A(new_n594), .B(new_n595), .C1(new_n596), .C2(new_n546), .ZN(G288));
  NAND2_X1  g172(.A1(G73), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G61), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n518), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G651), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n538), .A2(G48), .ZN(new_n603));
  INV_X1    g178(.A(G86), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n546), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(G305));
  AOI22_X1  g182(.A1(new_n539), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(new_n522), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n538), .A2(G47), .ZN(new_n610));
  INV_X1    g185(.A(G85), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n546), .B2(new_n611), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n609), .A2(new_n612), .ZN(G290));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  NOR2_X1   g189(.A1(G301), .A2(new_n614), .ZN(new_n615));
  AND2_X1   g190(.A1(G79), .A2(G543), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(new_n539), .B2(G66), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT80), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n617), .A2(new_n618), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n619), .A2(G651), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n550), .A2(KEYINPUT10), .A3(G92), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT10), .ZN(new_n623));
  INV_X1    g198(.A(G92), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n546), .B2(new_n624), .ZN(new_n625));
  AOI22_X1  g200(.A1(new_n622), .A2(new_n625), .B1(G54), .B2(new_n538), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT81), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n615), .B1(new_n628), .B2(new_n614), .ZN(G321));
  XOR2_X1   g204(.A(G321), .B(KEYINPUT82), .Z(G284));
  NOR2_X1   g205(.A1(G299), .A2(G868), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n631), .B1(G168), .B2(G868), .ZN(G297));
  XOR2_X1   g207(.A(G297), .B(KEYINPUT83), .Z(G280));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n628), .B1(new_n634), .B2(G860), .ZN(G148));
  NAND3_X1  g210(.A1(new_n628), .A2(new_n634), .A3(G868), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n576), .A2(new_n614), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT11), .Z(G282));
  INV_X1    g214(.A(new_n638), .ZN(G323));
  NAND2_X1  g215(.A1(new_n488), .A2(G2104), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT84), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT13), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT85), .B(G2100), .Z(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n482), .A2(G123), .ZN(new_n648));
  NOR2_X1   g223(.A1(G99), .A2(G2105), .ZN(new_n649));
  OAI21_X1  g224(.A(G2104), .B1(new_n481), .B2(G111), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(new_n492), .B2(G135), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2096), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n646), .A2(new_n647), .A3(new_n653), .ZN(G156));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n655), .B(new_n656), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT15), .B(G2435), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2438), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2427), .B(G2430), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(KEYINPUT14), .ZN(new_n663));
  AND2_X1   g238(.A1(new_n663), .A2(KEYINPUT87), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(KEYINPUT87), .ZN(new_n665));
  OAI22_X1  g240(.A1(new_n664), .A2(new_n665), .B1(new_n660), .B2(new_n661), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1341), .B(G1348), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n667), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n666), .B(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n673), .A2(new_n669), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n658), .B1(new_n671), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n669), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n668), .A2(new_n670), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n676), .A2(new_n677), .A3(new_n657), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n675), .A2(G14), .A3(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT88), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g256(.A1(new_n675), .A2(KEYINPUT88), .A3(G14), .A4(new_n678), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(G401));
  XOR2_X1   g259(.A(G2084), .B(G2090), .Z(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G2072), .B(G2078), .Z(new_n687));
  XNOR2_X1  g262(.A(G2067), .B(G2678), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NOR3_X1   g264(.A1(new_n686), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT18), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n688), .B1(new_n687), .B2(KEYINPUT89), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(KEYINPUT89), .B2(new_n687), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n687), .B(KEYINPUT17), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n693), .B(new_n686), .C1(new_n694), .C2(new_n689), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n694), .A2(new_n689), .A3(new_n685), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n691), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(G2096), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G2100), .ZN(G227));
  XOR2_X1   g274(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n700));
  XNOR2_X1  g275(.A(G1956), .B(G2474), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1961), .B(G1966), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(new_n703), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1971), .B(G1976), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT90), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT19), .ZN(new_n710));
  MUX2_X1   g285(.A(new_n703), .B(new_n706), .S(new_n710), .Z(new_n711));
  OR3_X1    g286(.A1(new_n710), .A2(KEYINPUT20), .A3(new_n705), .ZN(new_n712));
  OAI21_X1  g287(.A(KEYINPUT20), .B1(new_n710), .B2(new_n705), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT91), .B(G1986), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n711), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n715), .B1(new_n711), .B2(new_n714), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n700), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n711), .A2(new_n714), .ZN(new_n720));
  INV_X1    g295(.A(new_n715), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n700), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n722), .A2(new_n723), .A3(new_n716), .ZN(new_n724));
  XNOR2_X1  g299(.A(G1991), .B(G1996), .ZN(new_n725));
  INV_X1    g300(.A(G1981), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  AND3_X1   g302(.A1(new_n719), .A2(new_n724), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n727), .B1(new_n719), .B2(new_n724), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(G229));
  INV_X1    g306(.A(G16), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G24), .ZN(new_n733));
  INV_X1    g308(.A(G290), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n734), .A2(KEYINPUT94), .ZN(new_n735));
  OAI21_X1  g310(.A(G16), .B1(new_n734), .B2(KEYINPUT94), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n733), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n737), .A2(G1986), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n737), .A2(G1986), .ZN(new_n739));
  INV_X1    g314(.A(G29), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G25), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT92), .ZN(new_n742));
  OR2_X1    g317(.A1(G95), .A2(G2105), .ZN(new_n743));
  INV_X1    g318(.A(G107), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n466), .B1(new_n744), .B2(G2105), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n482), .A2(G119), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n492), .B2(G131), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT93), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n742), .B1(new_n749), .B2(new_n740), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT35), .B(G1991), .Z(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n739), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(G6), .A2(G16), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n606), .B2(G16), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT32), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G1981), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT95), .ZN(new_n758));
  NAND2_X1  g333(.A1(G288), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n550), .A2(G87), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n760), .A2(KEYINPUT95), .A3(new_n594), .A4(new_n595), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  MUX2_X1   g337(.A(G23), .B(new_n762), .S(G16), .Z(new_n763));
  XOR2_X1   g338(.A(KEYINPUT33), .B(G1976), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n757), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(G16), .A2(G22), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G166), .B2(G16), .ZN(new_n768));
  INV_X1    g343(.A(G1971), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n770), .A2(KEYINPUT96), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(KEYINPUT96), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n766), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  AOI211_X1 g348(.A(new_n738), .B(new_n753), .C1(new_n773), .C2(KEYINPUT34), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n773), .A2(KEYINPUT34), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n776), .A2(KEYINPUT36), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT36), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n774), .A2(new_n778), .A3(new_n775), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n732), .A2(G21), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G168), .B2(new_n732), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n782), .A2(G1966), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT100), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(G1966), .ZN(new_n785));
  INV_X1    g360(.A(G28), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n786), .A2(KEYINPUT30), .ZN(new_n787));
  AOI21_X1  g362(.A(G29), .B1(new_n786), .B2(KEYINPUT30), .ZN(new_n788));
  OR2_X1    g363(.A1(KEYINPUT31), .A2(G11), .ZN(new_n789));
  NAND2_X1  g364(.A1(KEYINPUT31), .A2(G11), .ZN(new_n790));
  AOI22_X1  g365(.A1(new_n787), .A2(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n652), .A2(G29), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(KEYINPUT99), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n732), .A2(G5), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G301), .B2(G16), .ZN(new_n795));
  INV_X1    g370(.A(G1961), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI211_X1 g372(.A(new_n793), .B(new_n797), .C1(KEYINPUT99), .C2(new_n792), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n784), .A2(new_n785), .A3(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT101), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n740), .A2(G27), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G164), .B2(new_n740), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(new_n443), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n740), .A2(G32), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n482), .A2(G129), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT98), .Z(new_n808));
  NAND3_X1  g383(.A1(new_n481), .A2(G105), .A3(G2104), .ZN(new_n809));
  NAND3_X1  g384(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT26), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n808), .B(new_n809), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n492), .A2(G141), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n806), .B1(new_n816), .B2(new_n740), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT27), .B(G1996), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT24), .ZN(new_n820));
  INV_X1    g395(.A(G34), .ZN(new_n821));
  AOI21_X1  g396(.A(G29), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n820), .B2(new_n821), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G160), .B2(new_n740), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n819), .B1(G2084), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n740), .A2(G33), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n481), .A2(G103), .A3(G2104), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT25), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n830), .B2(new_n481), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(new_n492), .B2(G139), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n826), .B1(new_n832), .B2(new_n740), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(new_n442), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n824), .A2(G2084), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT102), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(new_n796), .B2(new_n795), .ZN(new_n837));
  AND4_X1   g412(.A1(new_n805), .A2(new_n825), .A3(new_n834), .A4(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n801), .A2(new_n802), .A3(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT103), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n801), .A2(KEYINPUT103), .A3(new_n802), .A4(new_n838), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n732), .A2(G4), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n628), .B2(new_n732), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n844), .A2(G1348), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(G1348), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n732), .A2(G20), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT23), .Z(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(G299), .B2(G16), .ZN(new_n849));
  INV_X1    g424(.A(G1956), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n740), .A2(G35), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(G162), .B2(new_n740), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT29), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n851), .B1(G2090), .B2(new_n854), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n854), .A2(G2090), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n740), .A2(G26), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT28), .Z(new_n858));
  NAND2_X1  g433(.A1(new_n482), .A2(G128), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT97), .Z(new_n860));
  NAND2_X1  g435(.A1(new_n492), .A2(G140), .ZN(new_n861));
  NOR2_X1   g436(.A1(G104), .A2(G2105), .ZN(new_n862));
  OAI21_X1  g437(.A(G2104), .B1(new_n481), .B2(G116), .ZN(new_n863));
  OAI211_X1 g438(.A(new_n860), .B(new_n861), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n858), .B1(new_n864), .B2(G29), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(G2067), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n855), .A2(new_n856), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n732), .A2(G19), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n868), .B1(new_n576), .B2(new_n732), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(G1341), .ZN(new_n870));
  NOR4_X1   g445(.A1(new_n845), .A2(new_n846), .A3(new_n867), .A4(new_n870), .ZN(new_n871));
  AND4_X1   g446(.A1(new_n780), .A2(new_n841), .A3(new_n842), .A4(new_n871), .ZN(G311));
  NAND4_X1  g447(.A1(new_n780), .A2(new_n841), .A3(new_n842), .A4(new_n871), .ZN(G150));
  INV_X1    g448(.A(KEYINPUT107), .ZN(new_n874));
  AOI22_X1  g449(.A1(new_n539), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n875), .A2(new_n522), .ZN(new_n876));
  XNOR2_X1  g451(.A(KEYINPUT105), .B(G93), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n539), .A2(new_n526), .A3(new_n877), .ZN(new_n878));
  XOR2_X1   g453(.A(KEYINPUT104), .B(G55), .Z(new_n879));
  NAND2_X1  g454(.A1(new_n538), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT106), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n878), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n881), .B1(new_n878), .B2(new_n880), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n876), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n884), .A2(new_n572), .A3(new_n575), .ZN(new_n885));
  OAI221_X1 g460(.A(new_n876), .B1(new_n574), .B2(new_n566), .C1(new_n882), .C2(new_n883), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n874), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n885), .A2(new_n874), .A3(new_n886), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT38), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n628), .A2(G559), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n891), .B(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT39), .ZN(new_n894));
  AOI21_X1  g469(.A(G860), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n895), .B1(new_n894), .B2(new_n893), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n884), .A2(G860), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n897), .B(KEYINPUT37), .Z(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(G145));
  XOR2_X1   g474(.A(new_n652), .B(G160), .Z(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(G162), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n482), .A2(G130), .ZN(new_n902));
  NOR2_X1   g477(.A1(G106), .A2(G2105), .ZN(new_n903));
  OAI21_X1  g478(.A(G2104), .B1(new_n481), .B2(G118), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n905), .B1(new_n492), .B2(G142), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n642), .B(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n748), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n907), .A2(new_n908), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT109), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT109), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(new_n909), .B2(new_n910), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n832), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT108), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n508), .A2(new_n917), .ZN(new_n918));
  AOI22_X1  g493(.A1(new_n496), .A2(new_n501), .B1(new_n482), .B2(G126), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n919), .A2(KEYINPUT108), .A3(new_n506), .A4(new_n507), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n864), .B(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n816), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n922), .A2(new_n923), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n916), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n926), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n928), .A2(new_n832), .A3(new_n924), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n915), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n915), .B1(new_n927), .B2(new_n929), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n901), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(G37), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n927), .A2(new_n929), .A3(new_n911), .ZN(new_n934));
  INV_X1    g509(.A(new_n901), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n927), .A2(new_n929), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n934), .B(new_n935), .C1(new_n936), .C2(new_n915), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n932), .A2(new_n933), .A3(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g514(.A(new_n628), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n890), .B1(new_n940), .B2(G559), .ZN(new_n941));
  INV_X1    g516(.A(new_n889), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n942), .A2(new_n887), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n943), .A2(new_n634), .A3(new_n628), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT41), .ZN(new_n945));
  INV_X1    g520(.A(new_n627), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n946), .A2(G299), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n946), .A2(G299), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n945), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n627), .B(G299), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT41), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n941), .A2(new_n944), .A3(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n950), .B1(new_n941), .B2(new_n944), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT42), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT42), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n941), .A2(new_n944), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n957), .B(new_n953), .C1(new_n958), .C2(new_n950), .ZN(new_n959));
  XNOR2_X1  g534(.A(G166), .B(new_n734), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n762), .B(G305), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n960), .B(new_n961), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n956), .A2(new_n959), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n962), .B1(new_n956), .B2(new_n959), .ZN(new_n964));
  OAI21_X1  g539(.A(G868), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n884), .A2(new_n614), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n966), .B1(new_n965), .B2(new_n967), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(G295));
  NAND2_X1  g545(.A1(new_n965), .A2(new_n967), .ZN(G331));
  XNOR2_X1  g546(.A(G168), .B(G301), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n972), .A2(new_n888), .A3(new_n889), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT111), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT111), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n943), .A2(new_n975), .A3(new_n972), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n943), .A2(new_n972), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n952), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OR2_X1    g554(.A1(new_n943), .A2(new_n972), .ZN(new_n980));
  INV_X1    g555(.A(new_n950), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n980), .A2(new_n981), .A3(new_n973), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n962), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n978), .B1(new_n974), .B2(new_n976), .ZN(new_n984));
  INV_X1    g559(.A(new_n952), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n962), .B(new_n982), .C1(new_n984), .C2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n933), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n983), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n988), .A2(KEYINPUT43), .ZN(new_n989));
  INV_X1    g564(.A(new_n962), .ZN(new_n990));
  AOI211_X1 g565(.A(new_n950), .B(new_n978), .C1(new_n974), .C2(new_n976), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n985), .B1(new_n980), .B2(new_n973), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AND4_X1   g568(.A1(KEYINPUT43), .A2(new_n993), .A3(new_n933), .A4(new_n986), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT44), .B1(new_n989), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT43), .B1(new_n983), .B2(new_n987), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT43), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n993), .A2(new_n997), .A3(new_n933), .A4(new_n986), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n995), .B1(KEYINPUT44), .B2(new_n1000), .ZN(G397));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1002), .B1(new_n921), .B2(G1384), .ZN(new_n1003));
  NAND2_X1  g578(.A1(G113), .A2(G2104), .ZN(new_n1004));
  INV_X1    g579(.A(G125), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1005), .B1(new_n467), .B2(new_n468), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1004), .B1(new_n1006), .B2(KEYINPUT66), .ZN(new_n1007));
  INV_X1    g582(.A(new_n478), .ZN(new_n1008));
  OAI21_X1  g583(.A(G2105), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n472), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(G40), .A3(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1003), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n749), .A2(new_n751), .ZN(new_n1013));
  XOR2_X1   g588(.A(new_n864), .B(G2067), .Z(new_n1014));
  NAND2_X1  g589(.A1(new_n923), .A2(G1996), .ZN(new_n1015));
  INV_X1    g590(.A(G1996), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n816), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1014), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1013), .B1(new_n1018), .B2(new_n1012), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n864), .A2(G2067), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1012), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n748), .B(new_n751), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1012), .B1(new_n1018), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(G290), .A2(G1986), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1012), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1023), .B1(KEYINPUT48), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT48), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1012), .A2(new_n1016), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT46), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n1032), .B(KEYINPUT126), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1014), .A2(new_n816), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n1034), .A2(new_n1012), .B1(new_n1031), .B2(new_n1030), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT47), .ZN(new_n1037));
  OAI221_X1 g612(.A(new_n1021), .B1(new_n1027), .B2(new_n1029), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1038), .B1(new_n1037), .B2(new_n1036), .ZN(new_n1039));
  INV_X1    g614(.A(G1384), .ZN(new_n1040));
  NAND4_X1  g615(.A1(G160), .A2(G40), .A3(new_n1040), .A4(new_n508), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1041), .A2(G8), .ZN(new_n1042));
  INV_X1    g617(.A(G1976), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT52), .B1(G288), .B2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1042), .B(new_n1044), .C1(new_n762), .C2(new_n1043), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1042), .B1(new_n762), .B2(new_n1043), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT52), .ZN(new_n1047));
  OAI21_X1  g622(.A(G1981), .B1(new_n602), .B2(new_n605), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n602), .A2(new_n605), .A3(G1981), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT117), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1042), .B1(new_n1051), .B2(KEYINPUT49), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT49), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n606), .A2(new_n726), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n1048), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1053), .B1(new_n1055), .B2(KEYINPUT117), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1045), .B(new_n1047), .C1(new_n1052), .C2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1058), .A2(KEYINPUT114), .ZN(new_n1059));
  INV_X1    g634(.A(G8), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1060), .B1(KEYINPUT114), .B2(new_n1058), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1059), .B1(G166), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1059), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n534), .A2(new_n536), .A3(new_n1064), .A4(new_n1061), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n508), .A2(new_n1040), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1011), .B1(new_n1002), .B2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n918), .A2(KEYINPUT45), .A3(new_n920), .A4(new_n1040), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n769), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT50), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n508), .A2(new_n1072), .A3(new_n1040), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1067), .A2(KEYINPUT50), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1009), .A2(G40), .A3(new_n1010), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n508), .A2(KEYINPUT118), .A3(new_n1072), .A4(new_n1040), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1071), .B1(G2090), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(G8), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1057), .B1(new_n1066), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT116), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT113), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1073), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n1076), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1072), .B1(new_n508), .B2(new_n1040), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1011), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(G2090), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1086), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1071), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(G8), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT115), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1093), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1063), .A2(new_n1093), .A3(new_n1065), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1083), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1066), .A2(KEYINPUT115), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1060), .B1(new_n1071), .B2(new_n1090), .ZN(new_n1099));
  AND4_X1   g674(.A1(new_n1083), .A2(new_n1098), .A3(new_n1096), .A4(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1082), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n796), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n508), .A2(KEYINPUT45), .A3(new_n1040), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1105), .A2(G2078), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1068), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1067), .A2(new_n1002), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1069), .A2(new_n443), .A3(new_n1108), .A4(new_n1077), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(new_n1105), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1103), .A2(new_n1107), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1108), .A2(new_n1077), .A3(new_n1104), .ZN(new_n1112));
  INV_X1    g687(.A(G1966), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1114), .B(G168), .C1(new_n1102), .C2(G2084), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1115), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1114), .B1(new_n1102), .B2(G2084), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(G286), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT51), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1115), .A2(G8), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1116), .A2(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(G171), .B(new_n1111), .C1(new_n1121), .C2(KEYINPUT62), .ZN(new_n1122));
  OAI21_X1  g697(.A(KEYINPUT124), .B1(new_n1101), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(KEYINPUT62), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1098), .A2(new_n1096), .A3(new_n1099), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT116), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1095), .A2(new_n1083), .A3(new_n1096), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1111), .A2(G171), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1118), .A2(KEYINPUT51), .A3(G8), .A4(new_n1115), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1120), .A2(new_n1119), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1129), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1128), .A2(new_n1134), .A3(new_n1135), .A4(new_n1082), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1123), .A2(new_n1124), .A3(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1052), .A2(new_n1056), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1138), .A2(G1976), .A3(G288), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1042), .B1(new_n1139), .B2(new_n1050), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(new_n1128), .B2(new_n1057), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1117), .A2(G8), .A3(G168), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1099), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT63), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n1144), .A2(new_n1057), .A3(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1128), .A2(new_n1143), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1141), .B1(KEYINPUT63), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1142), .B1(new_n1128), .B2(new_n1146), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT123), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1103), .A2(G301), .A3(new_n1110), .A4(new_n1107), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(KEYINPUT54), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1069), .A2(new_n1077), .A3(new_n1106), .ZN(new_n1153));
  AOI22_X1  g728(.A1(new_n1153), .A2(new_n1003), .B1(new_n1109), .B2(new_n1105), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT121), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1155), .B1(new_n1102), .B2(new_n796), .ZN(new_n1156));
  AOI211_X1 g731(.A(KEYINPUT121), .B(G1961), .C1(new_n1086), .C2(new_n1088), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1154), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(G301), .B1(new_n1158), .B2(KEYINPUT122), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT122), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1160), .B(new_n1154), .C1(new_n1156), .C2(new_n1157), .ZN(new_n1161));
  AOI211_X1 g736(.A(new_n1150), .B(new_n1152), .C1(new_n1159), .C2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1158), .A2(KEYINPUT122), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1163), .A2(G171), .A3(new_n1161), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1152), .ZN(new_n1165));
  AOI21_X1  g740(.A(KEYINPUT123), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1162), .A2(new_n1166), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1069), .A2(new_n1108), .A3(new_n1077), .ZN(new_n1168));
  XNOR2_X1  g743(.A(KEYINPUT56), .B(G2072), .ZN(new_n1169));
  AOI22_X1  g744(.A1(new_n1168), .A2(new_n1169), .B1(new_n1079), .B2(new_n850), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT119), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT57), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(G299), .A2(new_n1174), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n587), .A2(new_n588), .A3(new_n590), .A4(new_n1173), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(KEYINPUT120), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT120), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1175), .A2(new_n1180), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1170), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1079), .A2(new_n850), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1068), .A2(new_n1069), .A3(new_n1169), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1184), .A2(new_n1185), .A3(new_n1178), .ZN(new_n1186));
  INV_X1    g761(.A(G1348), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1102), .A2(new_n1187), .ZN(new_n1188));
  OR2_X1    g763(.A1(new_n1041), .A2(G2067), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n627), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1183), .B1(new_n1186), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n1192));
  AND3_X1   g767(.A1(new_n1184), .A2(new_n1185), .A3(new_n1178), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1178), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1192), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n1069), .A2(new_n1016), .A3(new_n1108), .A4(new_n1077), .ZN(new_n1196));
  XOR2_X1   g771(.A(KEYINPUT58), .B(G1341), .Z(new_n1197));
  NAND2_X1  g772(.A1(new_n1041), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(new_n576), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT59), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1199), .A2(new_n1202), .A3(new_n576), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1204));
  OAI211_X1 g779(.A(KEYINPUT61), .B(new_n1186), .C1(new_n1170), .C2(new_n1182), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1195), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  AOI21_X1  g781(.A(KEYINPUT60), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1188), .A2(KEYINPUT60), .A3(new_n1189), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1208), .A2(new_n946), .ZN(new_n1209));
  NAND4_X1  g784(.A1(new_n1188), .A2(KEYINPUT60), .A3(new_n627), .A4(new_n1189), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1207), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1191), .B1(new_n1206), .B2(new_n1211), .ZN(new_n1212));
  OAI211_X1 g787(.A(G301), .B(new_n1154), .C1(new_n1156), .C2(new_n1157), .ZN(new_n1213));
  AOI21_X1  g788(.A(KEYINPUT54), .B1(new_n1213), .B2(new_n1129), .ZN(new_n1214));
  NOR2_X1   g789(.A1(new_n1132), .A2(new_n1214), .ZN(new_n1215));
  AND2_X1   g790(.A1(new_n1212), .A2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1149), .B1(new_n1167), .B2(new_n1216), .ZN(new_n1217));
  OAI211_X1 g792(.A(new_n1137), .B(new_n1148), .C1(new_n1217), .C2(new_n1101), .ZN(new_n1218));
  AND2_X1   g793(.A1(G290), .A2(G1986), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1012), .B1(new_n1219), .B2(new_n1024), .ZN(new_n1220));
  XNOR2_X1  g795(.A(new_n1220), .B(KEYINPUT112), .ZN(new_n1221));
  AND2_X1   g796(.A1(new_n1023), .A2(new_n1221), .ZN(new_n1222));
  AND3_X1   g797(.A1(new_n1218), .A2(KEYINPUT125), .A3(new_n1222), .ZN(new_n1223));
  AOI21_X1  g798(.A(KEYINPUT125), .B1(new_n1218), .B2(new_n1222), .ZN(new_n1224));
  OAI21_X1  g799(.A(new_n1039), .B1(new_n1223), .B2(new_n1224), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g800(.A(KEYINPUT127), .ZN(new_n1227));
  NOR2_X1   g801(.A1(G227), .A2(new_n463), .ZN(new_n1228));
  OAI21_X1  g802(.A(new_n1228), .B1(new_n728), .B2(new_n729), .ZN(new_n1229));
  AOI21_X1  g803(.A(new_n1229), .B1(new_n681), .B2(new_n682), .ZN(new_n1230));
  NAND2_X1  g804(.A1(new_n938), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g805(.A(new_n1231), .ZN(new_n1232));
  AOI21_X1  g806(.A(new_n1227), .B1(new_n999), .B2(new_n1232), .ZN(new_n1233));
  AOI211_X1 g807(.A(KEYINPUT127), .B(new_n1231), .C1(new_n996), .C2(new_n998), .ZN(new_n1234));
  NOR2_X1   g808(.A1(new_n1233), .A2(new_n1234), .ZN(G308));
  NAND2_X1  g809(.A1(new_n999), .A2(new_n1232), .ZN(G225));
endmodule


