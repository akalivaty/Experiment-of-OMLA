//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 1 1 0 0 0 1 0 1 1 0 0 1 0 0 1 1 0 1 1 0 1 0 0 0 1 1 1 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 0 1 1 0 0 1 0 0 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1265, new_n1266, new_n1267,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1334, new_n1335;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0006(.A(new_n201), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G50), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(KEYINPUT65), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G20), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n214), .B1(new_n215), .B2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(G13), .ZN(new_n217));
  NAND4_X1  g0017(.A1(new_n217), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(G250), .B1(G257), .B2(G264), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n213), .B1(new_n222), .B2(KEYINPUT0), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT0), .B2(new_n222), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT66), .ZN(new_n225));
  XOR2_X1   g0025(.A(KEYINPUT67), .B(G68), .Z(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G238), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n228), .A2(new_n229), .A3(KEYINPUT68), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G77), .A2(G244), .ZN(new_n231));
  AOI22_X1  g0031(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n232));
  NAND4_X1  g0032(.A1(new_n227), .A2(new_n230), .A3(new_n231), .A4(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(KEYINPUT68), .B1(new_n228), .B2(new_n229), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n215), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT1), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n225), .A2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT2), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G226), .ZN(new_n240));
  INV_X1    g0040(.A(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT69), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G68), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G87), .B(G97), .Z(new_n251));
  XOR2_X1   g0051(.A(G107), .B(G116), .Z(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  AND2_X1   g0055(.A1(new_n255), .A2(new_n210), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(KEYINPUT70), .A2(G1), .ZN(new_n258));
  NOR2_X1   g0058(.A1(KEYINPUT70), .A2(G1), .ZN(new_n259));
  NOR3_X1   g0059(.A1(new_n258), .A2(new_n259), .A3(new_n211), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G50), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT70), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(KEYINPUT70), .A2(G1), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n265), .A2(G13), .A3(G20), .A4(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n262), .B1(G50), .B2(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT8), .B(G58), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT72), .ZN(new_n271));
  INV_X1    g0071(.A(G33), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n271), .B1(new_n272), .B2(G20), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n211), .A2(KEYINPUT72), .A3(G33), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n270), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n256), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n268), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(new_n279), .B(KEYINPUT9), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT3), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n272), .ZN(new_n282));
  NAND2_X1  g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n284), .A2(G223), .A3(G1698), .ZN(new_n285));
  INV_X1    g0085(.A(G77), .ZN(new_n286));
  INV_X1    g0086(.A(G1698), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G222), .ZN(new_n289));
  OAI221_X1 g0089(.A(new_n285), .B1(new_n286), .B2(new_n284), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G41), .A2(G45), .ZN(new_n293));
  INV_X1    g0093(.A(G274), .ZN(new_n294));
  NOR3_X1   g0094(.A1(new_n293), .A2(G1), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G41), .ZN(new_n296));
  OAI211_X1 g0096(.A(G1), .B(G13), .C1(new_n272), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n265), .A2(new_n266), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n297), .B1(new_n298), .B2(new_n293), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n295), .B1(new_n300), .B2(G226), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n292), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT71), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n302), .A2(new_n303), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n280), .B1(new_n307), .B2(G200), .ZN(new_n308));
  OR2_X1    g0108(.A1(new_n305), .A2(new_n306), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G190), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT10), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT10), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n308), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n309), .A2(G179), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n307), .A2(G169), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n279), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT16), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n201), .B1(new_n226), .B2(G58), .ZN(new_n322));
  INV_X1    g0122(.A(G159), .ZN(new_n323));
  INV_X1    g0123(.A(new_n276), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n322), .A2(new_n211), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT67), .B(G68), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT7), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(new_n284), .B2(G20), .ZN(new_n328));
  AND2_X1   g0128(.A1(KEYINPUT3), .A2(G33), .ZN(new_n329));
  NOR2_X1   g0129(.A1(KEYINPUT3), .A2(G33), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n326), .B1(new_n328), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n321), .B1(new_n325), .B2(new_n333), .ZN(new_n334));
  NOR3_X1   g0134(.A1(new_n284), .A2(new_n327), .A3(G20), .ZN(new_n335));
  AOI21_X1  g0135(.A(KEYINPUT7), .B1(new_n331), .B2(new_n211), .ZN(new_n336));
  OAI21_X1  g0136(.A(G68), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G58), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n207), .B1(new_n326), .B2(new_n338), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n339), .A2(G20), .B1(G159), .B2(new_n276), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n337), .A2(new_n340), .A3(KEYINPUT16), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n334), .A2(new_n257), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n267), .A2(new_n269), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(new_n261), .B2(new_n269), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n295), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(new_n299), .B2(new_n241), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n284), .A2(G223), .A3(new_n287), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n284), .A2(G226), .A3(G1698), .ZN(new_n349));
  INV_X1    g0149(.A(G87), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n348), .B(new_n349), .C1(new_n272), .C2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n347), .B1(new_n291), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n352), .A2(G169), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n291), .ZN(new_n354));
  INV_X1    g0154(.A(G179), .ZN(new_n355));
  INV_X1    g0155(.A(new_n347), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n345), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(KEYINPUT18), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT18), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n345), .A2(new_n358), .A3(new_n361), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n284), .A2(G238), .A3(G1698), .ZN(new_n364));
  INV_X1    g0164(.A(G107), .ZN(new_n365));
  OAI221_X1 g0165(.A(new_n364), .B1(new_n365), .B2(new_n284), .C1(new_n288), .C2(new_n241), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n291), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n295), .B1(new_n300), .B2(G244), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G169), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n355), .B2(new_n369), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n273), .A2(new_n274), .ZN(new_n372));
  XNOR2_X1  g0172(.A(KEYINPUT15), .B(G87), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI22_X1  g0174(.A1(new_n269), .A2(new_n324), .B1(new_n211), .B2(new_n286), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n257), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n261), .A2(G77), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n376), .B(new_n377), .C1(G77), .C2(new_n267), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n371), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n369), .ZN(new_n381));
  INV_X1    g0181(.A(G190), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G200), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n369), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n378), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n380), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n354), .A2(new_n356), .A3(new_n382), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(G200), .B2(new_n352), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n389), .A2(new_n342), .A3(new_n344), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT17), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n389), .A2(new_n342), .A3(KEYINPUT17), .A4(new_n344), .ZN(new_n393));
  AND2_X1   g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n363), .A2(new_n387), .A3(new_n394), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n326), .A2(G20), .B1(G50), .B2(new_n276), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n286), .B2(new_n372), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n257), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT11), .ZN(new_n399));
  XNOR2_X1  g0199(.A(new_n398), .B(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT12), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n267), .A2(new_n226), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n402), .B1(new_n401), .B2(new_n267), .ZN(new_n403));
  OAI21_X1  g0203(.A(G68), .B1(new_n261), .B2(new_n401), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n400), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n284), .A2(G232), .A3(G1698), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G97), .ZN(new_n409));
  INV_X1    g0209(.A(G226), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n408), .B(new_n409), .C1(new_n288), .C2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n291), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n295), .B1(new_n300), .B2(G238), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT13), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT13), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n412), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(G179), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(G169), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(new_n415), .B2(new_n417), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT14), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n418), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n417), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n416), .B1(new_n412), .B2(new_n413), .ZN(new_n424));
  OAI21_X1  g0224(.A(G169), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n425), .A2(KEYINPUT14), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n407), .B1(new_n422), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(G200), .B1(new_n415), .B2(new_n417), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n423), .A2(new_n424), .A3(G190), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n406), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  NOR3_X1   g0231(.A1(new_n320), .A2(new_n395), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(G294), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n433), .A2(KEYINPUT83), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n433), .A2(KEYINPUT83), .ZN(new_n435));
  OAI21_X1  g0235(.A(G33), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI211_X1 g0236(.A(G250), .B(new_n287), .C1(new_n329), .C2(new_n330), .ZN(new_n437));
  OAI211_X1 g0237(.A(G257), .B(G1698), .C1(new_n329), .C2(new_n330), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(G45), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n258), .A2(new_n259), .A3(new_n440), .ZN(new_n441));
  XNOR2_X1  g0241(.A(KEYINPUT5), .B(G41), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n291), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n291), .A2(new_n439), .B1(new_n443), .B2(G264), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n441), .A2(G274), .A3(new_n297), .A4(new_n442), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n444), .A2(KEYINPUT84), .A3(new_n382), .A4(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT84), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n439), .A2(new_n291), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n265), .A2(G45), .A3(new_n266), .ZN(new_n449));
  AND2_X1   g0249(.A1(KEYINPUT5), .A2(G41), .ZN(new_n450));
  NOR2_X1   g0250(.A1(KEYINPUT5), .A2(G41), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI211_X1 g0252(.A(G264), .B(new_n297), .C1(new_n449), .C2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n448), .A2(new_n453), .A3(new_n445), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n447), .B1(new_n454), .B2(new_n384), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n454), .A2(G190), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n446), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT81), .ZN(new_n458));
  AND2_X1   g0258(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n459));
  OAI22_X1  g0259(.A1(new_n267), .A2(G107), .B1(KEYINPUT80), .B2(KEYINPUT25), .ZN(new_n460));
  NOR2_X1   g0260(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n260), .A2(G13), .A3(new_n365), .A4(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n459), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n265), .A2(G33), .A3(new_n266), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n267), .A2(new_n256), .A3(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(new_n365), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n458), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n466), .ZN(new_n468));
  AND2_X1   g0268(.A1(new_n460), .A2(new_n462), .ZN(new_n469));
  OAI211_X1 g0269(.A(KEYINPUT81), .B(new_n468), .C1(new_n469), .C2(new_n459), .ZN(new_n470));
  OR3_X1    g0270(.A1(new_n211), .A2(KEYINPUT23), .A3(G107), .ZN(new_n471));
  OAI21_X1  g0271(.A(KEYINPUT23), .B1(new_n211), .B2(G107), .ZN(new_n472));
  AND2_X1   g0272(.A1(KEYINPUT77), .A2(G116), .ZN(new_n473));
  NOR2_X1   g0273(.A1(KEYINPUT77), .A2(G116), .ZN(new_n474));
  OAI21_X1  g0274(.A(G33), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n471), .B(new_n472), .C1(new_n475), .C2(G20), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n211), .B(G87), .C1(new_n329), .C2(new_n330), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT22), .ZN(new_n478));
  AOI21_X1  g0278(.A(G20), .B1(new_n282), .B2(new_n283), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT22), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(new_n480), .A3(G87), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n476), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n256), .B1(new_n482), .B2(KEYINPUT24), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT24), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n481), .A2(new_n478), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n484), .B1(new_n485), .B2(new_n476), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n467), .A2(new_n470), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n457), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n470), .A2(new_n467), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n483), .A2(new_n486), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT82), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n492), .B1(new_n490), .B2(new_n491), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n454), .A2(new_n419), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(G179), .B2(new_n454), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n489), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(G107), .B1(new_n335), .B2(new_n336), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n365), .A2(KEYINPUT6), .A3(G97), .ZN(new_n501));
  INV_X1    g0301(.A(G97), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n502), .A2(new_n365), .ZN(new_n503));
  NOR2_X1   g0303(.A1(G97), .A2(G107), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n501), .B1(new_n505), .B2(KEYINPUT6), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G20), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n276), .A2(G77), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n500), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT73), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n260), .A2(new_n510), .A3(G13), .A4(new_n502), .ZN(new_n511));
  OAI21_X1  g0311(.A(KEYINPUT73), .B1(new_n267), .B2(G97), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n267), .A2(new_n464), .A3(new_n256), .A4(G97), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT74), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT74), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n511), .A2(new_n512), .A3(new_n513), .A4(new_n516), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n257), .A2(new_n509), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(G257), .B(new_n297), .C1(new_n449), .C2(new_n452), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n445), .A2(new_n519), .A3(KEYINPUT76), .ZN(new_n520));
  AOI21_X1  g0320(.A(KEYINPUT76), .B1(new_n445), .B2(new_n519), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT75), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT4), .ZN(new_n524));
  AOI21_X1  g0324(.A(G1698), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n523), .A2(new_n524), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n284), .A2(G244), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G283), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n284), .A2(G250), .A3(G1698), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(G244), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n531), .B1(new_n282), .B2(new_n283), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n526), .B1(new_n532), .B2(new_n525), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n291), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(G200), .B1(new_n522), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n445), .A2(new_n519), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT76), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n445), .A2(new_n519), .A3(KEYINPUT76), .ZN(new_n539));
  AND4_X1   g0339(.A1(new_n382), .A2(new_n534), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n518), .B1(new_n535), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n509), .A2(new_n257), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n515), .A2(new_n517), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n419), .B1(new_n522), .B2(new_n534), .ZN(new_n545));
  AND4_X1   g0345(.A1(G179), .A2(new_n534), .A3(new_n538), .A4(new_n539), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n541), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n267), .A2(new_n464), .A3(new_n256), .A4(G116), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n473), .A2(new_n474), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n260), .A2(G13), .A3(new_n550), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n528), .B1(new_n502), .B2(G33), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n211), .ZN(new_n554));
  OAI21_X1  g0354(.A(G20), .B1(new_n473), .B2(new_n474), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(KEYINPUT20), .B1(new_n556), .B2(new_n257), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT20), .ZN(new_n558));
  AOI211_X1 g0358(.A(new_n558), .B(new_n256), .C1(new_n554), .C2(new_n555), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n552), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(G264), .B(G1698), .C1(new_n329), .C2(new_n330), .ZN(new_n562));
  OAI211_X1 g0362(.A(G257), .B(new_n287), .C1(new_n329), .C2(new_n330), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n282), .A2(G303), .A3(new_n283), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT79), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT79), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n562), .A2(new_n563), .A3(new_n567), .A4(new_n564), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n291), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n291), .B1(new_n441), .B2(new_n294), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n449), .A2(new_n452), .ZN(new_n571));
  AOI22_X1  g0371(.A1(G270), .A2(new_n443), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n569), .A2(new_n572), .A3(new_n382), .ZN(new_n573));
  AOI21_X1  g0373(.A(G200), .B1(new_n569), .B2(new_n572), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n561), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n569), .A2(new_n572), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n576), .A2(G169), .A3(new_n560), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT21), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n576), .A2(KEYINPUT21), .A3(new_n560), .A4(G169), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n569), .A2(new_n572), .A3(G179), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n560), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n575), .A2(new_n579), .A3(new_n580), .A4(new_n582), .ZN(new_n583));
  OAI211_X1 g0383(.A(G244), .B(G1698), .C1(new_n329), .C2(new_n330), .ZN(new_n584));
  OAI211_X1 g0384(.A(G238), .B(new_n287), .C1(new_n329), .C2(new_n330), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n584), .A2(new_n585), .A3(new_n475), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT78), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n584), .A2(new_n585), .A3(KEYINPUT78), .A4(new_n475), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n588), .A2(new_n291), .A3(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n570), .B1(G250), .B2(new_n441), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n590), .A2(new_n355), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n260), .A2(G13), .A3(new_n373), .ZN(new_n593));
  OR2_X1    g0393(.A1(new_n465), .A2(new_n373), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT19), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n211), .B1(new_n409), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n350), .A2(new_n502), .A3(new_n365), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n479), .A2(G68), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n595), .B1(new_n372), .B2(new_n502), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n593), .B(new_n594), .C1(new_n600), .C2(new_n256), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n297), .B1(new_n449), .B2(G274), .ZN(new_n602));
  INV_X1    g0402(.A(G250), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n602), .B1(new_n603), .B2(new_n449), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n589), .A2(new_n291), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n604), .B1(new_n605), .B2(new_n588), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n592), .B(new_n601), .C1(new_n606), .C2(G169), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n586), .A2(new_n587), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n589), .A2(new_n291), .ZN(new_n609));
  OAI211_X1 g0409(.A(G190), .B(new_n591), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n256), .B1(new_n598), .B2(new_n599), .ZN(new_n611));
  INV_X1    g0411(.A(new_n593), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n465), .A2(new_n350), .ZN(new_n613));
  NOR3_X1   g0413(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n610), .B(new_n614), .C1(new_n606), .C2(new_n384), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n607), .A2(new_n615), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n548), .A2(new_n583), .A3(new_n616), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n432), .A2(new_n499), .A3(new_n617), .ZN(G372));
  INV_X1    g0418(.A(new_n427), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n619), .A2(new_n380), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n394), .A2(new_n430), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n363), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n318), .B1(new_n622), .B2(new_n315), .ZN(new_n623));
  INV_X1    g0423(.A(new_n432), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT87), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n490), .A2(new_n491), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT86), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n498), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(KEYINPUT86), .B1(new_n487), .B2(new_n497), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n579), .A2(new_n580), .A3(new_n582), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n625), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n631), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n633), .A2(KEYINPUT87), .A3(new_n628), .A4(new_n629), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n488), .A2(new_n541), .A3(new_n547), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n592), .A2(new_n601), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT85), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n637), .B1(new_n606), .B2(G169), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n590), .A2(new_n591), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n639), .A2(KEYINPUT85), .A3(new_n419), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n636), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n615), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n635), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n632), .A2(new_n634), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n641), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n534), .A2(new_n538), .A3(new_n539), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(G169), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n522), .A2(G179), .A3(new_n534), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n518), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n649), .A2(new_n607), .A3(new_n615), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n645), .B1(new_n650), .B2(KEYINPUT26), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT26), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n641), .A2(new_n649), .A3(new_n652), .A4(new_n615), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n644), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n623), .B1(new_n624), .B2(new_n656), .ZN(G369));
  NAND2_X1  g0457(.A1(new_n626), .A2(KEYINPUT82), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n487), .A2(new_n492), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(new_n659), .A3(new_n498), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n258), .A2(new_n259), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n217), .A2(G20), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G213), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G343), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n660), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n495), .A2(new_n668), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n671), .A2(new_n660), .A3(new_n488), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT88), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(KEYINPUT88), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n670), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n668), .A2(new_n560), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n631), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n677), .B1(new_n583), .B2(new_n676), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G330), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n630), .A2(new_n669), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n633), .A2(new_n668), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n673), .A2(new_n674), .A3(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n681), .A2(new_n682), .A3(new_n684), .ZN(G399));
  NOR2_X1   g0485(.A1(new_n220), .A2(G41), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(new_n264), .ZN(new_n687));
  NOR4_X1   g0487(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n687), .A2(new_n688), .B1(new_n209), .B2(new_n686), .ZN(new_n689));
  XOR2_X1   g0489(.A(new_n689), .B(KEYINPUT28), .Z(new_n690));
  AND3_X1   g0490(.A1(new_n534), .A2(new_n538), .A3(new_n539), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n590), .A2(new_n444), .A3(new_n591), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n581), .A2(new_n691), .A3(new_n692), .A4(KEYINPUT30), .ZN(new_n693));
  AOI21_X1  g0493(.A(G179), .B1(new_n444), .B2(new_n445), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n694), .A2(new_n646), .A3(new_n576), .A4(new_n639), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n590), .A2(new_n444), .A3(new_n591), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n646), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(KEYINPUT30), .B1(new_n698), .B2(new_n581), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n668), .B1(new_n696), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT31), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI211_X1 g0502(.A(KEYINPUT31), .B(new_n668), .C1(new_n696), .C2(new_n699), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(KEYINPUT89), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n617), .A2(new_n499), .A3(new_n669), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(KEYINPUT89), .B1(new_n702), .B2(new_n703), .ZN(new_n707));
  OAI21_X1  g0507(.A(G330), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT91), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n660), .A2(new_n633), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n645), .B1(new_n643), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n652), .B1(new_n547), .B2(new_n616), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT90), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n650), .A2(KEYINPUT90), .A3(new_n652), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n641), .A2(new_n649), .A3(KEYINPUT26), .A4(new_n615), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n712), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n710), .B1(new_n719), .B2(new_n669), .ZN(new_n720));
  AOI211_X1 g0520(.A(KEYINPUT91), .B(new_n668), .C1(new_n712), .C2(new_n718), .ZN(new_n721));
  OAI21_X1  g0521(.A(KEYINPUT29), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT29), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(new_n656), .B2(new_n668), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n709), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n690), .B1(new_n725), .B2(G1), .ZN(G364));
  NOR2_X1   g0526(.A1(G13), .A2(G33), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(G20), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n210), .B1(G20), .B2(new_n419), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n250), .A2(new_n440), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n208), .A2(new_n440), .ZN(new_n733));
  AOI211_X1 g0533(.A(new_n220), .B(new_n284), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(G355), .A2(new_n219), .A3(new_n284), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n735), .B1(G116), .B2(new_n219), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n731), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n662), .A2(G45), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n687), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n211), .A2(G190), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n743), .A2(new_n355), .A3(G200), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n745), .A2(KEYINPUT92), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(KEYINPUT92), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G77), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n211), .A2(new_n382), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n355), .A2(new_n384), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n202), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n384), .A2(G179), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n742), .A2(new_n755), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n756), .A2(new_n350), .B1(new_n757), .B2(new_n365), .ZN(new_n758));
  INV_X1    g0558(.A(new_n751), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n759), .A2(new_n355), .A3(G200), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n754), .B(new_n758), .C1(G58), .C2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G179), .A2(G200), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n211), .B1(new_n762), .B2(G190), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n502), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n752), .A2(new_n742), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n331), .B(new_n764), .C1(G68), .C2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n742), .A2(new_n762), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n323), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT32), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n750), .A2(new_n761), .A3(new_n766), .A4(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n765), .ZN(new_n771));
  XOR2_X1   g0571(.A(KEYINPUT33), .B(G317), .Z(new_n772));
  INV_X1    g0572(.A(G303), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n771), .A2(new_n772), .B1(new_n773), .B2(new_n756), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n284), .B(new_n774), .C1(G311), .C2(new_n744), .ZN(new_n775));
  INV_X1    g0575(.A(G283), .ZN(new_n776));
  INV_X1    g0576(.A(G329), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n757), .A2(new_n776), .B1(new_n767), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n778), .B1(G322), .B2(new_n760), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT94), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT93), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n753), .B(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n434), .A2(new_n435), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n763), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n783), .A2(G326), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n775), .B(new_n779), .C1(new_n780), .C2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n787), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(KEYINPUT94), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n770), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n741), .B1(new_n730), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n729), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n792), .B1(new_n678), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT95), .ZN(new_n795));
  INV_X1    g0595(.A(new_n679), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n740), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(G330), .B2(new_n678), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n795), .A2(new_n798), .ZN(G396));
  NAND2_X1  g0599(.A1(new_n668), .A2(new_n378), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT99), .Z(new_n801));
  OAI21_X1  g0601(.A(new_n379), .B1(new_n801), .B2(new_n386), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n380), .A2(new_n669), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(new_n655), .B2(new_n669), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n668), .B(new_n804), .C1(new_n644), .C2(new_n654), .ZN(new_n807));
  OR3_X1    g0607(.A1(new_n806), .A2(new_n807), .A3(new_n708), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n708), .B1(new_n806), .B2(new_n807), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n808), .A2(new_n739), .A3(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n730), .A2(new_n727), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n811), .B(KEYINPUT96), .Z(new_n812));
  OAI21_X1  g0612(.A(new_n740), .B1(G77), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n550), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n749), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n764), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n756), .A2(new_n365), .B1(new_n757), .B2(new_n350), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n284), .B(new_n817), .C1(G294), .C2(new_n760), .ZN(new_n818));
  INV_X1    g0618(.A(G311), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n771), .A2(new_n776), .B1(new_n767), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n753), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n820), .B1(G303), .B2(new_n821), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n815), .A2(new_n816), .A3(new_n818), .A4(new_n822), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n821), .A2(G137), .B1(new_n765), .B2(G150), .ZN(new_n824));
  INV_X1    g0624(.A(G143), .ZN(new_n825));
  INV_X1    g0625(.A(new_n760), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n824), .B1(new_n825), .B2(new_n826), .C1(new_n748), .C2(new_n323), .ZN(new_n827));
  XNOR2_X1  g0627(.A(KEYINPUT97), .B(KEYINPUT34), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n827), .B(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n756), .ZN(new_n830));
  INV_X1    g0630(.A(new_n757), .ZN(new_n831));
  AOI22_X1  g0631(.A1(G50), .A2(new_n830), .B1(new_n831), .B2(G68), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n338), .B2(new_n763), .ZN(new_n833));
  INV_X1    g0633(.A(G132), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n284), .B1(new_n767), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n835), .A2(KEYINPUT98), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n835), .A2(KEYINPUT98), .ZN(new_n837));
  OR3_X1    g0637(.A1(new_n833), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n823), .B1(new_n829), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n813), .B1(new_n839), .B2(new_n730), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n805), .B2(new_n728), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n810), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT100), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(G384));
  NOR2_X1   g0644(.A1(new_n661), .A2(new_n662), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n406), .A2(new_n669), .ZN(new_n846));
  AND3_X1   g0646(.A1(new_n427), .A2(KEYINPUT101), .A3(new_n430), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT101), .B1(new_n427), .B2(new_n430), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT101), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n431), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n846), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n427), .A2(new_n430), .A3(KEYINPUT101), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n849), .A2(new_n854), .A3(new_n805), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n360), .A2(new_n362), .A3(new_n393), .A4(new_n392), .ZN(new_n856));
  INV_X1    g0656(.A(new_n666), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n345), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n359), .A2(new_n858), .A3(new_n390), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT37), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT37), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n359), .A2(new_n858), .A3(new_n863), .A4(new_n390), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n860), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n337), .A2(new_n340), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n321), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n870), .A2(new_n257), .A3(new_n341), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n666), .B1(new_n871), .B2(new_n344), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n856), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n352), .A2(new_n355), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(G169), .B2(new_n352), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n875), .A2(new_n666), .B1(new_n344), .B2(new_n871), .ZN(new_n876));
  INV_X1    g0676(.A(new_n390), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT37), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n864), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n873), .A2(KEYINPUT38), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n868), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n705), .A2(new_n702), .A3(new_n703), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n855), .A2(KEYINPUT40), .A3(new_n881), .A4(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT40), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n849), .A2(new_n882), .A3(new_n854), .A4(new_n805), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n873), .A2(KEYINPUT38), .A3(new_n879), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT38), .B1(new_n873), .B2(new_n879), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n884), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n883), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n432), .A2(new_n882), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n890), .B(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(G330), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT39), .B1(new_n886), .B2(new_n887), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n868), .A2(new_n897), .A3(new_n880), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n619), .A2(new_n669), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n363), .A2(new_n857), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n849), .A2(new_n854), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n655), .A2(new_n669), .A3(new_n805), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n905), .B1(new_n906), .B2(new_n803), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n887), .B2(new_n886), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n722), .A2(new_n432), .A3(new_n724), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n623), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n909), .B(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n845), .B1(new_n895), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n912), .B2(new_n895), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n209), .B(G77), .C1(new_n338), .C2(new_n326), .ZN(new_n915));
  INV_X1    g0715(.A(G68), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n915), .B1(G50), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(new_n217), .A3(new_n298), .ZN(new_n918));
  OAI211_X1 g0718(.A(G116), .B(new_n212), .C1(new_n506), .C2(KEYINPUT35), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(KEYINPUT35), .B2(new_n506), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n920), .B(KEYINPUT36), .Z(new_n921));
  NAND3_X1  g0721(.A1(new_n914), .A2(new_n918), .A3(new_n921), .ZN(G367));
  OAI211_X1 g0722(.A(new_n541), .B(new_n547), .C1(new_n518), .C2(new_n669), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n684), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT42), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n547), .B1(new_n923), .B2(new_n660), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n924), .A2(new_n925), .B1(new_n669), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(KEYINPUT42), .B1(new_n684), .B2(new_n923), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n669), .A2(new_n614), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n641), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n929), .B1(new_n641), .B2(new_n615), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n927), .A2(new_n928), .B1(KEYINPUT43), .B2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n932), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT43), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n927), .A2(new_n935), .A3(new_n934), .A4(new_n928), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n923), .B1(new_n547), .B2(new_n669), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n681), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n939), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n937), .A2(new_n942), .A3(new_n938), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n686), .B(KEYINPUT41), .Z(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n675), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n679), .B(new_n684), .C1(new_n949), .C2(new_n683), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n670), .B(new_n683), .C1(new_n673), .C2(new_n674), .ZN(new_n951));
  INV_X1    g0751(.A(new_n684), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n796), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n725), .ZN(new_n955));
  AOI211_X1 g0755(.A(KEYINPUT44), .B(new_n940), .C1(new_n684), .C2(new_n682), .ZN(new_n956));
  NOR3_X1   g0756(.A1(new_n675), .A2(new_n679), .A3(KEYINPUT102), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n940), .B1(new_n684), .B2(new_n682), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT44), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n684), .A2(new_n682), .A3(new_n940), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT45), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n684), .A2(KEYINPUT45), .A3(new_n682), .A4(new_n940), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n958), .A2(new_n962), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n681), .A2(KEYINPUT102), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  NOR3_X1   g0771(.A1(new_n961), .A2(new_n956), .A3(new_n957), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n972), .A2(new_n967), .A3(new_n969), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n955), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n725), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n948), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n738), .A2(G1), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n946), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n731), .B1(new_n219), .B2(new_n373), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n220), .A2(new_n284), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n980), .B1(new_n245), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n982), .A2(new_n739), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n748), .A2(new_n202), .B1(new_n323), .B2(new_n771), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n984), .A2(KEYINPUT103), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(KEYINPUT103), .ZN(new_n986));
  INV_X1    g0786(.A(G137), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n284), .B1(new_n763), .B2(new_n916), .C1(new_n987), .C2(new_n767), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n760), .A2(G150), .B1(G77), .B2(new_n831), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n338), .B2(new_n756), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n988), .B(new_n990), .C1(G143), .C2(new_n783), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n985), .A2(new_n986), .A3(new_n991), .ZN(new_n992));
  AND3_X1   g0792(.A1(new_n830), .A2(KEYINPUT46), .A3(G116), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n826), .A2(new_n773), .B1(new_n784), .B2(new_n771), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n993), .B(new_n994), .C1(G97), .C2(new_n831), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n749), .A2(G283), .ZN(new_n996));
  INV_X1    g0796(.A(G317), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n331), .B1(new_n767), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(KEYINPUT46), .B1(new_n830), .B2(new_n814), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n998), .B(new_n999), .C1(G107), .C2(new_n786), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n783), .A2(G311), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n995), .A2(new_n996), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n992), .A2(KEYINPUT47), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n730), .ZN(new_n1004));
  AOI21_X1  g0804(.A(KEYINPUT47), .B1(new_n992), .B2(new_n1002), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n983), .B1(new_n932), .B2(new_n793), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n979), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(G387));
  INV_X1    g0809(.A(new_n955), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n686), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n725), .B2(new_n954), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n242), .A2(G45), .A3(new_n331), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n440), .B1(new_n916), .B2(new_n286), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n270), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT50), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n269), .B2(G50), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1015), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n688), .B1(new_n1019), .B2(new_n284), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n220), .B1(new_n1014), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n731), .B1(new_n365), .B2(new_n219), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n740), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n760), .A2(G317), .B1(G311), .B2(new_n765), .ZN(new_n1024));
  XOR2_X1   g0824(.A(KEYINPUT105), .B(G322), .Z(new_n1025));
  OAI221_X1 g0825(.A(new_n1024), .B1(new_n782), .B2(new_n1025), .C1(new_n748), .C2(new_n773), .ZN(new_n1026));
  AND2_X1   g0826(.A1(new_n1026), .A2(KEYINPUT106), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1026), .A2(KEYINPUT106), .ZN(new_n1028));
  OR3_X1    g0828(.A1(new_n1027), .A2(new_n1028), .A3(KEYINPUT48), .ZN(new_n1029));
  OAI21_X1  g0829(.A(KEYINPUT48), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n785), .A2(new_n830), .B1(G283), .B2(new_n786), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT49), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n742), .A2(G326), .A3(new_n762), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n284), .B1(new_n831), .B2(new_n814), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n763), .A2(new_n373), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(new_n760), .B2(G50), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT104), .ZN(new_n1041));
  INV_X1    g0841(.A(G150), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n745), .A2(new_n916), .B1(new_n767), .B2(new_n1042), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n331), .B(new_n1043), .C1(G97), .C2(new_n831), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n821), .A2(G159), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n830), .A2(G77), .B1(new_n765), .B2(new_n270), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1038), .B1(new_n1041), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1023), .B1(new_n1048), .B2(new_n730), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT107), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n675), .A2(new_n729), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1050), .A2(new_n1051), .B1(new_n954), .B2(new_n977), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1013), .A2(new_n1052), .ZN(G393));
  AOI21_X1  g0853(.A(new_n969), .B1(new_n972), .B2(new_n967), .ZN(new_n1054));
  AND4_X1   g0854(.A1(new_n967), .A2(new_n958), .A3(new_n962), .A4(new_n969), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1010), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n971), .A2(new_n973), .A3(new_n955), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1056), .A2(new_n686), .A3(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n977), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n253), .A2(new_n981), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n731), .B1(new_n502), .B2(new_n219), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n740), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n760), .A2(G159), .B1(new_n821), .B2(G150), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT51), .Z(new_n1064));
  OAI22_X1  g0864(.A1(new_n756), .A2(new_n326), .B1(new_n767), .B2(new_n825), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n284), .B1(new_n763), .B2(new_n286), .C1(new_n350), .C2(new_n757), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(G50), .C2(new_n765), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1064), .B(new_n1067), .C1(new_n269), .C2(new_n748), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1068), .A2(KEYINPUT108), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(KEYINPUT108), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n331), .B1(new_n757), .B2(new_n365), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n745), .A2(new_n433), .B1(new_n773), .B2(new_n771), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(new_n814), .C2(new_n786), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n760), .A2(G311), .B1(new_n821), .B2(G317), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT52), .Z(new_n1075));
  OAI22_X1  g0875(.A1(new_n1025), .A2(new_n767), .B1(new_n756), .B2(new_n776), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT109), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1073), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1069), .A2(new_n1070), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1062), .B1(new_n1079), .B2(new_n730), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n940), .B2(new_n793), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1058), .A2(new_n1059), .A3(new_n1081), .ZN(G390));
  AND2_X1   g0882(.A1(new_n896), .A2(new_n898), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n907), .B2(new_n901), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n709), .A2(new_n855), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n802), .B1(new_n720), .B2(new_n721), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n905), .B1(new_n1086), .B2(new_n803), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n881), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n900), .B(KEYINPUT110), .Z(new_n1089));
  NOR2_X1   g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1084), .B(new_n1085), .C1(new_n1087), .C2(new_n1091), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n849), .A2(new_n854), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n803), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1093), .B1(new_n807), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n899), .B1(new_n1095), .B2(new_n900), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n802), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n719), .A2(new_n669), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(KEYINPUT91), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n719), .A2(new_n710), .A3(new_n669), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1097), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1093), .B1(new_n1101), .B2(new_n1094), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1096), .B1(new_n1102), .B2(new_n1090), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n849), .A2(new_n854), .A3(new_n805), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n882), .A2(G330), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n977), .B(new_n1092), .C1(new_n1103), .C2(new_n1107), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n1108), .A2(KEYINPUT112), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1084), .B1(new_n1087), .B2(new_n1091), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n1106), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT112), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1111), .A2(new_n1112), .A3(new_n977), .A4(new_n1092), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n740), .B1(new_n270), .B2(new_n812), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n771), .A2(new_n365), .B1(new_n767), .B2(new_n433), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(G116), .B2(new_n760), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n748), .B2(new_n502), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n763), .A2(new_n286), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n331), .B1(new_n756), .B2(new_n350), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n753), .A2(new_n776), .B1(new_n757), .B2(new_n916), .ZN(new_n1120));
  NOR4_X1   g0920(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n1121), .A2(KEYINPUT113), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(KEYINPUT113), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n760), .A2(G132), .B1(G50), .B2(new_n831), .ZN(new_n1124));
  INV_X1    g0924(.A(G125), .ZN(new_n1125));
  INV_X1    g0925(.A(G128), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n1124), .B1(new_n1125), .B2(new_n767), .C1(new_n1126), .C2(new_n753), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n284), .B1(new_n323), .B2(new_n763), .C1(new_n771), .C2(new_n987), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n756), .A2(new_n1042), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT53), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT54), .B(G143), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1129), .B(new_n1131), .C1(new_n748), .C2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1122), .A2(new_n1123), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1114), .B1(new_n1134), .B2(new_n730), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n899), .B2(new_n728), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1113), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(KEYINPUT114), .B1(new_n1109), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1108), .A2(KEYINPUT112), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT114), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1139), .A2(new_n1140), .A3(new_n1113), .A4(new_n1136), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1111), .A2(new_n1092), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n432), .A2(G330), .A3(new_n882), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n910), .A2(new_n623), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n807), .A2(new_n1094), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT111), .ZN(new_n1147));
  OAI211_X1 g0947(.A(G330), .B(new_n805), .C1(new_n706), .C2(new_n707), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1147), .B1(new_n1148), .B2(new_n905), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1149), .A2(new_n1106), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1148), .A2(new_n1147), .A3(new_n905), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1146), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n882), .A2(G330), .A3(new_n805), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n709), .A2(new_n855), .B1(new_n905), .B2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1154), .A2(new_n803), .A3(new_n1086), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1145), .B1(new_n1152), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1011), .B1(new_n1142), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n1142), .B2(new_n1157), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1138), .A2(new_n1141), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(KEYINPUT115), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT115), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1138), .A2(new_n1141), .A3(new_n1162), .A4(new_n1159), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(G378));
  NAND3_X1  g0965(.A1(new_n883), .A2(new_n889), .A3(G330), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n279), .A2(new_n666), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n315), .B2(new_n319), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n1167), .B(new_n318), .C1(new_n312), .C2(new_n314), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  XOR2_X1   g0972(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1170), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1173), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1166), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT119), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1180), .A2(new_n883), .A3(new_n889), .A4(G330), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1178), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT120), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(new_n909), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n904), .A2(new_n1183), .A3(new_n908), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(new_n1179), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1178), .A2(new_n1181), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1185), .A2(new_n977), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n739), .B1(new_n202), .B2(new_n811), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT118), .Z(new_n1192));
  INV_X1    g0992(.A(new_n730), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n284), .A2(G41), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(G33), .A2(G41), .ZN(new_n1195));
  OR3_X1    g0995(.A1(new_n1194), .A2(G50), .A3(new_n1195), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n821), .A2(G116), .B1(new_n831), .B2(G58), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1197), .B1(new_n286), .B2(new_n756), .C1(new_n502), .C2(new_n771), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1194), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G107), .B2(new_n760), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1200), .B1(new_n776), .B2(new_n767), .C1(new_n373), .C2(new_n745), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1198), .B(new_n1201), .C1(G68), .C2(new_n786), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1196), .B1(new_n1202), .B2(KEYINPUT58), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT116), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n826), .A2(new_n1126), .B1(new_n834), .B2(new_n771), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n745), .A2(new_n987), .B1(new_n1125), .B2(new_n753), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n756), .A2(new_n1132), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n1208), .A2(KEYINPUT117), .B1(G150), .B2(new_n786), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1207), .B(new_n1209), .C1(KEYINPUT117), .C2(new_n1208), .ZN(new_n1210));
  OR2_X1    g1010(.A1(new_n1210), .A2(KEYINPUT59), .ZN(new_n1211));
  INV_X1    g1011(.A(G124), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1195), .B1(new_n767), .B2(new_n1212), .C1(new_n323), .C2(new_n757), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n1210), .B2(KEYINPUT59), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n1202), .A2(KEYINPUT58), .B1(new_n1211), .B2(new_n1214), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1204), .A2(new_n1215), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1192), .B1(new_n1193), .B2(new_n1216), .C1(new_n1180), .C2(new_n728), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1190), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT121), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1144), .B(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n1142), .B2(new_n1157), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1221), .A2(new_n1185), .A3(new_n1189), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT57), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1188), .A2(new_n908), .A3(new_n904), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n909), .A2(new_n1178), .A3(new_n1181), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1225), .A2(KEYINPUT57), .A3(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1011), .B1(new_n1227), .B2(new_n1221), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1218), .B1(new_n1224), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(G375));
  NAND2_X1  g1030(.A1(new_n1148), .A2(new_n905), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(KEYINPUT111), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1232), .A2(new_n1107), .A3(new_n1151), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1146), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1101), .A2(new_n1094), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1233), .A2(new_n1234), .B1(new_n1235), .B2(new_n1154), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1236), .A2(new_n978), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n748), .A2(new_n365), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n331), .B1(new_n757), .B2(new_n286), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n771), .A2(new_n550), .B1(new_n767), .B2(new_n773), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n753), .A2(new_n433), .B1(new_n756), .B2(new_n502), .ZN(new_n1241));
  NOR4_X1   g1041(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .A4(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1039), .B1(new_n760), .B2(G283), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1243), .B(KEYINPUT122), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n745), .A2(new_n1042), .B1(new_n767), .B2(new_n1126), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n771), .A2(new_n1132), .B1(new_n323), .B2(new_n756), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n284), .B1(new_n757), .B2(new_n338), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n826), .A2(new_n987), .B1(new_n753), .B2(new_n834), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n1248), .B(new_n1249), .C1(G50), .C2(new_n786), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1242), .A2(new_n1244), .B1(new_n1247), .B2(new_n1250), .ZN(new_n1251));
  OAI221_X1 g1051(.A(new_n740), .B1(G68), .B2(new_n812), .C1(new_n1251), .C2(new_n1193), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n905), .B2(new_n727), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1237), .A2(new_n1253), .ZN(new_n1254));
  AND3_X1   g1054(.A1(new_n1148), .A2(new_n1147), .A3(new_n905), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1255), .A2(new_n1149), .A3(new_n1106), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1144), .B(new_n1155), .C1(new_n1256), .C2(new_n1146), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1157), .A2(new_n948), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1254), .A2(new_n1258), .ZN(G381));
  INV_X1    g1059(.A(G396), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1013), .A2(new_n1052), .A3(new_n1260), .ZN(new_n1261));
  NOR4_X1   g1061(.A1(G387), .A2(G384), .A3(G390), .A4(new_n1261), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(G375), .A2(new_n1160), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1262), .A2(new_n1258), .A3(new_n1254), .A4(new_n1263), .ZN(G407));
  INV_X1    g1064(.A(G213), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1265), .A2(G343), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1263), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(G407), .A2(G213), .A3(new_n1267), .ZN(G409));
  AND3_X1   g1068(.A1(new_n1058), .A2(new_n1059), .A3(new_n1081), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n979), .B2(new_n1007), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT125), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1260), .B1(new_n1013), .B2(new_n1052), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1271), .B1(new_n1273), .B2(new_n1261), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1056), .A2(new_n725), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n977), .B1(new_n1275), .B2(new_n948), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1006), .B(G390), .C1(new_n1276), .C2(new_n946), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1270), .A2(new_n1274), .A3(new_n1277), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1008), .A2(G390), .A3(new_n1261), .A4(new_n1273), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n1013), .A2(new_n1052), .A3(new_n1260), .ZN(new_n1280));
  OAI21_X1  g1080(.A(KEYINPUT125), .B1(new_n1280), .B2(new_n1272), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1281), .B(new_n1269), .C1(new_n979), .C2(new_n1007), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1278), .A2(new_n1279), .A3(new_n1282), .ZN(new_n1283));
  XNOR2_X1  g1083(.A(new_n1283), .B(KEYINPUT127), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1161), .A2(new_n1163), .A3(new_n1229), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1225), .A2(new_n977), .A3(new_n1226), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1217), .B(new_n1286), .C1(new_n1222), .C2(new_n947), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1287), .A2(new_n1141), .A3(new_n1138), .A4(new_n1159), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1266), .B1(new_n1285), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT62), .ZN(new_n1290));
  AOI21_X1  g1090(.A(KEYINPUT60), .B1(new_n1236), .B2(new_n1144), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1236), .A2(new_n1144), .ZN(new_n1292));
  OAI21_X1  g1092(.A(KEYINPUT123), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1294), .A2(KEYINPUT60), .A3(new_n1144), .A4(new_n1155), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(KEYINPUT124), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT124), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1236), .A2(new_n1297), .A3(KEYINPUT60), .A4(new_n1144), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1296), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1293), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT60), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1257), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT123), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1302), .A2(new_n1303), .A3(new_n1157), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n686), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1254), .B1(new_n1300), .B2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n843), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1293), .A2(new_n1299), .A3(new_n1304), .A4(new_n686), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1308), .A2(G384), .A3(new_n1254), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1307), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1289), .A2(new_n1290), .A3(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT61), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1309), .ZN(new_n1314));
  AOI21_X1  g1114(.A(G384), .B1(new_n1308), .B2(new_n1254), .ZN(new_n1315));
  OAI211_X1 g1115(.A(G2897), .B(new_n1266), .C1(new_n1314), .C2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(G2897), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1266), .ZN(new_n1318));
  OAI211_X1 g1118(.A(new_n1307), .B(new_n1309), .C1(new_n1317), .C2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1316), .A2(new_n1319), .ZN(new_n1320));
  OAI211_X1 g1120(.A(new_n1312), .B(new_n1313), .C1(new_n1289), .C2(new_n1320), .ZN(new_n1321));
  AOI211_X1 g1121(.A(new_n1266), .B(new_n1310), .C1(new_n1285), .C2(new_n1288), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1322), .A2(new_n1290), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1284), .B1(new_n1321), .B2(new_n1323), .ZN(new_n1324));
  OAI21_X1  g1124(.A(KEYINPUT63), .B1(new_n1289), .B2(new_n1320), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1289), .A2(new_n1311), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1283), .A2(new_n1313), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1328), .B1(new_n1322), .B2(KEYINPUT63), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT126), .ZN(new_n1330));
  AND3_X1   g1130(.A1(new_n1327), .A2(new_n1329), .A3(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1330), .B1(new_n1327), .B2(new_n1329), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1324), .B1(new_n1331), .B2(new_n1332), .ZN(G405));
  XNOR2_X1  g1133(.A(new_n1283), .B(new_n1310), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1285), .B1(new_n1160), .B2(new_n1229), .ZN(new_n1335));
  XNOR2_X1  g1135(.A(new_n1334), .B(new_n1335), .ZN(G402));
endmodule


