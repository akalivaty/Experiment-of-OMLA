

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582;

  XNOR2_X1 U323 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U324 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U325 ( .A(n405), .B(n404), .ZN(n408) );
  XNOR2_X1 U326 ( .A(n445), .B(KEYINPUT123), .ZN(n446) );
  XOR2_X1 U327 ( .A(n416), .B(n415), .Z(n453) );
  XOR2_X1 U328 ( .A(KEYINPUT41), .B(n453), .Z(n546) );
  XOR2_X1 U329 ( .A(n440), .B(n310), .Z(n515) );
  XNOR2_X1 U330 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U331 ( .A(n452), .B(n451), .ZN(G1349GAT) );
  XOR2_X1 U332 ( .A(G183GAT), .B(KEYINPUT83), .Z(n292) );
  XNOR2_X1 U333 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n291) );
  XNOR2_X1 U334 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U335 ( .A(n293), .B(KEYINPUT17), .Z(n295) );
  XNOR2_X1 U336 ( .A(KEYINPUT82), .B(G190GAT), .ZN(n294) );
  XNOR2_X1 U337 ( .A(n295), .B(n294), .ZN(n440) );
  XOR2_X1 U338 ( .A(KEYINPUT20), .B(G99GAT), .Z(n297) );
  XNOR2_X1 U339 ( .A(G43GAT), .B(G15GAT), .ZN(n296) );
  XNOR2_X1 U340 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U341 ( .A(n298), .B(KEYINPUT84), .Z(n300) );
  XOR2_X1 U342 ( .A(G120GAT), .B(G71GAT), .Z(n414) );
  XNOR2_X1 U343 ( .A(G169GAT), .B(n414), .ZN(n299) );
  XNOR2_X1 U344 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U345 ( .A(KEYINPUT80), .B(G176GAT), .Z(n302) );
  NAND2_X1 U346 ( .A1(G227GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U347 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U348 ( .A(n304), .B(n303), .Z(n309) );
  XOR2_X1 U349 ( .A(KEYINPUT79), .B(G134GAT), .Z(n306) );
  XNOR2_X1 U350 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n305) );
  XNOR2_X1 U351 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U352 ( .A(G113GAT), .B(n307), .Z(n344) );
  XNOR2_X1 U353 ( .A(n344), .B(KEYINPUT81), .ZN(n308) );
  XNOR2_X1 U354 ( .A(n309), .B(n308), .ZN(n310) );
  INV_X1 U355 ( .A(n515), .ZN(n525) );
  XOR2_X1 U356 ( .A(G204GAT), .B(KEYINPUT22), .Z(n312) );
  XNOR2_X1 U357 ( .A(G50GAT), .B(KEYINPUT24), .ZN(n311) );
  XNOR2_X1 U358 ( .A(n312), .B(n311), .ZN(n322) );
  XOR2_X1 U359 ( .A(G155GAT), .B(KEYINPUT3), .Z(n314) );
  XNOR2_X1 U360 ( .A(G162GAT), .B(KEYINPUT2), .ZN(n313) );
  XNOR2_X1 U361 ( .A(n314), .B(n313), .ZN(n334) );
  XOR2_X1 U362 ( .A(G141GAT), .B(G22GAT), .Z(n386) );
  XOR2_X1 U363 ( .A(n334), .B(n386), .Z(n316) );
  NAND2_X1 U364 ( .A1(G228GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U365 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U366 ( .A(n317), .B(KEYINPUT85), .Z(n320) );
  XNOR2_X1 U367 ( .A(G106GAT), .B(G78GAT), .ZN(n318) );
  XNOR2_X1 U368 ( .A(n318), .B(G148GAT), .ZN(n406) );
  XNOR2_X1 U369 ( .A(n406), .B(KEYINPUT23), .ZN(n319) );
  XNOR2_X1 U370 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n327) );
  XNOR2_X1 U372 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n323) );
  XNOR2_X1 U373 ( .A(n323), .B(KEYINPUT86), .ZN(n324) );
  XOR2_X1 U374 ( .A(n324), .B(KEYINPUT87), .Z(n326) );
  XNOR2_X1 U375 ( .A(G197GAT), .B(G218GAT), .ZN(n325) );
  XOR2_X1 U376 ( .A(n326), .B(n325), .Z(n435) );
  XNOR2_X1 U377 ( .A(n327), .B(n435), .ZN(n462) );
  XOR2_X1 U378 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n329) );
  XNOR2_X1 U379 ( .A(G141GAT), .B(KEYINPUT89), .ZN(n328) );
  XNOR2_X1 U380 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U381 ( .A(G57GAT), .B(KEYINPUT4), .Z(n331) );
  XNOR2_X1 U382 ( .A(KEYINPUT5), .B(KEYINPUT88), .ZN(n330) );
  XNOR2_X1 U383 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U384 ( .A(n333), .B(n332), .Z(n339) );
  XOR2_X1 U385 ( .A(G85GAT), .B(n334), .Z(n336) );
  XNOR2_X1 U386 ( .A(G29GAT), .B(G148GAT), .ZN(n335) );
  XNOR2_X1 U387 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U388 ( .A(G120GAT), .B(n337), .ZN(n338) );
  XNOR2_X1 U389 ( .A(n339), .B(n338), .ZN(n343) );
  XOR2_X1 U390 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n341) );
  NAND2_X1 U391 ( .A1(G225GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U392 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U393 ( .A(n343), .B(n342), .Z(n346) );
  XNOR2_X1 U394 ( .A(G1GAT), .B(n344), .ZN(n345) );
  XOR2_X1 U395 ( .A(n346), .B(n345), .Z(n461) );
  INV_X1 U396 ( .A(n461), .ZN(n508) );
  INV_X1 U397 ( .A(KEYINPUT54), .ZN(n443) );
  INV_X1 U398 ( .A(KEYINPUT47), .ZN(n421) );
  XOR2_X1 U399 ( .A(G99GAT), .B(G85GAT), .Z(n401) );
  XOR2_X1 U400 ( .A(G162GAT), .B(G218GAT), .Z(n348) );
  XNOR2_X1 U401 ( .A(G134GAT), .B(G190GAT), .ZN(n347) );
  XNOR2_X1 U402 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U403 ( .A(n401), .B(n349), .ZN(n351) );
  AND2_X1 U404 ( .A1(G232GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U405 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U406 ( .A(KEYINPUT9), .B(G92GAT), .Z(n353) );
  XNOR2_X1 U407 ( .A(G36GAT), .B(G106GAT), .ZN(n352) );
  XNOR2_X1 U408 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U409 ( .A(n355), .B(n354), .ZN(n364) );
  XNOR2_X1 U410 ( .A(G43GAT), .B(KEYINPUT67), .ZN(n356) );
  XNOR2_X1 U411 ( .A(n356), .B(G29GAT), .ZN(n357) );
  XOR2_X1 U412 ( .A(n357), .B(KEYINPUT7), .Z(n359) );
  XNOR2_X1 U413 ( .A(G50GAT), .B(KEYINPUT8), .ZN(n358) );
  XNOR2_X1 U414 ( .A(n359), .B(n358), .ZN(n398) );
  XOR2_X1 U415 ( .A(KEYINPUT11), .B(KEYINPUT75), .Z(n361) );
  XNOR2_X1 U416 ( .A(KEYINPUT74), .B(KEYINPUT10), .ZN(n360) );
  XNOR2_X1 U417 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U418 ( .A(n398), .B(n362), .ZN(n363) );
  XNOR2_X1 U419 ( .A(n364), .B(n363), .ZN(n561) );
  INV_X1 U420 ( .A(n561), .ZN(n554) );
  XOR2_X1 U421 ( .A(G78GAT), .B(G71GAT), .Z(n366) );
  XNOR2_X1 U422 ( .A(G127GAT), .B(G183GAT), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U424 ( .A(G57GAT), .B(KEYINPUT13), .Z(n413) );
  XOR2_X1 U425 ( .A(n367), .B(n413), .Z(n369) );
  XNOR2_X1 U426 ( .A(G22GAT), .B(G211GAT), .ZN(n368) );
  XNOR2_X1 U427 ( .A(n369), .B(n368), .ZN(n374) );
  XNOR2_X1 U428 ( .A(G15GAT), .B(G1GAT), .ZN(n370) );
  XNOR2_X1 U429 ( .A(n370), .B(KEYINPUT68), .ZN(n394) );
  XOR2_X1 U430 ( .A(n394), .B(KEYINPUT12), .Z(n372) );
  NAND2_X1 U431 ( .A1(G231GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U432 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U433 ( .A(n374), .B(n373), .Z(n382) );
  XOR2_X1 U434 ( .A(KEYINPUT78), .B(G64GAT), .Z(n376) );
  XNOR2_X1 U435 ( .A(G8GAT), .B(G155GAT), .ZN(n375) );
  XNOR2_X1 U436 ( .A(n376), .B(n375), .ZN(n380) );
  XOR2_X1 U437 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n378) );
  XNOR2_X1 U438 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n377) );
  XNOR2_X1 U439 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U440 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U441 ( .A(n382), .B(n381), .Z(n576) );
  INV_X1 U442 ( .A(n576), .ZN(n551) );
  NAND2_X1 U443 ( .A1(n554), .A2(n551), .ZN(n419) );
  XOR2_X1 U444 ( .A(KEYINPUT64), .B(KEYINPUT66), .Z(n384) );
  XNOR2_X1 U445 ( .A(G113GAT), .B(G197GAT), .ZN(n383) );
  XNOR2_X1 U446 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U447 ( .A(n386), .B(n385), .Z(n388) );
  NAND2_X1 U448 ( .A1(G229GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U449 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U450 ( .A(KEYINPUT30), .B(KEYINPUT69), .Z(n390) );
  XNOR2_X1 U451 ( .A(KEYINPUT29), .B(KEYINPUT65), .ZN(n389) );
  XNOR2_X1 U452 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U453 ( .A(n392), .B(n391), .Z(n396) );
  XNOR2_X1 U454 ( .A(G169GAT), .B(G36GAT), .ZN(n393) );
  XNOR2_X1 U455 ( .A(n393), .B(G8GAT), .ZN(n436) );
  XNOR2_X1 U456 ( .A(n436), .B(n394), .ZN(n395) );
  XNOR2_X1 U457 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U458 ( .A(n398), .B(n397), .Z(n569) );
  XOR2_X1 U459 ( .A(G64GAT), .B(G92GAT), .Z(n400) );
  XNOR2_X1 U460 ( .A(G176GAT), .B(G204GAT), .ZN(n399) );
  XNOR2_X1 U461 ( .A(n400), .B(n399), .ZN(n433) );
  XNOR2_X1 U462 ( .A(n433), .B(n401), .ZN(n405) );
  AND2_X1 U463 ( .A1(G230GAT), .A2(G233GAT), .ZN(n403) );
  INV_X1 U464 ( .A(KEYINPUT33), .ZN(n402) );
  XNOR2_X1 U465 ( .A(n406), .B(KEYINPUT31), .ZN(n407) );
  XNOR2_X1 U466 ( .A(n408), .B(n407), .ZN(n412) );
  XOR2_X1 U467 ( .A(KEYINPUT32), .B(KEYINPUT73), .Z(n410) );
  XNOR2_X1 U468 ( .A(KEYINPUT72), .B(KEYINPUT71), .ZN(n409) );
  XOR2_X1 U469 ( .A(n410), .B(n409), .Z(n411) );
  XNOR2_X1 U470 ( .A(n412), .B(n411), .ZN(n416) );
  XNOR2_X1 U471 ( .A(n414), .B(n413), .ZN(n415) );
  NOR2_X1 U472 ( .A1(n569), .A2(n546), .ZN(n417) );
  XNOR2_X1 U473 ( .A(n417), .B(KEYINPUT46), .ZN(n418) );
  NOR2_X1 U474 ( .A1(n419), .A2(n418), .ZN(n420) );
  XNOR2_X1 U475 ( .A(n421), .B(n420), .ZN(n429) );
  XOR2_X1 U476 ( .A(KEYINPUT70), .B(n569), .Z(n557) );
  INV_X1 U477 ( .A(n453), .ZN(n572) );
  XOR2_X1 U478 ( .A(KEYINPUT45), .B(KEYINPUT108), .Z(n423) );
  XNOR2_X1 U479 ( .A(n554), .B(KEYINPUT36), .ZN(n579) );
  NOR2_X1 U480 ( .A1(n551), .A2(n579), .ZN(n422) );
  XNOR2_X1 U481 ( .A(n423), .B(n422), .ZN(n424) );
  NOR2_X1 U482 ( .A1(n572), .A2(n424), .ZN(n425) );
  XNOR2_X1 U483 ( .A(n425), .B(KEYINPUT109), .ZN(n426) );
  NOR2_X1 U484 ( .A1(n557), .A2(n426), .ZN(n427) );
  XNOR2_X1 U485 ( .A(KEYINPUT110), .B(n427), .ZN(n428) );
  NOR2_X1 U486 ( .A1(n429), .A2(n428), .ZN(n430) );
  XNOR2_X1 U487 ( .A(n430), .B(KEYINPUT48), .ZN(n522) );
  XOR2_X1 U488 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n432) );
  NAND2_X1 U489 ( .A1(G226GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U490 ( .A(n432), .B(n431), .ZN(n434) );
  XOR2_X1 U491 ( .A(n434), .B(n433), .Z(n438) );
  XOR2_X1 U492 ( .A(n436), .B(n435), .Z(n437) );
  XNOR2_X1 U493 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X2 U494 ( .A(n440), .B(n439), .Z(n511) );
  XOR2_X1 U495 ( .A(KEYINPUT122), .B(n511), .Z(n441) );
  NOR2_X1 U496 ( .A1(n522), .A2(n441), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n444) );
  NOR2_X1 U498 ( .A1(n508), .A2(n444), .ZN(n568) );
  AND2_X1 U499 ( .A1(n462), .A2(n568), .ZN(n447) );
  INV_X1 U500 ( .A(KEYINPUT55), .ZN(n445) );
  NOR2_X1 U501 ( .A1(n525), .A2(n448), .ZN(n562) );
  INV_X1 U502 ( .A(n546), .ZN(n529) );
  NAND2_X1 U503 ( .A1(n562), .A2(n529), .ZN(n452) );
  XOR2_X1 U504 ( .A(G176GAT), .B(KEYINPUT56), .Z(n450) );
  XNOR2_X1 U505 ( .A(KEYINPUT124), .B(KEYINPUT57), .ZN(n449) );
  NAND2_X1 U506 ( .A1(n557), .A2(n453), .ZN(n483) );
  NOR2_X1 U507 ( .A1(n551), .A2(n561), .ZN(n454) );
  XNOR2_X1 U508 ( .A(KEYINPUT16), .B(n454), .ZN(n468) );
  NAND2_X1 U509 ( .A1(n515), .A2(n511), .ZN(n455) );
  NAND2_X1 U510 ( .A1(n462), .A2(n455), .ZN(n456) );
  XOR2_X1 U511 ( .A(KEYINPUT25), .B(n456), .Z(n459) );
  XNOR2_X1 U512 ( .A(n511), .B(KEYINPUT27), .ZN(n463) );
  NOR2_X1 U513 ( .A1(n462), .A2(n515), .ZN(n457) );
  XNOR2_X1 U514 ( .A(n457), .B(KEYINPUT26), .ZN(n567) );
  NAND2_X1 U515 ( .A1(n463), .A2(n567), .ZN(n458) );
  NAND2_X1 U516 ( .A1(n459), .A2(n458), .ZN(n460) );
  NAND2_X1 U517 ( .A1(n461), .A2(n460), .ZN(n466) );
  XOR2_X1 U518 ( .A(KEYINPUT28), .B(n462), .Z(n518) );
  INV_X1 U519 ( .A(n518), .ZN(n524) );
  NAND2_X1 U520 ( .A1(n508), .A2(n463), .ZN(n521) );
  NOR2_X1 U521 ( .A1(n515), .A2(n521), .ZN(n464) );
  NAND2_X1 U522 ( .A1(n524), .A2(n464), .ZN(n465) );
  NAND2_X1 U523 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U524 ( .A(KEYINPUT94), .B(n467), .ZN(n478) );
  NAND2_X1 U525 ( .A1(n468), .A2(n478), .ZN(n494) );
  NOR2_X1 U526 ( .A1(n483), .A2(n494), .ZN(n476) );
  NAND2_X1 U527 ( .A1(n476), .A2(n508), .ZN(n472) );
  XOR2_X1 U528 ( .A(KEYINPUT34), .B(KEYINPUT96), .Z(n470) );
  XNOR2_X1 U529 ( .A(G1GAT), .B(KEYINPUT95), .ZN(n469) );
  XNOR2_X1 U530 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U531 ( .A(n472), .B(n471), .ZN(G1324GAT) );
  NAND2_X1 U532 ( .A1(n476), .A2(n511), .ZN(n473) );
  XNOR2_X1 U533 ( .A(n473), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U534 ( .A(G15GAT), .B(KEYINPUT35), .Z(n475) );
  NAND2_X1 U535 ( .A1(n476), .A2(n515), .ZN(n474) );
  XNOR2_X1 U536 ( .A(n475), .B(n474), .ZN(G1326GAT) );
  NAND2_X1 U537 ( .A1(n518), .A2(n476), .ZN(n477) );
  XNOR2_X1 U538 ( .A(n477), .B(G22GAT), .ZN(G1327GAT) );
  AND2_X1 U539 ( .A1(n551), .A2(n478), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n479), .B(KEYINPUT97), .ZN(n480) );
  NOR2_X1 U541 ( .A1(n579), .A2(n480), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n481), .B(KEYINPUT98), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n482), .B(KEYINPUT37), .ZN(n507) );
  NOR2_X1 U544 ( .A1(n483), .A2(n507), .ZN(n484) );
  XNOR2_X1 U545 ( .A(n484), .B(KEYINPUT38), .ZN(n490) );
  NAND2_X1 U546 ( .A1(n508), .A2(n490), .ZN(n486) );
  XOR2_X1 U547 ( .A(G29GAT), .B(KEYINPUT39), .Z(n485) );
  XNOR2_X1 U548 ( .A(n486), .B(n485), .ZN(G1328GAT) );
  NAND2_X1 U549 ( .A1(n490), .A2(n511), .ZN(n487) );
  XNOR2_X1 U550 ( .A(n487), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U551 ( .A1(n490), .A2(n515), .ZN(n488) );
  XNOR2_X1 U552 ( .A(n488), .B(KEYINPUT40), .ZN(n489) );
  XNOR2_X1 U553 ( .A(G43GAT), .B(n489), .ZN(G1330GAT) );
  NAND2_X1 U554 ( .A1(n518), .A2(n490), .ZN(n491) );
  XNOR2_X1 U555 ( .A(G50GAT), .B(n491), .ZN(G1331GAT) );
  XNOR2_X1 U556 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n492) );
  XNOR2_X1 U557 ( .A(n492), .B(KEYINPUT100), .ZN(n493) );
  XOR2_X1 U558 ( .A(KEYINPUT99), .B(n493), .Z(n496) );
  NAND2_X1 U559 ( .A1(n569), .A2(n529), .ZN(n506) );
  NOR2_X1 U560 ( .A1(n506), .A2(n494), .ZN(n501) );
  NAND2_X1 U561 ( .A1(n501), .A2(n508), .ZN(n495) );
  XNOR2_X1 U562 ( .A(n496), .B(n495), .ZN(G1332GAT) );
  NAND2_X1 U563 ( .A1(n501), .A2(n511), .ZN(n497) );
  XNOR2_X1 U564 ( .A(n497), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n499) );
  NAND2_X1 U566 ( .A1(n501), .A2(n515), .ZN(n498) );
  XNOR2_X1 U567 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U568 ( .A(G71GAT), .B(n500), .ZN(G1334GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT104), .B(KEYINPUT43), .Z(n503) );
  NAND2_X1 U570 ( .A1(n501), .A2(n518), .ZN(n502) );
  XNOR2_X1 U571 ( .A(n503), .B(n502), .ZN(n505) );
  XOR2_X1 U572 ( .A(G78GAT), .B(KEYINPUT103), .Z(n504) );
  XNOR2_X1 U573 ( .A(n505), .B(n504), .ZN(G1335GAT) );
  XOR2_X1 U574 ( .A(G85GAT), .B(KEYINPUT105), .Z(n510) );
  NOR2_X1 U575 ( .A1(n507), .A2(n506), .ZN(n517) );
  NAND2_X1 U576 ( .A1(n517), .A2(n508), .ZN(n509) );
  XNOR2_X1 U577 ( .A(n510), .B(n509), .ZN(G1336GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n513) );
  NAND2_X1 U579 ( .A1(n517), .A2(n511), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U581 ( .A(G92GAT), .B(n514), .ZN(G1337GAT) );
  NAND2_X1 U582 ( .A1(n517), .A2(n515), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n516), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U584 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n519), .B(KEYINPUT44), .ZN(n520) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n520), .ZN(G1339GAT) );
  NOR2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n523) );
  XOR2_X1 U588 ( .A(KEYINPUT111), .B(n523), .Z(n541) );
  NAND2_X1 U589 ( .A1(n541), .A2(n524), .ZN(n526) );
  NOR2_X1 U590 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U591 ( .A(n527), .B(KEYINPUT112), .ZN(n536) );
  NAND2_X1 U592 ( .A1(n536), .A2(n557), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n528), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT49), .B(KEYINPUT113), .Z(n531) );
  NAND2_X1 U595 ( .A1(n529), .A2(n536), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U597 ( .A(G120GAT), .B(n532), .Z(G1341GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n534) );
  NAND2_X1 U599 ( .A1(n536), .A2(n576), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U601 ( .A(G127GAT), .B(n535), .Z(G1342GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n538) );
  NAND2_X1 U603 ( .A1(n536), .A2(n561), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(n540) );
  XOR2_X1 U605 ( .A(G134GAT), .B(KEYINPUT115), .Z(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  NAND2_X1 U607 ( .A1(n541), .A2(n567), .ZN(n553) );
  NOR2_X1 U608 ( .A1(n569), .A2(n553), .ZN(n543) );
  XNOR2_X1 U609 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(G1344GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT120), .B(KEYINPUT119), .Z(n545) );
  XNOR2_X1 U612 ( .A(KEYINPUT52), .B(KEYINPUT53), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(n550) );
  NOR2_X1 U614 ( .A1(n546), .A2(n553), .ZN(n548) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(G1345GAT) );
  NOR2_X1 U618 ( .A1(n551), .A2(n553), .ZN(n552) );
  XOR2_X1 U619 ( .A(G155GAT), .B(n552), .Z(G1346GAT) );
  NOR2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n556) );
  XNOR2_X1 U621 ( .A(G162GAT), .B(KEYINPUT121), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1347GAT) );
  NAND2_X1 U623 ( .A1(n557), .A2(n562), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G169GAT), .B(n558), .ZN(G1348GAT) );
  XOR2_X1 U625 ( .A(G183GAT), .B(KEYINPUT125), .Z(n560) );
  NAND2_X1 U626 ( .A1(n562), .A2(n576), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1350GAT) );
  XNOR2_X1 U628 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n564) );
  NAND2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1351GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT126), .B(KEYINPUT59), .Z(n566) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n571) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n578) );
  NOR2_X1 U635 ( .A1(n569), .A2(n578), .ZN(n570) );
  XOR2_X1 U636 ( .A(n571), .B(n570), .Z(G1352GAT) );
  XOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .Z(n574) );
  INV_X1 U638 ( .A(n578), .ZN(n575) );
  NAND2_X1 U639 ( .A1(n575), .A2(n572), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n577), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U644 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

