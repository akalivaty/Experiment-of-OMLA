//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0 1 0 0 0 0 1 0 0 1 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n853, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980;
  INV_X1    g000(.A(KEYINPUT90), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT36), .ZN(new_n203));
  XOR2_X1   g002(.A(G15gat), .B(G43gat), .Z(new_n204));
  XNOR2_X1  g003(.A(G71gat), .B(G99gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G227gat), .A2(G233gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT26), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT67), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT67), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n213), .A2(new_n217), .A3(new_n214), .ZN(new_n218));
  INV_X1    g017(.A(G183gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT27), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT27), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G183gat), .ZN(new_n222));
  INV_X1    g021(.A(G190gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n220), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT28), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(KEYINPUT27), .B(G183gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(KEYINPUT28), .A3(new_n223), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n216), .A2(new_n218), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT25), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(new_n214), .ZN(new_n233));
  NAND3_X1  g032(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n212), .A2(KEYINPUT23), .ZN(new_n236));
  INV_X1    g035(.A(G169gat), .ZN(new_n237));
  INV_X1    g036(.A(G176gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n235), .A2(new_n240), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n208), .A2(KEYINPUT64), .A3(KEYINPUT23), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT64), .B1(new_n208), .B2(KEYINPUT23), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n231), .B1(new_n241), .B2(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n231), .B1(new_n208), .B2(KEYINPUT23), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n240), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT65), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n234), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g048(.A1(KEYINPUT65), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n249), .A2(new_n250), .B1(new_n214), .B2(new_n232), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT66), .B1(new_n245), .B2(new_n252), .ZN(new_n253));
  AOI22_X1  g052(.A1(new_n233), .A2(new_n234), .B1(new_n239), .B2(new_n236), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n237), .A2(new_n238), .A3(KEYINPUT23), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT64), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n208), .A2(KEYINPUT64), .A3(KEYINPUT23), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT25), .B1(new_n254), .B2(new_n259), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n247), .A2(new_n251), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT66), .ZN(new_n262));
  NOR3_X1   g061(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n230), .B1(new_n253), .B2(new_n263), .ZN(new_n264));
  XOR2_X1   g063(.A(G127gat), .B(G134gat), .Z(new_n265));
  XNOR2_X1  g064(.A(G113gat), .B(G120gat), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n266), .A2(KEYINPUT68), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT1), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n268), .B1(new_n266), .B2(KEYINPUT68), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n265), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n265), .A2(KEYINPUT1), .ZN(new_n271));
  INV_X1    g070(.A(G120gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(G113gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT69), .B(G113gat), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n273), .B1(new_n274), .B2(new_n272), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT70), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n270), .A2(new_n279), .A3(new_n276), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n245), .A2(new_n252), .A3(KEYINPUT66), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n262), .B1(new_n260), .B2(new_n261), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n285), .A2(new_n278), .A3(new_n280), .A4(new_n230), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n207), .B1(new_n282), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n206), .B1(new_n287), .B2(KEYINPUT33), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT32), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n282), .A2(new_n286), .ZN(new_n292));
  INV_X1    g091(.A(new_n207), .ZN(new_n293));
  AOI221_X4 g092(.A(new_n289), .B1(KEYINPUT33), .B2(new_n206), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT71), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n282), .A2(new_n207), .A3(new_n286), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT34), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  NOR3_X1   g097(.A1(new_n291), .A2(new_n298), .A3(new_n294), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n296), .B(KEYINPUT34), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n264), .A2(new_n281), .ZN(new_n301));
  AOI22_X1  g100(.A1(new_n285), .A2(new_n230), .B1(new_n278), .B2(new_n280), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n293), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT32), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT33), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n304), .A2(new_n306), .A3(new_n206), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n288), .A2(new_n290), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n300), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n295), .B1(new_n299), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n307), .A2(new_n308), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n311), .A2(KEYINPUT71), .A3(new_n300), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n203), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n298), .B1(new_n291), .B2(new_n294), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n307), .A2(new_n308), .A3(new_n300), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n316), .A2(KEYINPUT36), .ZN(new_n317));
  NAND2_X1  g116(.A1(G228gat), .A2(G233gat), .ZN(new_n318));
  XOR2_X1   g117(.A(new_n318), .B(KEYINPUT81), .Z(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G197gat), .B(G204gat), .ZN(new_n321));
  INV_X1    g120(.A(G211gat), .ZN(new_n322));
  INV_X1    g121(.A(G218gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n321), .B1(KEYINPUT22), .B2(new_n324), .ZN(new_n325));
  XOR2_X1   g124(.A(G211gat), .B(G218gat), .Z(new_n326));
  XNOR2_X1  g125(.A(new_n325), .B(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT29), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT3), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT77), .ZN(new_n331));
  XNOR2_X1  g130(.A(KEYINPUT74), .B(G141gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G148gat), .ZN(new_n333));
  OR2_X1    g132(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n334), .A2(G141gat), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G155gat), .ZN(new_n338));
  INV_X1    g137(.A(G162gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(G155gat), .A2(G162gat), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT2), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n337), .A2(new_n345), .ZN(new_n346));
  XOR2_X1   g145(.A(G141gat), .B(G148gat), .Z(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n343), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n340), .A2(new_n342), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n331), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  AOI211_X1 g150(.A(new_n340), .B(new_n342), .C1(new_n347), .C2(new_n343), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n333), .A2(new_n336), .B1(new_n341), .B2(new_n344), .ZN(new_n353));
  NOR3_X1   g152(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT77), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n330), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n352), .A2(new_n353), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT3), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT29), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OR2_X1    g157(.A1(new_n358), .A2(new_n327), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n320), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  OAI211_X1 g159(.A(G228gat), .B(G233gat), .C1(new_n329), .C2(new_n356), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n358), .A2(new_n327), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(G22gat), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n354), .A2(new_n351), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n365), .A2(new_n329), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n319), .B1(new_n366), .B2(new_n362), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT82), .B(G22gat), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n367), .B(new_n368), .C1(new_n362), .C2(new_n361), .ZN(new_n369));
  XNOR2_X1  g168(.A(G78gat), .B(G106gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT31), .B(G50gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  AND3_X1   g171(.A1(new_n364), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n372), .B(KEYINPUT80), .ZN(new_n374));
  INV_X1    g173(.A(new_n368), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n375), .B1(new_n360), .B2(new_n363), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n374), .B1(new_n376), .B2(new_n369), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(G225gat), .A2(G233gat), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT76), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n277), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n346), .A2(new_n350), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT3), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n270), .A2(KEYINPUT76), .A3(new_n276), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n346), .A2(new_n357), .A3(new_n350), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n382), .A2(new_n384), .A3(new_n385), .A4(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT4), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n270), .A2(new_n279), .A3(new_n276), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n279), .B1(new_n270), .B2(new_n276), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n388), .B1(new_n391), .B2(new_n365), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n356), .A2(new_n388), .A3(new_n270), .A4(new_n276), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT78), .ZN(new_n394));
  INV_X1    g193(.A(new_n277), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT78), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n395), .A2(new_n396), .A3(new_n388), .A4(new_n356), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n380), .B(new_n387), .C1(new_n392), .C2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT5), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n382), .A2(new_n383), .A3(new_n385), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n395), .A2(new_n356), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n380), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n400), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT4), .B1(new_n391), .B2(new_n365), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n395), .A2(KEYINPUT4), .A3(new_n356), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n387), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n404), .A2(KEYINPUT5), .ZN(new_n410));
  AOI22_X1  g209(.A1(new_n399), .A2(new_n405), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  XOR2_X1   g210(.A(G1gat), .B(G29gat), .Z(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G57gat), .B(G85gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT6), .B1(new_n411), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n406), .ZN(new_n419));
  INV_X1    g218(.A(new_n408), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n419), .A2(new_n420), .A3(new_n410), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n387), .A2(new_n380), .ZN(new_n422));
  INV_X1    g221(.A(new_n398), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n391), .A2(new_n365), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT4), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n422), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n403), .A2(new_n404), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT5), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n421), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n416), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n418), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n429), .A2(KEYINPUT6), .A3(new_n416), .ZN(new_n432));
  XNOR2_X1  g231(.A(G8gat), .B(G36gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(G64gat), .B(G92gat), .ZN(new_n434));
  XOR2_X1   g233(.A(new_n433), .B(new_n434), .Z(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n245), .A2(new_n252), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n230), .ZN(new_n438));
  NAND2_X1  g237(.A1(G226gat), .A2(G233gat), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n216), .A2(new_n218), .A3(new_n229), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n443), .B1(new_n284), .B2(new_n283), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n439), .B1(new_n444), .B2(KEYINPUT29), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n442), .B1(new_n445), .B2(KEYINPUT72), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT72), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n447), .B(new_n439), .C1(new_n444), .C2(KEYINPUT29), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n327), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n327), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n285), .A2(new_n440), .A3(new_n230), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n438), .A2(new_n328), .A3(new_n439), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n436), .B1(new_n449), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT29), .B1(new_n285), .B2(new_n230), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT72), .B1(new_n455), .B2(new_n440), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n456), .A2(new_n448), .A3(new_n441), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n450), .ZN(new_n458));
  INV_X1    g257(.A(new_n453), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n458), .A2(new_n459), .A3(new_n435), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT30), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n461), .A2(KEYINPUT73), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n454), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n453), .B1(new_n457), .B2(new_n450), .ZN(new_n464));
  XNOR2_X1  g263(.A(KEYINPUT73), .B(KEYINPUT30), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(new_n435), .A3(new_n465), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n431), .A2(new_n432), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  OAI22_X1  g266(.A1(new_n313), .A2(new_n317), .B1(new_n379), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n463), .A2(new_n466), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT83), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT86), .B1(new_n411), .B2(new_n417), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT86), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n429), .A2(new_n472), .A3(new_n416), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n404), .B1(new_n406), .B2(new_n408), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  XOR2_X1   g275(.A(KEYINPUT84), .B(KEYINPUT39), .Z(new_n477));
  AOI21_X1  g276(.A(new_n416), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT85), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n479), .B1(new_n403), .B2(new_n404), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n401), .A2(KEYINPUT85), .A3(new_n402), .A4(new_n380), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n475), .A2(KEYINPUT39), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT40), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT40), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n478), .A2(new_n485), .A3(new_n482), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n474), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT83), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n463), .A2(new_n488), .A3(new_n466), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n470), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT37), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n436), .B1(new_n464), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT89), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g293(.A(KEYINPUT89), .B(new_n436), .C1(new_n464), .C2(new_n491), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT38), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n496), .B1(new_n464), .B2(new_n491), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n451), .A2(new_n450), .A3(new_n452), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT88), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT88), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n451), .A2(new_n452), .A3(new_n501), .A4(new_n450), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n456), .A2(new_n327), .A3(new_n448), .A4(new_n441), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n503), .B1(KEYINPUT87), .B2(new_n504), .ZN(new_n505));
  OR2_X1    g304(.A1(new_n504), .A2(KEYINPUT87), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n491), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n458), .A2(new_n491), .A3(new_n459), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(new_n436), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n496), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n498), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n471), .A2(new_n418), .A3(new_n473), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n512), .A2(new_n432), .A3(new_n460), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n378), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n468), .B1(new_n490), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT35), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(new_n373), .B2(new_n377), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n517), .B1(new_n512), .B2(new_n432), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n463), .A2(new_n488), .A3(new_n466), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n488), .B1(new_n463), .B2(new_n466), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n518), .B(new_n316), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n378), .B1(new_n310), .B2(new_n312), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n516), .B1(new_n523), .B2(new_n467), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n202), .B1(new_n515), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n513), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n527), .A2(new_n490), .A3(new_n379), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n314), .A2(new_n315), .B1(KEYINPUT71), .B2(new_n311), .ZN(new_n529));
  INV_X1    g328(.A(new_n312), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT36), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n317), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n431), .A2(new_n432), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(new_n469), .ZN(new_n534));
  AOI22_X1  g333(.A1(new_n531), .A2(new_n532), .B1(new_n534), .B2(new_n378), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n528), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n536), .B(KEYINPUT90), .C1(new_n524), .C2(new_n522), .ZN(new_n537));
  XOR2_X1   g336(.A(KEYINPUT91), .B(G29gat), .Z(new_n538));
  XOR2_X1   g337(.A(KEYINPUT92), .B(G36gat), .Z(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NOR3_X1   g341(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n540), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G43gat), .B(G50gat), .Z(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n544), .A2(KEYINPUT15), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT93), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n543), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n543), .A2(new_n548), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n542), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n546), .A2(KEYINPUT15), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT15), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n545), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n552), .A2(new_n540), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n547), .B1(new_n551), .B2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT17), .ZN(new_n557));
  XNOR2_X1  g356(.A(G15gat), .B(G22gat), .ZN(new_n558));
  AND2_X1   g357(.A1(KEYINPUT94), .A2(G1gat), .ZN(new_n559));
  OAI21_X1  g358(.A(KEYINPUT16), .B1(KEYINPUT94), .B2(G1gat), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n561), .B(KEYINPUT95), .C1(G1gat), .C2(new_n558), .ZN(new_n562));
  INV_X1    g361(.A(G8gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n557), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G229gat), .A2(G233gat), .ZN(new_n566));
  INV_X1    g365(.A(new_n564), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(new_n556), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n565), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT18), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n564), .B(new_n556), .Z(new_n571));
  XOR2_X1   g370(.A(new_n566), .B(KEYINPUT13), .Z(new_n572));
  AOI22_X1  g371(.A1(new_n569), .A2(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n565), .A2(KEYINPUT18), .A3(new_n566), .A4(new_n568), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G113gat), .B(G141gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(G197gat), .ZN(new_n577));
  XOR2_X1   g376(.A(KEYINPUT11), .B(G169gat), .Z(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n579), .B(KEYINPUT12), .Z(new_n580));
  NAND2_X1  g379(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n580), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n573), .A2(new_n582), .A3(new_n574), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT96), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n581), .A2(KEYINPUT96), .A3(new_n583), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n526), .A2(new_n537), .A3(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(G71gat), .A2(G78gat), .ZN(new_n590));
  NOR2_X1   g389(.A1(G71gat), .A2(G78gat), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G57gat), .B(G64gat), .Z(new_n593));
  AOI21_X1  g392(.A(new_n592), .B1(new_n593), .B2(KEYINPUT97), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n593), .B1(KEYINPUT9), .B2(new_n590), .ZN(new_n595));
  OR2_X1    g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n595), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n598), .A2(KEYINPUT21), .ZN(new_n599));
  NAND2_X1  g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(G127gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n567), .B1(KEYINPUT21), .B2(new_n598), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(G155gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(G183gat), .B(G211gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n605), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT99), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT7), .ZN(new_n615));
  OAI211_X1 g414(.A(G85gat), .B(G92gat), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT100), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n618), .B1(KEYINPUT99), .B2(KEYINPUT7), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n616), .B(KEYINPUT100), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n620), .A2(new_n614), .A3(new_n615), .ZN(new_n621));
  NAND2_X1  g420(.A1(G99gat), .A2(G106gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(KEYINPUT8), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n623), .B1(G85gat), .B2(G92gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT101), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n619), .A2(new_n621), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(G99gat), .B(G106gat), .Z(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n627), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n619), .A2(new_n621), .A3(new_n629), .A4(new_n625), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n628), .A2(new_n556), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT41), .ZN(new_n632));
  NAND2_X1  g431(.A1(G232gat), .A2(G233gat), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n628), .A2(new_n630), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n634), .B1(new_n557), .B2(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(G190gat), .B(G218gat), .Z(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n633), .A2(new_n632), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT98), .ZN(new_n640));
  XOR2_X1   g439(.A(G134gat), .B(G162gat), .Z(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n638), .A2(new_n642), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(KEYINPUT102), .B1(new_n613), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n645), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n647), .A2(new_n612), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n598), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT10), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n628), .A2(new_n598), .A3(new_n630), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  OR2_X1    g454(.A1(new_n654), .A2(new_n653), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n655), .A2(KEYINPUT103), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT103), .B1(new_n655), .B2(new_n656), .ZN(new_n659));
  NAND2_X1  g458(.A1(G230gat), .A2(G233gat), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n658), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n652), .A2(new_n654), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n661), .ZN(new_n665));
  XNOR2_X1  g464(.A(G120gat), .B(G148gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(G176gat), .B(G204gat), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n666), .B(new_n667), .Z(new_n668));
  NAND3_X1  g467(.A1(new_n663), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n655), .A2(new_n656), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(new_n660), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n665), .ZN(new_n672));
  INV_X1    g471(.A(new_n668), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n650), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n589), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n677), .A2(new_n533), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n678), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g478(.A1(new_n519), .A2(new_n520), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT104), .B(KEYINPUT16), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(G8gat), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n685), .A2(KEYINPUT42), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(KEYINPUT42), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n686), .B(new_n687), .C1(new_n563), .C2(new_n682), .ZN(G1325gat));
  NOR2_X1   g487(.A1(new_n313), .A2(new_n317), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(G15gat), .B1(new_n677), .B2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n316), .ZN(new_n692));
  OR2_X1    g491(.A1(new_n692), .A2(G15gat), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n691), .B1(new_n677), .B2(new_n693), .ZN(G1326gat));
  NOR2_X1   g493(.A1(new_n677), .A2(new_n379), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT105), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT43), .B(G22gat), .Z(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1327gat));
  INV_X1    g497(.A(new_n675), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n589), .A2(new_n613), .A3(new_n645), .A4(new_n699), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n700), .A2(new_n533), .A3(new_n538), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n701), .B(KEYINPUT45), .Z(new_n702));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n703), .B1(new_n522), .B2(new_n524), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n379), .B1(new_n529), .B2(new_n530), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT35), .B1(new_n705), .B2(new_n534), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n706), .A2(KEYINPUT108), .A3(new_n521), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n704), .A2(new_n536), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n645), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n647), .A2(new_n710), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n526), .A2(new_n537), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n675), .B(KEYINPUT107), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT106), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n584), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n581), .A2(KEYINPUT106), .A3(new_n583), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n716), .A2(new_n613), .A3(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n714), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n538), .B1(new_n723), .B2(new_n533), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n702), .A2(new_n724), .ZN(G1328gat));
  NOR3_X1   g524(.A1(new_n700), .A2(new_n681), .A3(new_n539), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT46), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n539), .B1(new_n723), .B2(new_n681), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(G1329gat));
  NAND3_X1  g528(.A1(new_n722), .A2(G43gat), .A3(new_n689), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n700), .A2(new_n692), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n730), .B1(new_n731), .B2(G43gat), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g532(.A(G50gat), .B1(new_n723), .B2(new_n379), .ZN(new_n734));
  AOI21_X1  g533(.A(KEYINPUT48), .B1(new_n734), .B2(KEYINPUT109), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n379), .A2(G50gat), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n700), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n735), .B(new_n737), .ZN(G1331gat));
  NOR3_X1   g537(.A1(new_n650), .A2(new_n716), .A3(new_n720), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n739), .A2(new_n708), .ZN(new_n740));
  INV_X1    g539(.A(new_n533), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g542(.A1(new_n740), .A2(new_n680), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n745));
  XOR2_X1   g544(.A(KEYINPUT49), .B(G64gat), .Z(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n744), .B2(new_n746), .ZN(G1333gat));
  NAND3_X1  g546(.A1(new_n740), .A2(G71gat), .A3(new_n689), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT110), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n740), .A2(new_n316), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(G71gat), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g551(.A1(new_n740), .A2(new_n378), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g553(.A1(new_n720), .A2(new_n612), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n675), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT111), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n711), .A2(new_n713), .A3(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(G85gat), .B1(new_n759), .B2(new_n533), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n708), .A2(new_n645), .A3(new_n755), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n708), .A2(KEYINPUT51), .A3(new_n645), .A4(new_n755), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n699), .A2(G85gat), .A3(new_n533), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT112), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n760), .B1(new_n766), .B2(new_n768), .ZN(G1336gat));
  INV_X1    g568(.A(KEYINPUT115), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n711), .A2(new_n680), .A3(new_n713), .A4(new_n757), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G92gat), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n716), .A2(G92gat), .A3(new_n681), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n765), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n772), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  AOI22_X1  g578(.A1(G92gat), .A2(new_n771), .B1(new_n765), .B2(new_n774), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT113), .B1(new_n780), .B2(new_n773), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n772), .A2(KEYINPUT113), .A3(new_n775), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT52), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n770), .B(new_n779), .C1(new_n781), .C2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n778), .B1(new_n780), .B2(KEYINPUT113), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n776), .A2(new_n777), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n770), .B1(new_n788), .B2(new_n779), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n785), .A2(new_n789), .ZN(G1337gat));
  OAI21_X1  g589(.A(G99gat), .B1(new_n759), .B2(new_n690), .ZN(new_n791));
  OR3_X1    g590(.A1(new_n699), .A2(G99gat), .A3(new_n692), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n766), .B2(new_n792), .ZN(G1338gat));
  NAND2_X1  g592(.A1(new_n758), .A2(new_n378), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(G106gat), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT116), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n379), .A2(G106gat), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n765), .A2(new_n715), .A3(new_n800), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n795), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n799), .B1(new_n795), .B2(new_n801), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n798), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n795), .A2(new_n801), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(KEYINPUT117), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT53), .B1(new_n795), .B2(KEYINPUT116), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n795), .A2(new_n799), .A3(new_n801), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n804), .A2(new_n809), .ZN(G1339gat));
  AOI21_X1  g609(.A(new_n566), .B1(new_n565), .B2(new_n568), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n571), .A2(new_n572), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n579), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n583), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n675), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n673), .B1(new_n671), .B2(KEYINPUT54), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(KEYINPUT54), .B1(new_n670), .B2(new_n660), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n817), .B1(new_n662), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n817), .B(KEYINPUT55), .C1(new_n662), .C2(new_n818), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n821), .A2(new_n669), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n718), .A2(new_n719), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n815), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT118), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI211_X1 g626(.A(KEYINPUT118), .B(new_n815), .C1(new_n823), .C2(new_n824), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n827), .A2(new_n647), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n823), .A2(new_n647), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n814), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n612), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n650), .A2(new_n675), .A3(new_n720), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n834), .A2(new_n379), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n680), .A2(new_n692), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n835), .A2(new_n741), .A3(new_n836), .A4(new_n588), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n837), .A2(KEYINPUT119), .A3(G113gat), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(KEYINPUT119), .B1(new_n837), .B2(G113gat), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n835), .A2(new_n741), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n680), .B1(new_n312), .B2(new_n310), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n824), .A2(new_n274), .ZN(new_n845));
  OAI22_X1  g644(.A1(new_n839), .A2(new_n840), .B1(new_n844), .B2(new_n845), .ZN(G1340gat));
  NAND4_X1  g645(.A1(new_n835), .A2(new_n741), .A3(new_n836), .A4(new_n715), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(KEYINPUT120), .A3(G120gat), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT120), .B1(new_n847), .B2(G120gat), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n675), .A2(new_n272), .ZN(new_n851));
  OAI22_X1  g650(.A1(new_n849), .A2(new_n850), .B1(new_n844), .B2(new_n851), .ZN(G1341gat));
  NAND2_X1  g651(.A1(new_n842), .A2(new_n836), .ZN(new_n853));
  OAI21_X1  g652(.A(G127gat), .B1(new_n853), .B2(new_n613), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n612), .A2(new_n602), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n854), .B1(new_n844), .B2(new_n855), .ZN(G1342gat));
  XOR2_X1   g655(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n647), .A2(G134gat), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n858), .B1(new_n844), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(G134gat), .B1(new_n853), .B2(new_n647), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n842), .A2(new_n843), .A3(new_n859), .A4(new_n857), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(G1343gat));
  INV_X1    g663(.A(KEYINPUT58), .ZN(new_n865));
  INV_X1    g664(.A(new_n332), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n867), .B(new_n378), .C1(new_n832), .C2(new_n833), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n689), .A2(new_n533), .A3(new_n680), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n822), .A2(new_n669), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n871));
  AOI21_X1  g670(.A(KEYINPUT55), .B1(new_n819), .B2(new_n871), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n817), .B(KEYINPUT122), .C1(new_n662), .C2(new_n818), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT123), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n659), .A2(new_n661), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n818), .B1(new_n875), .B2(new_n657), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n871), .B1(new_n876), .B2(new_n816), .ZN(new_n877));
  AND4_X1   g676(.A1(KEYINPUT123), .A2(new_n873), .A3(new_n877), .A4(new_n820), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n588), .B(new_n870), .C1(new_n874), .C2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n645), .B1(new_n879), .B2(new_n815), .ZN(new_n880));
  INV_X1    g679(.A(new_n831), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n613), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(new_n833), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n379), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n868), .B(new_n869), .C1(new_n884), .C2(new_n867), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n866), .B1(new_n885), .B2(new_n824), .ZN(new_n886));
  INV_X1    g685(.A(new_n588), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n887), .A2(G141gat), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n834), .A2(new_n378), .A3(new_n869), .A4(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n865), .B1(new_n886), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n865), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n882), .A2(new_n883), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n378), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(KEYINPUT57), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n894), .A2(new_n588), .A3(new_n868), .A4(new_n869), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n891), .B1(new_n895), .B2(new_n866), .ZN(new_n896));
  OAI21_X1  g695(.A(KEYINPUT124), .B1(new_n890), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n866), .B1(new_n885), .B2(new_n887), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n865), .A3(new_n889), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT124), .ZN(new_n900));
  INV_X1    g699(.A(new_n889), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n894), .A2(new_n720), .A3(new_n868), .A4(new_n869), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n901), .B1(new_n902), .B2(new_n866), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n899), .B(new_n900), .C1(new_n903), .C2(new_n865), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n897), .A2(new_n904), .ZN(G1344gat));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n834), .A2(new_n378), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT57), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n879), .A2(new_n815), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n647), .ZN(new_n910));
  OR3_X1    g709(.A1(new_n823), .A2(KEYINPUT125), .A3(new_n647), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT125), .B1(new_n823), .B2(new_n647), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(new_n814), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n612), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n650), .A2(new_n588), .A3(new_n675), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n867), .B(new_n378), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n908), .A2(new_n916), .A3(new_n675), .A4(new_n869), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n906), .B1(new_n917), .B2(G148gat), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n885), .A2(new_n699), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n334), .A2(new_n335), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n919), .A2(KEYINPUT59), .A3(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n907), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(new_n869), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n675), .A2(new_n921), .ZN(new_n925));
  OAI22_X1  g724(.A1(new_n918), .A2(new_n922), .B1(new_n924), .B2(new_n925), .ZN(G1345gat));
  OAI21_X1  g725(.A(G155gat), .B1(new_n885), .B2(new_n613), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n612), .A2(new_n338), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n924), .B2(new_n928), .ZN(G1346gat));
  OAI21_X1  g728(.A(G162gat), .B1(new_n885), .B2(new_n647), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n645), .A2(new_n339), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n930), .B1(new_n924), .B2(new_n931), .ZN(G1347gat));
  NOR2_X1   g731(.A1(new_n681), .A2(new_n741), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n934), .A2(new_n692), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n835), .A2(new_n935), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n936), .A2(new_n237), .A3(new_n887), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n834), .A2(new_n523), .A3(new_n933), .ZN(new_n938));
  AOI21_X1  g737(.A(G169gat), .B1(new_n938), .B2(new_n720), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n937), .A2(new_n939), .ZN(G1348gat));
  OAI21_X1  g739(.A(G176gat), .B1(new_n936), .B2(new_n716), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n938), .A2(new_n238), .A3(new_n675), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(G1349gat));
  OAI21_X1  g742(.A(G183gat), .B1(new_n936), .B2(new_n613), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n938), .A2(new_n227), .A3(new_n612), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(KEYINPUT60), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT60), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n944), .A2(new_n948), .A3(new_n945), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n949), .ZN(G1350gat));
  NAND3_X1  g749(.A1(new_n938), .A2(new_n223), .A3(new_n645), .ZN(new_n951));
  OAI21_X1  g750(.A(G190gat), .B1(new_n936), .B2(new_n647), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n952), .A2(KEYINPUT61), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n952), .A2(KEYINPUT61), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(G1351gat));
  AND2_X1   g754(.A1(new_n908), .A2(new_n916), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n934), .A2(new_n689), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(G197gat), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n887), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n923), .A2(new_n957), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT126), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n923), .A2(KEYINPUT126), .A3(new_n957), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n964), .A2(new_n720), .A3(new_n965), .ZN(new_n966));
  AOI22_X1  g765(.A1(new_n959), .A2(new_n961), .B1(new_n966), .B2(new_n960), .ZN(G1352gat));
  NOR2_X1   g766(.A1(new_n699), .A2(G204gat), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n923), .A2(new_n957), .A3(new_n968), .ZN(new_n969));
  XOR2_X1   g768(.A(new_n969), .B(KEYINPUT62), .Z(new_n970));
  OAI21_X1  g769(.A(G204gat), .B1(new_n958), .B2(new_n716), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(G1353gat));
  NAND4_X1  g771(.A1(new_n908), .A2(new_n916), .A3(new_n612), .A4(new_n957), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n973), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT63), .B1(new_n973), .B2(G211gat), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n964), .A2(new_n965), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n612), .A2(new_n322), .ZN(new_n977));
  OAI22_X1  g776(.A1(new_n974), .A2(new_n975), .B1(new_n976), .B2(new_n977), .ZN(G1354gat));
  OAI21_X1  g777(.A(G218gat), .B1(new_n958), .B2(new_n647), .ZN(new_n979));
  NAND4_X1  g778(.A1(new_n964), .A2(new_n323), .A3(new_n645), .A4(new_n965), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(G1355gat));
endmodule


