//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 0 0 0 1 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G140), .ZN(new_n189));
  INV_X1    g003(.A(G227), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G953), .ZN(new_n191));
  XOR2_X1   g005(.A(new_n189), .B(new_n191), .Z(new_n192));
  INV_X1    g006(.A(G101), .ZN(new_n193));
  INV_X1    g007(.A(G104), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G107), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G104), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n193), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT80), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n199), .B1(new_n196), .B2(G104), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT3), .B1(new_n194), .B2(G107), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(new_n196), .A3(G104), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n194), .A2(KEYINPUT80), .A3(G107), .ZN(new_n204));
  AND4_X1   g018(.A1(new_n200), .A2(new_n201), .A3(new_n203), .A4(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n198), .B1(new_n205), .B2(new_n193), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  AND2_X1   g021(.A1(KEYINPUT64), .A2(G143), .ZN(new_n208));
  NOR2_X1   g022(.A1(KEYINPUT64), .A2(G143), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT1), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n207), .A2(KEYINPUT65), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G146), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(new_n214), .A3(G143), .ZN(new_n215));
  OR2_X1    g029(.A1(KEYINPUT64), .A2(G143), .ZN(new_n216));
  NAND2_X1  g030(.A1(KEYINPUT64), .A2(G143), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(G146), .A3(new_n217), .ZN(new_n218));
  AOI22_X1  g032(.A1(new_n211), .A2(G128), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT1), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n218), .A2(new_n215), .A3(new_n220), .A4(G128), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n206), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT10), .ZN(new_n224));
  AOI21_X1  g038(.A(G146), .B1(new_n216), .B2(new_n217), .ZN(new_n225));
  AOI21_X1  g039(.A(G143), .B1(new_n212), .B2(new_n214), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G128), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n228), .B1(new_n215), .B2(KEYINPUT1), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n221), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n198), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n200), .A2(new_n201), .A3(new_n203), .A4(new_n204), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n231), .B(KEYINPUT10), .C1(new_n232), .C2(G101), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n223), .A2(new_n224), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  XOR2_X1   g049(.A(KEYINPUT82), .B(KEYINPUT4), .Z(new_n236));
  INV_X1    g050(.A(KEYINPUT81), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n201), .A2(new_n203), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n194), .A2(KEYINPUT80), .A3(G107), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT80), .B1(new_n194), .B2(G107), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n237), .B1(new_n238), .B2(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n232), .A2(KEYINPUT81), .ZN(new_n243));
  OAI211_X1 g057(.A(G101), .B(new_n236), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  XOR2_X1   g058(.A(KEYINPUT0), .B(G128), .Z(new_n245));
  OAI21_X1  g059(.A(new_n245), .B1(new_n225), .B2(new_n226), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n218), .A2(new_n215), .A3(KEYINPUT0), .A4(G128), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n205), .A2(new_n237), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n232), .A2(KEYINPUT81), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n193), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(KEYINPUT4), .B1(new_n232), .B2(G101), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n244), .B(new_n248), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n235), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT11), .ZN(new_n255));
  INV_X1    g069(.A(G134), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n255), .B1(new_n256), .B2(G137), .ZN(new_n257));
  INV_X1    g071(.A(G137), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT11), .A3(G134), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n256), .A2(G137), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G131), .ZN(new_n262));
  INV_X1    g076(.A(G131), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n257), .A2(new_n259), .A3(new_n263), .A4(new_n260), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n254), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT83), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n254), .A2(KEYINPUT83), .A3(new_n265), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n265), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n235), .A2(new_n253), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n192), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(KEYINPUT65), .B(G146), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n220), .B1(new_n274), .B2(G143), .ZN(new_n275));
  OAI22_X1  g089(.A1(new_n275), .A2(new_n228), .B1(new_n225), .B2(new_n226), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n231), .B1(new_n232), .B2(G101), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(new_n221), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n271), .B1(new_n223), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT12), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n279), .B(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n272), .A2(new_n192), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n187), .B(new_n188), .C1(new_n273), .C2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n282), .B1(new_n268), .B2(new_n269), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n279), .B(KEYINPUT12), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n192), .B1(new_n286), .B2(new_n272), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n188), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT84), .B1(new_n288), .B2(G469), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n272), .A2(new_n192), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT83), .B1(new_n254), .B2(new_n265), .ZN(new_n291));
  AOI211_X1 g105(.A(new_n267), .B(new_n271), .C1(new_n235), .C2(new_n253), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n192), .ZN(new_n294));
  INV_X1    g108(.A(new_n272), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n294), .B1(new_n281), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(G902), .B1(new_n293), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT84), .ZN(new_n298));
  NOR3_X1   g112(.A1(new_n297), .A2(new_n298), .A3(new_n187), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n284), .B1(new_n289), .B2(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT9), .B(G234), .ZN(new_n301));
  OAI21_X1  g115(.A(G221), .B1(new_n301), .B2(G902), .ZN(new_n302));
  XOR2_X1   g116(.A(new_n302), .B(KEYINPUT79), .Z(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(G113), .B(G122), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n305), .B(new_n194), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n216), .A2(new_n217), .ZN(new_n307));
  INV_X1    g121(.A(G237), .ZN(new_n308));
  INV_X1    g122(.A(G953), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n308), .A2(new_n309), .A3(G214), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT88), .ZN(new_n311));
  NOR2_X1   g125(.A1(G237), .A2(G953), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G214), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT88), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n307), .B1(new_n311), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n310), .A2(G143), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  OAI211_X1 g132(.A(KEYINPUT18), .B(G131), .C1(new_n316), .C2(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n208), .A2(new_n209), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n313), .A2(new_n314), .ZN(new_n321));
  AOI21_X1  g135(.A(KEYINPUT88), .B1(new_n312), .B2(G214), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(KEYINPUT18), .A2(G131), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(new_n317), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G140), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G125), .ZN(new_n327));
  INV_X1    g141(.A(G125), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G140), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n274), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n331), .B1(new_n207), .B2(new_n330), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n319), .A2(new_n325), .A3(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(G131), .B1(new_n316), .B2(new_n318), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT17), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n323), .A2(new_n263), .A3(new_n317), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  OAI211_X1 g151(.A(KEYINPUT17), .B(G131), .C1(new_n316), .C2(new_n318), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n327), .A2(new_n329), .A3(KEYINPUT16), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT76), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n327), .A2(new_n329), .A3(KEYINPUT76), .A4(KEYINPUT16), .ZN(new_n342));
  OR2_X1    g156(.A1(new_n327), .A2(KEYINPUT16), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n207), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n341), .A2(G146), .A3(new_n342), .A4(new_n343), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n338), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n306), .B(new_n333), .C1(new_n337), .C2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n350), .A2(new_n345), .A3(new_n346), .A4(new_n338), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n306), .B1(new_n351), .B2(new_n333), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n188), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G475), .ZN(new_n354));
  INV_X1    g168(.A(new_n306), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n319), .A2(new_n325), .A3(new_n332), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n327), .A2(new_n329), .A3(KEYINPUT19), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT19), .B1(new_n327), .B2(new_n329), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n274), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n346), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n360), .B1(new_n334), .B2(new_n336), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n355), .B1(new_n356), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n348), .ZN(new_n363));
  NOR2_X1   g177(.A1(G475), .A2(G902), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n363), .B(new_n364), .C1(KEYINPUT89), .C2(KEYINPUT20), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n354), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT91), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n363), .A2(new_n364), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n363), .A2(KEYINPUT89), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT20), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n320), .A2(G128), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n228), .A2(G143), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n256), .A3(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(G116), .B(G122), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(new_n196), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n373), .B1(new_n307), .B2(new_n228), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT13), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(G134), .B1(new_n372), .B2(KEYINPUT13), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n374), .B(new_n376), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G122), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G116), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n196), .B1(new_n383), .B2(KEYINPUT14), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(new_n375), .ZN(new_n385));
  INV_X1    g199(.A(new_n374), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n256), .B1(new_n372), .B2(new_n373), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G217), .ZN(new_n389));
  NOR3_X1   g203(.A1(new_n301), .A2(new_n389), .A3(G953), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n381), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n390), .B1(new_n381), .B2(new_n388), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n188), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G478), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n394), .A2(KEYINPUT15), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n395), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n188), .B(new_n397), .C1(new_n391), .C2(new_n392), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  AOI211_X1 g213(.A(new_n188), .B(new_n309), .C1(G234), .C2(G237), .ZN(new_n400));
  XNOR2_X1  g214(.A(KEYINPUT21), .B(G898), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OR2_X1    g216(.A1(KEYINPUT90), .A2(G952), .ZN(new_n403));
  NAND2_X1  g217(.A1(KEYINPUT90), .A2(G952), .ZN(new_n404));
  AOI21_X1  g218(.A(G953), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G234), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n405), .B1(new_n406), .B2(new_n308), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n399), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n366), .A2(new_n367), .A3(new_n371), .A4(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n371), .A2(new_n354), .A3(new_n365), .ZN(new_n411));
  INV_X1    g225(.A(new_n409), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT91), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(G214), .B1(G237), .B2(G902), .ZN(new_n415));
  XOR2_X1   g229(.A(new_n415), .B(KEYINPUT85), .Z(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT2), .ZN(new_n418));
  INV_X1    g232(.A(G113), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT67), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT67), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(KEYINPUT2), .A3(G113), .ZN(new_n422));
  AOI22_X1  g236(.A1(new_n420), .A2(new_n422), .B1(new_n418), .B2(new_n419), .ZN(new_n423));
  XNOR2_X1  g237(.A(G116), .B(G119), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n423), .B(new_n424), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n244), .B(new_n425), .C1(new_n251), .C2(new_n252), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n420), .A2(new_n422), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n418), .A2(new_n419), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n428), .A3(new_n424), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n424), .A2(KEYINPUT5), .ZN(new_n430));
  INV_X1    g244(.A(G116), .ZN(new_n431));
  NOR3_X1   g245(.A1(new_n431), .A2(KEYINPUT5), .A3(G119), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n432), .A2(new_n419), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n206), .A2(new_n429), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n426), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(G110), .B(G122), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n426), .A2(new_n435), .A3(new_n437), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(KEYINPUT6), .A3(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT6), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n436), .A2(new_n442), .A3(new_n438), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n246), .A2(G125), .A3(new_n247), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n230), .A2(new_n328), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n309), .A2(G224), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n447), .B(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n441), .A2(new_n443), .A3(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G210), .B1(G237), .B2(G902), .ZN(new_n451));
  XOR2_X1   g265(.A(new_n437), .B(KEYINPUT8), .Z(new_n452));
  INV_X1    g266(.A(new_n429), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n277), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT86), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n433), .A2(new_n455), .B1(KEYINPUT5), .B2(new_n424), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n456), .B1(new_n455), .B2(new_n433), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n434), .A2(new_n429), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n277), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT87), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n454), .A2(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n458), .A2(KEYINPUT87), .A3(new_n277), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n452), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(G125), .B1(new_n276), .B2(new_n221), .ZN(new_n464));
  OAI211_X1 g278(.A(KEYINPUT7), .B(new_n448), .C1(new_n464), .C2(new_n444), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n448), .A2(KEYINPUT7), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n445), .A2(new_n446), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(G902), .B1(new_n469), .B2(new_n440), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n450), .A2(new_n451), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n451), .B1(new_n450), .B2(new_n470), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n417), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n300), .A2(new_n304), .A3(new_n414), .A4(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT92), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n474), .B1(new_n410), .B2(new_n413), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n479), .A2(KEYINPUT92), .A3(new_n304), .A4(new_n300), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n260), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n256), .A2(G137), .ZN(new_n483));
  OAI21_X1  g297(.A(G131), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n264), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n485), .B1(new_n276), .B2(new_n221), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n265), .A2(new_n247), .A3(new_n246), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n425), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n485), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n230), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n423), .A2(new_n424), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n453), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n265), .A2(new_n247), .A3(new_n246), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n490), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n488), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(KEYINPUT28), .ZN(new_n496));
  AOI21_X1  g310(.A(KEYINPUT72), .B1(new_n490), .B2(new_n493), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n490), .A2(KEYINPUT72), .A3(new_n493), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n425), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n496), .B1(new_n500), .B2(KEYINPUT28), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT27), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n312), .A2(new_n502), .A3(G210), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n502), .B1(new_n312), .B2(G210), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT69), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n505), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT69), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n508), .A3(new_n503), .ZN(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT26), .B(G101), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n506), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n510), .B1(new_n506), .B2(new_n509), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(KEYINPUT29), .B1(new_n501), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT28), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n516), .B1(new_n488), .B2(new_n494), .ZN(new_n517));
  INV_X1    g331(.A(new_n499), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n492), .B1(new_n518), .B2(new_n497), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n517), .B1(new_n519), .B2(new_n516), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT29), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n513), .B(KEYINPUT71), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n515), .A2(new_n524), .ZN(new_n525));
  XOR2_X1   g339(.A(KEYINPUT66), .B(KEYINPUT30), .Z(new_n526));
  OAI21_X1  g340(.A(new_n526), .B1(new_n486), .B2(new_n487), .ZN(new_n527));
  NOR2_X1   g341(.A1(KEYINPUT66), .A2(KEYINPUT30), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n490), .A2(new_n493), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(KEYINPUT68), .B1(new_n530), .B2(new_n425), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT68), .ZN(new_n532));
  AOI211_X1 g346(.A(new_n532), .B(new_n492), .C1(new_n527), .C2(new_n529), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n513), .B1(new_n534), .B2(new_n494), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n188), .B1(new_n525), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(G472), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n494), .A2(KEYINPUT70), .A3(new_n513), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT70), .B1(new_n494), .B2(new_n513), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n540), .B1(new_n531), .B2(new_n533), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT31), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT73), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n543), .B1(new_n520), .B2(new_n523), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n501), .A2(KEYINPUT73), .A3(new_n522), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT31), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n540), .B(new_n546), .C1(new_n531), .C2(new_n533), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n542), .A2(new_n544), .A3(new_n545), .A4(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT32), .ZN(new_n549));
  NOR2_X1   g363(.A1(G472), .A2(G902), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n549), .B1(new_n548), .B2(new_n550), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n537), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT74), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n345), .A2(new_n346), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n228), .A2(G119), .ZN(new_n556));
  INV_X1    g370(.A(G119), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(G128), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT24), .B(G110), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT23), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n562), .B1(new_n557), .B2(G128), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n228), .A2(KEYINPUT23), .A3(G119), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n558), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(G110), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT75), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n565), .A2(KEYINPUT75), .A3(G110), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n561), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n555), .A2(new_n570), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n559), .A2(new_n560), .ZN(new_n572));
  XOR2_X1   g386(.A(KEYINPUT77), .B(G110), .Z(new_n573));
  NOR2_X1   g387(.A1(new_n565), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n346), .B(new_n331), .C1(new_n572), .C2(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(KEYINPUT22), .B(G137), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n309), .A2(G221), .A3(G234), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n571), .A2(new_n575), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n579), .B1(new_n571), .B2(new_n575), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n188), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n188), .B(new_n583), .C1(new_n580), .C2(new_n581), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n389), .B1(G234), .B2(new_n188), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n587), .A2(G902), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n589), .B1(new_n580), .B2(new_n581), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT74), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n537), .B(new_n593), .C1(new_n551), .C2(new_n552), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n554), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n481), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(new_n193), .ZN(G3));
  INV_X1    g411(.A(KEYINPUT33), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n598), .B1(new_n391), .B2(new_n392), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n394), .A2(G902), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT95), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT94), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n381), .A2(new_n388), .ZN(new_n603));
  INV_X1    g417(.A(new_n390), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n381), .A2(new_n388), .A3(new_n390), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(KEYINPUT33), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n392), .A2(new_n602), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n601), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI211_X1 g424(.A(KEYINPUT33), .B(new_n606), .C1(new_n392), .C2(new_n602), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n392), .A2(new_n602), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n611), .A2(new_n612), .A3(KEYINPUT95), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n599), .B(new_n600), .C1(new_n610), .C2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT96), .B(G478), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n393), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n617), .A2(new_n411), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n471), .A2(KEYINPUT93), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n450), .A2(new_n470), .ZN(new_n620));
  INV_X1    g434(.A(new_n451), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT93), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n450), .A2(new_n470), .A3(new_n623), .A4(new_n451), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n619), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n408), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n618), .A2(new_n625), .A3(new_n626), .A4(new_n417), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT97), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n548), .A2(new_n188), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(G472), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n548), .A2(new_n550), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n288), .A2(KEYINPUT84), .A3(G469), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n298), .B1(new_n297), .B2(new_n187), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n272), .B1(new_n291), .B2(new_n292), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n294), .ZN(new_n637));
  INV_X1    g451(.A(new_n283), .ZN(new_n638));
  AOI21_X1  g452(.A(G902), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AOI22_X1  g453(.A1(new_n634), .A2(new_n635), .B1(new_n187), .B2(new_n639), .ZN(new_n640));
  NOR4_X1   g454(.A1(new_n633), .A2(new_n640), .A3(new_n591), .A4(new_n303), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n629), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  NAND2_X1  g458(.A1(new_n625), .A2(new_n417), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n354), .A2(new_n399), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n368), .B(KEYINPUT20), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(new_n408), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n641), .A2(new_n646), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT98), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT35), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT99), .B(G107), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  NAND2_X1  g469(.A1(new_n571), .A2(new_n575), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n656), .B1(KEYINPUT36), .B2(new_n579), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n579), .A2(KEYINPUT36), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n571), .A2(new_n575), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n589), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n588), .A2(KEYINPUT100), .A3(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(KEYINPUT100), .B1(new_n588), .B2(new_n662), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n633), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n478), .A2(new_n480), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT101), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT102), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT37), .B(G110), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G12));
  INV_X1    g486(.A(new_n407), .ZN(new_n673));
  INV_X1    g487(.A(G900), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n673), .B1(new_n674), .B2(new_n400), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n647), .A2(new_n648), .A3(new_n676), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n640), .A2(new_n677), .A3(new_n303), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n645), .A2(new_n666), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n554), .A2(new_n678), .A3(new_n594), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G128), .ZN(G30));
  XNOR2_X1  g495(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n675), .B(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n300), .A2(new_n304), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n684), .B(KEYINPUT40), .Z(new_n685));
  NAND2_X1  g499(.A1(new_n632), .A2(KEYINPUT32), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI22_X1  g502(.A1(new_n534), .A2(new_n540), .B1(new_n495), .B2(new_n522), .ZN(new_n689));
  OAI21_X1  g503(.A(G472), .B1(new_n689), .B2(G902), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n472), .A2(new_n473), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT38), .ZN(new_n693));
  INV_X1    g507(.A(new_n666), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n411), .A2(new_n399), .ZN(new_n695));
  NOR4_X1   g509(.A1(new_n693), .A2(new_n416), .A3(new_n694), .A4(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n685), .A2(new_n691), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(new_n307), .ZN(G45));
  NAND3_X1  g512(.A1(new_n617), .A2(new_n411), .A3(new_n676), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n640), .A2(new_n303), .A3(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n554), .A2(new_n594), .A3(new_n700), .A4(new_n679), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G146), .ZN(G48));
  INV_X1    g516(.A(new_n302), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n283), .B1(new_n636), .B2(new_n294), .ZN(new_n704));
  OAI21_X1  g518(.A(G469), .B1(new_n704), .B2(G902), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT104), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n284), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  OAI211_X1 g521(.A(KEYINPUT104), .B(G469), .C1(new_n704), .C2(G902), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n703), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n554), .A2(new_n592), .A3(new_n594), .A4(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n710), .A2(new_n628), .ZN(new_n711));
  XOR2_X1   g525(.A(KEYINPUT41), .B(G113), .Z(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G15));
  NAND2_X1  g527(.A1(new_n646), .A2(new_n650), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(new_n431), .ZN(G18));
  AOI221_X4 g530(.A(new_n703), .B1(new_n410), .B2(new_n413), .C1(new_n707), .C2(new_n708), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n717), .A2(new_n554), .A3(new_n594), .A4(new_n679), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G119), .ZN(G21));
  AOI211_X1 g533(.A(new_n703), .B(new_n408), .C1(new_n707), .C2(new_n708), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n695), .A2(KEYINPUT106), .ZN(new_n721));
  OR2_X1    g535(.A1(new_n695), .A2(KEYINPUT106), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n645), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(G472), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n724), .B1(new_n548), .B2(new_n188), .ZN(new_n725));
  INV_X1    g539(.A(new_n550), .ZN(new_n726));
  AOI22_X1  g540(.A1(new_n541), .A2(KEYINPUT31), .B1(new_n501), .B2(new_n522), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n726), .B1(new_n727), .B2(new_n547), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(KEYINPUT105), .B1(new_n729), .B2(new_n592), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT105), .ZN(new_n731));
  NOR4_X1   g545(.A1(new_n725), .A2(new_n731), .A3(new_n728), .A4(new_n591), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n720), .B(new_n723), .C1(new_n730), .C2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G122), .ZN(G24));
  NOR4_X1   g548(.A1(new_n666), .A2(new_n725), .A3(new_n699), .A4(new_n728), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n646), .A3(new_n709), .ZN(new_n736));
  XOR2_X1   g550(.A(KEYINPUT107), .B(G125), .Z(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G27));
  XNOR2_X1  g552(.A(KEYINPUT109), .B(KEYINPUT42), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n622), .A2(new_n417), .A3(new_n471), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT108), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n288), .A2(G469), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n284), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n622), .A2(KEYINPUT108), .A3(new_n417), .A4(new_n471), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n742), .A2(new_n302), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n554), .A2(new_n747), .A3(new_n592), .A4(new_n594), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n739), .B1(new_n748), .B2(new_n699), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT42), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n699), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n553), .A2(new_n592), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g566(.A(KEYINPUT110), .B1(new_n752), .B2(new_n746), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n591), .B1(new_n688), .B2(new_n537), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT110), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n754), .A2(new_n747), .A3(new_n755), .A4(new_n751), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n749), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G131), .ZN(G33));
  NOR2_X1   g573(.A1(new_n748), .A2(new_n677), .ZN(new_n760));
  XNOR2_X1  g574(.A(KEYINPUT111), .B(G134), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(G36));
  NAND2_X1  g576(.A1(new_n293), .A2(new_n296), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(KEYINPUT112), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n187), .B1(new_n763), .B2(new_n764), .ZN(new_n767));
  AOI22_X1  g581(.A1(new_n766), .A2(new_n767), .B1(G469), .B2(G902), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n768), .A2(KEYINPUT46), .ZN(new_n769));
  AOI22_X1  g583(.A1(new_n768), .A2(KEYINPUT46), .B1(new_n187), .B2(new_n639), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n703), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n771), .A2(new_n683), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n742), .A2(new_n745), .ZN(new_n773));
  INV_X1    g587(.A(new_n411), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n617), .ZN(new_n775));
  XOR2_X1   g589(.A(new_n775), .B(KEYINPUT43), .Z(new_n776));
  NAND3_X1  g590(.A1(new_n776), .A2(new_n633), .A3(new_n694), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT44), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n772), .A2(new_n773), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G137), .ZN(G39));
  NAND2_X1  g594(.A1(new_n769), .A2(new_n770), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT47), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n781), .A2(new_n302), .A3(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n782), .A2(KEYINPUT47), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n785), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n771), .A2(new_n783), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n773), .A2(new_n591), .A3(new_n618), .A4(new_n676), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n790), .B1(new_n554), .B2(new_n594), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  NAND2_X1  g607(.A1(new_n399), .A2(KEYINPUT114), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n396), .A2(new_n795), .A3(new_n398), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n411), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n618), .A2(new_n797), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n798), .A2(new_n408), .A3(new_n474), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n641), .A2(new_n799), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n668), .B(new_n800), .C1(new_n481), .C2(new_n595), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AND4_X1   g616(.A1(new_n354), .A2(new_n794), .A3(new_n676), .A4(new_n796), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n648), .B(new_n803), .C1(new_n664), .C2(new_n665), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n640), .A2(new_n804), .A3(new_n303), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n554), .A2(new_n805), .A3(new_n594), .A4(new_n773), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n747), .A2(new_n735), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n806), .B(new_n807), .C1(new_n748), .C2(new_n677), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n802), .A2(new_n758), .A3(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n588), .A2(new_n302), .A3(new_n662), .A4(new_n676), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT115), .B1(new_n744), .B2(new_n812), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n744), .A2(KEYINPUT115), .A3(new_n812), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n691), .B(new_n723), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n680), .A2(new_n701), .A3(new_n815), .A4(new_n736), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n816), .B(new_n817), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n718), .B(new_n733), .C1(new_n710), .C2(new_n628), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n715), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n810), .A2(KEYINPUT53), .A3(new_n818), .A4(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n801), .A2(new_n808), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n823), .A2(new_n820), .A3(new_n758), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n816), .B(KEYINPUT52), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n822), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n821), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT116), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n821), .A2(new_n826), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT54), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n830), .A2(KEYINPUT116), .A3(KEYINPUT54), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n707), .A2(new_n708), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n303), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n786), .A2(new_n788), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n730), .A2(new_n732), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n776), .A2(new_n673), .ZN(new_n838));
  INV_X1    g652(.A(new_n773), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n773), .A2(new_n302), .A3(new_n834), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n688), .A2(new_n592), .A3(new_n690), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n842), .A2(new_n407), .A3(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n844), .A2(new_n774), .A3(new_n614), .A4(new_n616), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n838), .A2(new_n842), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(new_n694), .A3(new_n729), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n837), .A2(new_n838), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n693), .A2(new_n709), .A3(new_n416), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT117), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n849), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT50), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI211_X1 g670(.A(KEYINPUT50), .B(new_n849), .C1(new_n852), .C2(new_n853), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n848), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n841), .A2(new_n858), .A3(KEYINPUT51), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT51), .B1(new_n841), .B2(new_n858), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n846), .A2(new_n754), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT48), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n844), .A2(new_n618), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n849), .A2(new_n646), .A3(new_n709), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n862), .A2(new_n405), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n859), .A2(new_n860), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n832), .A2(new_n833), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(KEYINPUT118), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT118), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n832), .A2(new_n866), .A3(new_n869), .A4(new_n833), .ZN(new_n870));
  OR2_X1    g684(.A1(G952), .A2(G953), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n868), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n834), .B(KEYINPUT49), .ZN(new_n873));
  INV_X1    g687(.A(new_n843), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n775), .A2(new_n303), .A3(new_n416), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n873), .A2(new_n693), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n872), .A2(new_n876), .ZN(G75));
  NOR2_X1   g691(.A1(new_n309), .A2(G952), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n830), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n880), .A2(new_n188), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT56), .B1(new_n881), .B2(G210), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n441), .A2(new_n443), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(new_n449), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT55), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n879), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n882), .B2(new_n885), .ZN(G51));
  AOI211_X1 g701(.A(KEYINPUT119), .B(new_n827), .C1(new_n821), .C2(new_n826), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n828), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n888), .B1(new_n831), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(G469), .A2(G902), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT57), .ZN(new_n893));
  OAI22_X1  g707(.A1(new_n891), .A2(new_n893), .B1(new_n273), .B2(new_n283), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n881), .A2(new_n766), .A3(new_n767), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n878), .B1(new_n894), .B2(new_n895), .ZN(G54));
  NAND3_X1  g710(.A1(new_n881), .A2(KEYINPUT58), .A3(G475), .ZN(new_n897));
  INV_X1    g711(.A(new_n363), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n897), .A2(new_n898), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n899), .A2(new_n900), .A3(new_n878), .ZN(G60));
  OR2_X1    g715(.A1(new_n610), .A2(new_n613), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n902), .A2(new_n599), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n832), .A2(new_n833), .ZN(new_n904));
  NAND2_X1  g718(.A1(G478), .A2(G902), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT59), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n903), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n903), .A2(new_n906), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n879), .B1(new_n891), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n907), .A2(new_n909), .ZN(G63));
  NAND2_X1  g724(.A1(G217), .A2(G902), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT60), .Z(new_n912));
  NAND2_X1  g726(.A1(new_n830), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n580), .A2(new_n581), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n878), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT120), .ZN(new_n916));
  INV_X1    g730(.A(new_n913), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n916), .B1(new_n917), .B2(new_n661), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n913), .A2(KEYINPUT120), .A3(new_n660), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n915), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI211_X1 g736(.A(KEYINPUT61), .B(new_n915), .C1(new_n918), .C2(new_n919), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(G66));
  INV_X1    g738(.A(G224), .ZN(new_n925));
  OAI21_X1  g739(.A(G953), .B1(new_n401), .B2(new_n925), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT121), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n801), .A2(new_n819), .A3(new_n715), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n927), .B1(new_n928), .B2(G953), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n883), .B1(G898), .B2(new_n309), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT122), .Z(new_n931));
  XNOR2_X1  g745(.A(new_n929), .B(new_n931), .ZN(G69));
  NOR2_X1   g746(.A1(new_n357), .A2(new_n358), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n530), .B(new_n933), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT123), .ZN(new_n935));
  OR4_X1    g749(.A1(new_n595), .A2(new_n684), .A3(new_n839), .A4(new_n798), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n792), .A2(new_n779), .A3(new_n936), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n680), .A2(new_n701), .A3(new_n736), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n697), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT62), .Z(new_n940));
  NAND2_X1  g754(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n935), .B1(new_n941), .B2(new_n309), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n792), .A2(new_n758), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n772), .A2(new_n723), .A3(new_n754), .ZN(new_n944));
  INV_X1    g758(.A(new_n760), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n779), .A2(new_n944), .A3(new_n945), .A4(new_n938), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n309), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n674), .A2(G953), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT125), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n934), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n942), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(G953), .B1(new_n190), .B2(new_n674), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT124), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n951), .B(new_n953), .Z(G72));
  NAND2_X1  g768(.A1(new_n534), .A2(new_n494), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT126), .Z(new_n956));
  NAND3_X1  g770(.A1(new_n937), .A2(new_n928), .A3(new_n940), .ZN(new_n957));
  NAND2_X1  g771(.A1(G472), .A2(G902), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT63), .Z(new_n959));
  AOI211_X1 g773(.A(new_n514), .B(new_n956), .C1(new_n957), .C2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n959), .ZN(new_n961));
  INV_X1    g775(.A(new_n535), .ZN(new_n962));
  AOI211_X1 g776(.A(new_n961), .B(new_n880), .C1(new_n962), .C2(new_n541), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n943), .A2(new_n946), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n961), .B1(new_n964), .B2(new_n928), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n956), .A2(new_n514), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n879), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT127), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI211_X1 g783(.A(KEYINPUT127), .B(new_n879), .C1(new_n965), .C2(new_n966), .ZN(new_n970));
  AOI211_X1 g784(.A(new_n960), .B(new_n963), .C1(new_n969), .C2(new_n970), .ZN(G57));
endmodule


