//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 1 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1292, new_n1293, new_n1295, new_n1296, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1361, new_n1362, new_n1363, new_n1364;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT64), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(new_n206), .ZN(new_n213));
  NAND2_X1  g0013(.A1(KEYINPUT64), .A2(G20), .ZN(new_n214));
  AND2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n208), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n211), .B(new_n220), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT65), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT66), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT67), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G58), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  INV_X1    g0047(.A(G13), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n248), .A2(G1), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G20), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n216), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n205), .A2(G20), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI22_X1  g0059(.A1(new_n255), .A2(new_n259), .B1(new_n250), .B2(new_n257), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OR2_X1    g0061(.A1(G223), .A2(G1698), .ZN(new_n262));
  INV_X1    g0062(.A(G1698), .ZN(new_n263));
  AND2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  OAI221_X1 g0065(.A(new_n262), .B1(G226), .B2(new_n263), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G87), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n216), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  INV_X1    g0072(.A(G41), .ZN(new_n273));
  INV_X1    g0073(.A(G45), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n271), .A2(new_n272), .B1(new_n275), .B2(new_n205), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT68), .B(G45), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n273), .ZN(new_n278));
  INV_X1    g0078(.A(G274), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(G1), .ZN(new_n280));
  AOI22_X1  g0080(.A1(G232), .A2(new_n276), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G190), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n270), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G200), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n278), .A2(new_n280), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n271), .A2(new_n272), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n275), .A2(new_n205), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(new_n287), .A3(G232), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n286), .B1(new_n266), .B2(new_n267), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n284), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n283), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT76), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT3), .ZN(new_n294));
  INV_X1    g0094(.A(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(KEYINPUT3), .A2(G33), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n213), .A2(new_n296), .A3(new_n214), .A4(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT7), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n293), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n264), .A2(new_n265), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n215), .A2(KEYINPUT76), .A3(KEYINPUT7), .A4(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT75), .ZN(new_n304));
  NOR3_X1   g0104(.A1(new_n264), .A2(new_n265), .A3(G20), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n304), .B1(new_n305), .B2(KEYINPUT7), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n296), .A2(new_n297), .ZN(new_n307));
  OAI211_X1 g0107(.A(KEYINPUT75), .B(new_n299), .C1(new_n307), .C2(G20), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n303), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G68), .ZN(new_n311));
  AND2_X1   g0111(.A1(G58), .A2(G68), .ZN(new_n312));
  NOR2_X1   g0112(.A1(G58), .A2(G68), .ZN(new_n313));
  OAI211_X1 g0113(.A(KEYINPUT73), .B(G20), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(G20), .A2(G33), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G159), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g0117(.A(G58), .B(G68), .ZN(new_n318));
  AOI21_X1  g0118(.A(KEYINPUT73), .B1(new_n318), .B2(G20), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(KEYINPUT16), .B1(new_n311), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT74), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(new_n317), .B2(new_n319), .ZN(new_n323));
  OAI21_X1  g0123(.A(G20), .B1(new_n312), .B2(new_n313), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT73), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n326), .A2(KEYINPUT74), .A3(new_n316), .A4(new_n314), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G68), .ZN(new_n329));
  AND4_X1   g0129(.A1(new_n213), .A2(new_n296), .A3(new_n214), .A4(new_n297), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n329), .B1(new_n330), .B2(new_n299), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT7), .B1(new_n307), .B2(G20), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n328), .A2(KEYINPUT16), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n253), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n261), .B(new_n292), .C1(new_n321), .C2(new_n335), .ZN(new_n336));
  XNOR2_X1  g0136(.A(KEYINPUT77), .B(KEYINPUT17), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT77), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(KEYINPUT17), .ZN(new_n340));
  INV_X1    g0140(.A(new_n253), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n323), .A2(new_n327), .B1(new_n331), .B2(new_n332), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n341), .B1(new_n342), .B2(KEYINPUT16), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT16), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n329), .B1(new_n303), .B2(new_n309), .ZN(new_n345));
  INV_X1    g0145(.A(new_n320), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n260), .B1(new_n343), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n340), .B1(new_n348), .B2(new_n292), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n338), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n261), .B1(new_n321), .B2(new_n335), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT18), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n270), .A2(new_n281), .A3(G179), .ZN(new_n353));
  OAI21_X1  g0153(.A(G169), .B1(new_n289), .B2(new_n290), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n351), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n355), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT18), .B1(new_n348), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n350), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n263), .B1(new_n296), .B2(new_n297), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n361), .A2(G223), .B1(new_n301), .B2(G77), .ZN(new_n362));
  INV_X1    g0162(.A(G222), .ZN(new_n363));
  AOI21_X1  g0163(.A(G1698), .B1(new_n296), .B2(new_n297), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n362), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n269), .ZN(new_n367));
  INV_X1    g0167(.A(new_n285), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(G226), .B2(new_n276), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G169), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n315), .A2(G150), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n215), .A2(G33), .ZN(new_n374));
  OAI221_X1 g0174(.A(new_n373), .B1(new_n206), .B2(new_n201), .C1(new_n374), .C2(new_n256), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n253), .ZN(new_n376));
  INV_X1    g0176(.A(G50), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n377), .B1(new_n205), .B2(G20), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n254), .A2(new_n378), .B1(new_n377), .B2(new_n251), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n372), .B(new_n380), .C1(G179), .C2(new_n370), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n276), .A2(G244), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n361), .A2(G238), .B1(new_n301), .B2(G107), .ZN(new_n383));
  INV_X1    g0183(.A(G232), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n383), .B1(new_n384), .B2(new_n365), .ZN(new_n385));
  AOI211_X1 g0185(.A(new_n368), .B(new_n382), .C1(new_n385), .C2(new_n269), .ZN(new_n386));
  INV_X1    g0186(.A(G179), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n213), .A2(new_n214), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n257), .A2(new_n315), .B1(new_n389), .B2(G77), .ZN(new_n390));
  XNOR2_X1  g0190(.A(KEYINPUT15), .B(G87), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n390), .B1(new_n374), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n253), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n258), .A2(G77), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n254), .A2(new_n395), .B1(new_n202), .B2(new_n251), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n388), .B(new_n397), .C1(G169), .C2(new_n386), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n386), .A2(G190), .ZN(new_n399));
  INV_X1    g0199(.A(new_n397), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n399), .B(new_n400), .C1(new_n284), .C2(new_n386), .ZN(new_n401));
  AND2_X1   g0201(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n380), .A2(KEYINPUT9), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT9), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n376), .A2(new_n404), .A3(new_n379), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n403), .A2(new_n405), .B1(G200), .B2(new_n370), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT10), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT69), .ZN(new_n408));
  INV_X1    g0208(.A(new_n370), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n408), .B1(new_n409), .B2(G190), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n406), .A2(new_n407), .A3(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n407), .B1(new_n406), .B2(new_n410), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n381), .B(new_n402), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT70), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n413), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n411), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n418), .A2(KEYINPUT70), .A3(new_n381), .A4(new_n402), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n384), .A2(G1698), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n307), .B(new_n420), .C1(G226), .C2(G1698), .ZN(new_n421));
  NAND2_X1  g0221(.A1(G33), .A2(G97), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n286), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n276), .A2(G238), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n285), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT71), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT13), .ZN(new_n427));
  OAI22_X1  g0227(.A1(new_n423), .A2(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n423), .ZN(new_n429));
  INV_X1    g0229(.A(new_n425), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(new_n430), .A3(KEYINPUT13), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n428), .B1(new_n431), .B2(new_n426), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(G179), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n427), .B1(new_n423), .B2(new_n425), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n431), .A2(G169), .A3(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT14), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n436), .A2(KEYINPUT72), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n435), .A2(new_n437), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n315), .A2(G50), .B1(G20), .B2(new_n329), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n374), .B2(new_n202), .ZN(new_n442));
  AOI21_X1  g0242(.A(KEYINPUT11), .B1(new_n442), .B2(new_n253), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(KEYINPUT11), .A3(new_n253), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n258), .A2(G68), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT12), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n446), .B1(new_n251), .B2(new_n329), .ZN(new_n447));
  NOR3_X1   g0247(.A1(new_n250), .A2(KEYINPUT12), .A3(G68), .ZN(new_n448));
  OAI221_X1 g0248(.A(new_n444), .B1(new_n255), .B2(new_n445), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  OAI22_X1  g0249(.A1(new_n439), .A2(new_n440), .B1(new_n443), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n449), .A2(new_n443), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n432), .A2(G190), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n431), .A2(G200), .A3(new_n434), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  AND4_X1   g0255(.A1(new_n360), .A2(new_n416), .A3(new_n419), .A4(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT80), .ZN(new_n458));
  NOR3_X1   g0258(.A1(new_n202), .A2(G20), .A3(G33), .ZN(new_n459));
  OR2_X1    g0259(.A1(new_n459), .A2(KEYINPUT78), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(KEYINPUT78), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g0262(.A(G97), .B(G107), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT6), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G97), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n464), .A2(new_n466), .A3(G107), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n462), .B1(new_n468), .B2(new_n215), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n310), .A2(G107), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n469), .B1(new_n470), .B2(KEYINPUT79), .ZN(new_n471));
  INV_X1    g0271(.A(G107), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n472), .B1(new_n303), .B2(new_n309), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT79), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n341), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n250), .A2(G97), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n205), .A2(G33), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n341), .A2(new_n250), .A3(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n477), .B1(new_n480), .B2(G97), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n458), .B1(new_n476), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n475), .ZN(new_n484));
  OR2_X1    g0284(.A1(new_n465), .A2(new_n467), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n485), .A2(new_n389), .B1(new_n460), .B2(new_n461), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(new_n473), .B2(new_n474), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n253), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(KEYINPUT80), .A3(new_n481), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n307), .A2(G244), .A3(new_n263), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT4), .ZN(new_n491));
  OAI21_X1  g0291(.A(KEYINPUT82), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT82), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n364), .A2(new_n493), .A3(KEYINPUT4), .A4(G244), .ZN(new_n494));
  XNOR2_X1  g0294(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n361), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n492), .A2(new_n494), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n269), .ZN(new_n499));
  XNOR2_X1  g0299(.A(KEYINPUT5), .B(G41), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n274), .A2(G1), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n502), .A2(G257), .A3(new_n286), .ZN(new_n503));
  NOR3_X1   g0303(.A1(new_n274), .A2(new_n279), .A3(G1), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n286), .A2(new_n500), .A3(new_n504), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n503), .A2(KEYINPUT83), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT83), .B1(new_n503), .B2(new_n505), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n499), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n503), .A2(new_n505), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n510), .B1(new_n498), .B2(new_n269), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n509), .A2(G200), .B1(G190), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n483), .A2(new_n489), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n488), .A2(new_n481), .ZN(new_n514));
  INV_X1    g0314(.A(new_n509), .ZN(new_n515));
  INV_X1    g0315(.A(new_n510), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n499), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n515), .A2(new_n387), .B1(new_n371), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n391), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n520), .A2(new_n250), .ZN(new_n521));
  INV_X1    g0321(.A(G87), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n479), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(new_n466), .A3(new_n472), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT19), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n422), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n524), .B1(new_n389), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n213), .A2(G33), .A3(G97), .A4(new_n214), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n525), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n213), .B(new_n214), .C1(new_n264), .C2(new_n265), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n527), .B(new_n529), .C1(new_n329), .C2(new_n530), .ZN(new_n531));
  AOI211_X1 g0331(.A(new_n521), .B(new_n523), .C1(new_n531), .C2(new_n253), .ZN(new_n532));
  INV_X1    g0332(.A(new_n504), .ZN(new_n533));
  OAI21_X1  g0333(.A(G250), .B1(new_n274), .B2(G1), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n269), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI211_X1 g0335(.A(G238), .B(new_n263), .C1(new_n264), .C2(new_n265), .ZN(new_n536));
  OAI211_X1 g0336(.A(G244), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n537));
  INV_X1    g0337(.A(G116), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n536), .B(new_n537), .C1(new_n295), .C2(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n535), .B1(new_n539), .B2(new_n269), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G190), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n532), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n539), .A2(new_n269), .ZN(new_n543));
  INV_X1    g0343(.A(new_n535), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G200), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n371), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n540), .A2(new_n387), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n521), .B1(new_n531), .B2(new_n253), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n480), .A2(new_n520), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n542), .A2(new_n546), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n513), .A2(new_n519), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n295), .A2(G97), .ZN(new_n555));
  NAND2_X1  g0355(.A1(G33), .A2(G283), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n213), .A2(new_n555), .A3(new_n214), .A4(new_n556), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n252), .A2(new_n216), .B1(G20), .B2(new_n538), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(KEYINPUT84), .A2(KEYINPUT20), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(KEYINPUT84), .A2(KEYINPUT20), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n559), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n557), .A2(new_n558), .A3(new_n560), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n251), .A2(new_n538), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n479), .B2(new_n538), .ZN(new_n567));
  OR2_X1    g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n502), .A2(G270), .A3(new_n286), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n569), .A2(new_n505), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n307), .A2(G264), .A3(G1698), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n307), .A2(G257), .A3(new_n263), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n301), .A2(G303), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n269), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n568), .A2(G169), .A3(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT21), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n568), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n569), .A2(new_n505), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n269), .B2(new_n574), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(G190), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n580), .B(new_n583), .C1(new_n284), .C2(new_n582), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n576), .A2(new_n387), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n568), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n568), .A2(KEYINPUT21), .A3(G169), .A4(new_n576), .ZN(new_n587));
  AND4_X1   g0387(.A1(new_n579), .A2(new_n584), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(KEYINPUT22), .B1(new_n530), .B2(new_n522), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT22), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n215), .A2(new_n590), .A3(G87), .A4(new_n307), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(KEYINPUT23), .A2(G107), .ZN(new_n593));
  AOI21_X1  g0393(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n593), .B1(new_n594), .B2(G20), .ZN(new_n595));
  NOR2_X1   g0395(.A1(KEYINPUT23), .A2(G107), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n595), .B1(new_n389), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g0398(.A(KEYINPUT85), .B(KEYINPUT24), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n599), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n592), .A2(new_n597), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n341), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n251), .A2(KEYINPUT25), .A3(new_n472), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT25), .B1(new_n251), .B2(new_n472), .ZN(new_n606));
  OAI22_X1  g0406(.A1(new_n605), .A2(new_n606), .B1(new_n479), .B2(new_n472), .ZN(new_n607));
  OAI21_X1  g0407(.A(KEYINPUT86), .B1(new_n603), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n602), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n601), .B1(new_n592), .B2(new_n597), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n253), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT86), .ZN(new_n612));
  INV_X1    g0412(.A(new_n607), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n502), .A2(G264), .A3(new_n286), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT87), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n269), .B1(new_n501), .B2(new_n500), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n618), .A2(KEYINPUT87), .A3(G264), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n307), .A2(G257), .A3(G1698), .ZN(new_n621));
  NAND2_X1  g0421(.A1(G33), .A2(G294), .ZN(new_n622));
  OAI211_X1 g0422(.A(G250), .B(new_n263), .C1(new_n264), .C2(new_n265), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n269), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n620), .A2(new_n505), .A3(new_n625), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n625), .A2(new_n505), .A3(new_n615), .ZN(new_n627));
  OAI22_X1  g0427(.A1(new_n626), .A2(new_n387), .B1(new_n627), .B2(new_n371), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n608), .A2(new_n614), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n611), .A2(new_n613), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n284), .A2(new_n626), .B1(new_n627), .B2(new_n282), .ZN(new_n631));
  OR2_X1    g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n588), .A2(new_n629), .A3(new_n632), .ZN(new_n633));
  NOR3_X1   g0433(.A1(new_n457), .A2(new_n554), .A3(new_n633), .ZN(G372));
  NOR2_X1   g0434(.A1(new_n630), .A2(new_n631), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n545), .A2(KEYINPUT88), .A3(G200), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT88), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n637), .B1(new_n540), .B2(new_n284), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n532), .A2(new_n636), .A3(new_n541), .A4(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n552), .A2(new_n547), .A3(new_n548), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT89), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n639), .A2(new_n640), .A3(KEYINPUT89), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n635), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n579), .A2(new_n586), .A3(new_n587), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n630), .A2(new_n628), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n513), .A2(new_n645), .A3(new_n648), .A4(new_n519), .ZN(new_n649));
  INV_X1    g0449(.A(new_n640), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n553), .A2(new_n514), .A3(new_n518), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n650), .B1(new_n651), .B2(KEYINPUT26), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n483), .A2(new_n489), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n643), .A2(new_n644), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n653), .A2(new_n654), .A3(new_n518), .A4(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n649), .A2(new_n652), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n456), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n398), .A2(KEYINPUT90), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n386), .A2(G169), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT90), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n660), .A2(new_n661), .A3(new_n388), .A4(new_n397), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n659), .A2(new_n454), .A3(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n350), .B1(new_n663), .B2(new_n450), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n418), .B1(new_n664), .B2(new_n359), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n665), .A2(new_n381), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n658), .A2(new_n666), .ZN(G369));
  INV_X1    g0467(.A(G330), .ZN(new_n668));
  INV_X1    g0468(.A(new_n646), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n215), .A2(new_n249), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n669), .A2(new_n568), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n675), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n588), .B1(new_n580), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n679), .A2(KEYINPUT91), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(KEYINPUT91), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n668), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT92), .ZN(new_n683));
  INV_X1    g0483(.A(new_n629), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n675), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n608), .A2(new_n614), .A3(new_n675), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n629), .A2(new_n632), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n683), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n685), .A2(new_n683), .A3(new_n687), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n682), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n646), .A2(new_n675), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n685), .A2(new_n683), .A3(new_n687), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n693), .B1(new_n694), .B2(new_n688), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n630), .A2(new_n628), .A3(new_n677), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n692), .A2(new_n697), .ZN(G399));
  INV_X1    g0498(.A(new_n209), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(G41), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n524), .A2(G116), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(G1), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n218), .B2(new_n701), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT28), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n653), .A2(new_n518), .A3(new_n655), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(KEYINPUT26), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n646), .A2(new_n629), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n513), .A2(new_n645), .A3(new_n708), .A4(new_n519), .ZN(new_n709));
  INV_X1    g0509(.A(new_n651), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n650), .B1(new_n710), .B2(new_n654), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n707), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n712), .A2(KEYINPUT29), .A3(new_n677), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n657), .A2(new_n677), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n713), .B1(new_n714), .B2(KEYINPUT29), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT30), .ZN(new_n716));
  AOI22_X1  g0516(.A1(new_n617), .A2(new_n619), .B1(new_n269), .B2(new_n624), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n582), .A2(new_n717), .A3(G179), .A4(new_n540), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n716), .B1(new_n718), .B2(new_n517), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n717), .A2(new_n540), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n720), .A2(KEYINPUT30), .A3(new_n585), .A4(new_n511), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n540), .A2(G179), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n509), .A2(new_n626), .A3(new_n576), .A4(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n719), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n724), .A2(KEYINPUT31), .A3(new_n675), .ZN(new_n725));
  AOI21_X1  g0525(.A(KEYINPUT31), .B1(new_n724), .B2(new_n675), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n588), .A2(new_n629), .A3(new_n632), .A4(new_n677), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n727), .B1(new_n554), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G330), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT93), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n729), .A2(KEYINPUT93), .A3(G330), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n715), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n705), .B1(new_n736), .B2(G1), .ZN(G364));
  INV_X1    g0537(.A(new_n682), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n389), .A2(new_n248), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G45), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G1), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n700), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n680), .A2(new_n668), .A3(new_n681), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n738), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n248), .A2(new_n295), .A3(KEYINPUT95), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT95), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(G13), .B2(G33), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n216), .B1(G20), .B2(new_n371), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n699), .A2(new_n307), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n246), .A2(new_n274), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n756), .B(new_n757), .C1(new_n219), .C2(new_n277), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT94), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n209), .A2(new_n307), .ZN(new_n760));
  INV_X1    g0560(.A(G355), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n760), .A2(new_n761), .B1(G116), .B2(new_n209), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n758), .B1(new_n759), .B2(new_n762), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n762), .A2(new_n759), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n754), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n284), .A2(G179), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n766), .A2(G20), .A3(G190), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n307), .B1(new_n768), .B2(G303), .ZN(new_n769));
  INV_X1    g0569(.A(G329), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G179), .A2(G200), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n389), .A2(new_n282), .A3(new_n771), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n769), .A2(KEYINPUT100), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n389), .A2(new_n282), .A3(new_n766), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n771), .A2(G190), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n389), .A2(new_n776), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n775), .A2(G283), .B1(G294), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n215), .A2(new_n387), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G190), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  XOR2_X1   g0582(.A(KEYINPUT33), .B(G317), .Z(new_n783));
  OAI21_X1  g0583(.A(new_n778), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n773), .B(new_n784), .C1(KEYINPUT100), .C2(new_n769), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n779), .A2(KEYINPUT96), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G200), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n779), .A2(KEYINPUT96), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n282), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT98), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(new_n780), .B2(new_n282), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n779), .A2(KEYINPUT98), .A3(G190), .A4(G200), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n790), .A2(G322), .B1(G326), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G311), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n787), .A2(new_n282), .A3(new_n788), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n785), .B(new_n795), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n790), .B(KEYINPUT97), .Z(new_n799));
  INV_X1    g0599(.A(G58), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n777), .A2(G97), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n782), .B2(new_n329), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT99), .ZN(new_n804));
  INV_X1    g0604(.A(new_n797), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G77), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n794), .A2(G50), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n775), .A2(G107), .ZN(new_n808));
  INV_X1    g0608(.A(G159), .ZN(new_n809));
  OAI21_X1  g0609(.A(KEYINPUT32), .B1(new_n772), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n301), .B1(new_n768), .B2(G87), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n808), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NOR3_X1   g0612(.A1(new_n772), .A2(KEYINPUT32), .A3(new_n809), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n804), .A2(new_n806), .A3(new_n807), .A4(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n798), .B1(new_n801), .B2(new_n815), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n765), .B(new_n743), .C1(new_n816), .C2(new_n752), .ZN(new_n817));
  INV_X1    g0617(.A(new_n751), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n679), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n745), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(G396));
  NAND4_X1  g0621(.A1(new_n659), .A2(new_n397), .A3(new_n662), .A4(new_n675), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n398), .B(new_n401), .C1(new_n400), .C2(new_n677), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n714), .B(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n742), .B1(new_n826), .B2(new_n734), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n734), .B2(new_n826), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n749), .A2(new_n752), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n743), .B1(new_n202), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n775), .A2(G87), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n307), .B1(new_n768), .B2(G107), .ZN(new_n832));
  AND3_X1   g0632(.A1(new_n831), .A2(new_n802), .A3(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(G283), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n833), .B1(new_n796), .B2(new_n772), .C1(new_n782), .C2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n790), .ZN(new_n836));
  INV_X1    g0636(.A(G294), .ZN(new_n837));
  INV_X1    g0637(.A(G303), .ZN(new_n838));
  INV_X1    g0638(.A(new_n794), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n836), .A2(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n835), .B(new_n840), .C1(G116), .C2(new_n805), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n794), .A2(G137), .B1(G150), .B2(new_n781), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n809), .B2(new_n797), .ZN(new_n843));
  INV_X1    g0643(.A(new_n799), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n843), .B1(new_n844), .B2(G143), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(KEYINPUT34), .Z(new_n846));
  NAND2_X1  g0646(.A1(new_n775), .A2(G68), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n301), .B1(new_n768), .B2(G50), .ZN(new_n848));
  INV_X1    g0648(.A(new_n777), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n847), .B(new_n848), .C1(new_n800), .C2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n772), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n850), .B1(G132), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n841), .B1(new_n846), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n752), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n830), .B1(new_n750), .B2(new_n825), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n828), .A2(new_n855), .ZN(G384));
  NOR2_X1   g0656(.A1(new_n739), .A2(new_n205), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n358), .B(new_n356), .C1(new_n338), .C2(new_n349), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n328), .A2(new_n333), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n344), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n260), .B1(new_n343), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT101), .B1(new_n861), .B2(new_n673), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n342), .A2(KEYINPUT16), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n261), .B1(new_n335), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT101), .ZN(new_n865));
  INV_X1    g0665(.A(new_n673), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n858), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n864), .A2(new_n355), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT102), .B1(new_n871), .B2(new_n336), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n872), .A2(new_n868), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n871), .A2(KEYINPUT102), .A3(new_n336), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n870), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n351), .A2(new_n355), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n673), .B(KEYINPUT103), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n351), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n876), .A2(new_n879), .A3(new_n870), .A4(new_n336), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  OAI211_X1 g0681(.A(KEYINPUT38), .B(new_n869), .C1(new_n875), .C2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n348), .A2(new_n877), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n336), .B1(new_n348), .B2(new_n357), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT37), .B1(new_n884), .B2(new_n883), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n858), .A2(new_n883), .B1(new_n885), .B2(new_n880), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT104), .B1(new_n886), .B2(KEYINPUT38), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n858), .A2(new_n883), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n885), .A2(new_n880), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT104), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n882), .A2(new_n887), .A3(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT39), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n450), .A2(new_n675), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n862), .A2(new_n867), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT102), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n283), .A2(new_n291), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n260), .B(new_n900), .C1(new_n347), .C2(new_n343), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n343), .A2(new_n860), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n357), .B1(new_n902), .B2(new_n261), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n899), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n898), .A2(new_n874), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n881), .B1(new_n905), .B2(KEYINPUT37), .ZN(new_n906));
  INV_X1    g0706(.A(new_n869), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n892), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(new_n882), .A3(KEYINPUT39), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n896), .A2(new_n897), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n450), .A2(new_n454), .ZN(new_n911));
  INV_X1    g0711(.A(new_n451), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n911), .A2(new_n912), .A3(new_n675), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n450), .B(new_n454), .C1(new_n451), .C2(new_n677), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n657), .A2(new_n677), .A3(new_n825), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n398), .A2(new_n675), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n916), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n908), .A2(new_n882), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n920), .A2(new_n921), .B1(new_n359), .B2(new_n877), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n910), .A2(new_n922), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n456), .B(new_n713), .C1(new_n714), .C2(KEYINPUT29), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n666), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n923), .B(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n824), .B1(new_n914), .B2(new_n913), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n927), .A2(KEYINPUT40), .A3(new_n729), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n894), .A2(new_n928), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n927), .A2(new_n729), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT40), .B1(new_n921), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n456), .A2(new_n729), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n668), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n933), .B2(new_n932), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n857), .B1(new_n926), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n926), .B2(new_n935), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n485), .A2(KEYINPUT35), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n485), .A2(KEYINPUT35), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n938), .A2(G116), .A3(new_n217), .A4(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT36), .ZN(new_n941));
  NOR3_X1   g0741(.A1(new_n218), .A2(new_n312), .A3(new_n202), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n329), .A2(G50), .ZN(new_n943));
  OAI211_X1 g0743(.A(G1), .B(new_n248), .C1(new_n942), .C2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n937), .A2(new_n941), .A3(new_n944), .ZN(G367));
  NOR2_X1   g0745(.A1(new_n677), .A2(new_n532), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n643), .B2(new_n644), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(new_n650), .B2(new_n946), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n751), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n754), .B1(new_n699), .B2(new_n520), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n755), .A2(new_n238), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n743), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n805), .A2(G50), .B1(G143), .B2(new_n794), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n775), .A2(G77), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n851), .A2(G137), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n777), .A2(G68), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n301), .B1(new_n768), .B2(G58), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n954), .A2(new_n955), .A3(new_n956), .A4(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(G159), .B2(new_n781), .ZN(new_n959));
  INV_X1    g0759(.A(G150), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n953), .B(new_n959), .C1(new_n960), .C2(new_n836), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT113), .Z(new_n962));
  NAND2_X1  g0762(.A1(new_n844), .A2(G303), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT46), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n767), .B2(new_n538), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n768), .A2(KEYINPUT46), .A3(G116), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n965), .B(new_n966), .C1(new_n782), .C2(new_n837), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n967), .A2(KEYINPUT111), .B1(new_n805), .B2(G283), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n796), .B2(new_n839), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n967), .A2(KEYINPUT111), .B1(new_n472), .B2(new_n849), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n775), .A2(G97), .ZN(new_n971));
  INV_X1    g0771(.A(G317), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n971), .B(new_n301), .C1(new_n972), .C2(new_n772), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT112), .Z(new_n974));
  NOR3_X1   g0774(.A1(new_n969), .A2(new_n970), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n962), .B1(new_n963), .B2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT47), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n949), .B(new_n952), .C1(new_n977), .C2(new_n854), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n741), .B(KEYINPUT110), .Z(new_n979));
  INV_X1    g0779(.A(new_n692), .ZN(new_n980));
  AND3_X1   g0780(.A1(new_n488), .A2(KEYINPUT80), .A3(new_n481), .ZN(new_n981));
  AOI21_X1  g0781(.A(KEYINPUT80), .B1(new_n488), .B2(new_n481), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n675), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n983), .A2(new_n513), .A3(new_n519), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(KEYINPUT105), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT105), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n983), .A2(new_n986), .A3(new_n513), .A4(new_n519), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n518), .B(new_n675), .C1(new_n981), .C2(new_n982), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n985), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(KEYINPUT106), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n695), .A2(new_n696), .ZN(new_n991));
  INV_X1    g0791(.A(new_n988), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(new_n984), .B2(KEYINPUT105), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT106), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n993), .A2(new_n994), .A3(new_n987), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n990), .A2(new_n991), .A3(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT44), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n990), .A2(KEYINPUT44), .A3(new_n991), .A4(new_n995), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AND3_X1   g0800(.A1(new_n993), .A2(new_n994), .A3(new_n987), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n994), .B1(new_n993), .B2(new_n987), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n697), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n990), .A2(new_n995), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1007), .A2(new_n697), .A3(new_n1004), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  OAI211_X1 g0809(.A(KEYINPUT109), .B(new_n980), .C1(new_n1000), .C2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n695), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n691), .A2(new_n693), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n738), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1012), .A2(new_n1011), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n682), .ZN(new_n1015));
  AND2_X1   g0815(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1016), .A2(new_n736), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n998), .A2(new_n999), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1018), .A2(new_n692), .A3(new_n1008), .A4(new_n1006), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1010), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1018), .A2(new_n1008), .A3(new_n1006), .ZN(new_n1021));
  AOI21_X1  g0821(.A(KEYINPUT109), .B1(new_n1021), .B2(new_n980), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n736), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n700), .B(KEYINPUT41), .Z(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n979), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT43), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n948), .A2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n948), .A2(new_n1027), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT107), .ZN(new_n1031));
  NOR3_X1   g0831(.A1(new_n1001), .A2(new_n1002), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(KEYINPUT107), .B1(new_n990), .B2(new_n995), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n684), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n675), .B1(new_n1034), .B2(new_n519), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n695), .B1(new_n990), .B2(new_n995), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT42), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1036), .B(new_n1037), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1028), .B(new_n1030), .C1(new_n1035), .C2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1007), .A2(new_n1031), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n990), .A2(KEYINPUT107), .A3(new_n995), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n629), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n519), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n677), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1036), .B(KEYINPUT42), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1044), .A2(new_n1027), .A3(new_n948), .A4(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1039), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n980), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1049), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1039), .A2(new_n1046), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n978), .B1(new_n1026), .B2(new_n1053), .ZN(G387));
  NAND2_X1  g0854(.A1(new_n1016), .A2(new_n979), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT114), .Z(new_n1056));
  NAND3_X1  g0856(.A1(new_n689), .A2(new_n690), .A3(new_n751), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n760), .A2(new_n702), .B1(G107), .B2(new_n209), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT115), .Z(new_n1059));
  INV_X1    g0859(.A(new_n277), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n234), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n702), .ZN(new_n1062));
  AOI211_X1 g0862(.A(G45), .B(new_n1062), .C1(G68), .C2(G77), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n256), .A2(G50), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT50), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n756), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1059), .B1(new_n1061), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n742), .B1(new_n1067), .B2(new_n754), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n781), .A2(new_n257), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(KEYINPUT116), .B(G150), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n851), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n307), .B1(new_n767), .B2(new_n202), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n520), .B2(new_n777), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1069), .A2(new_n971), .A3(new_n1071), .A4(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(G50), .B2(new_n790), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n839), .A2(KEYINPUT117), .A3(new_n809), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT117), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n794), .B2(G159), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1075), .B1(new_n329), .B2(new_n797), .C1(new_n1076), .C2(new_n1078), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n794), .A2(G322), .B1(G311), .B2(new_n781), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1080), .B1(new_n838), .B2(new_n797), .C1(new_n799), .C2(new_n972), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT48), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G294), .A2(new_n768), .B1(new_n777), .B2(G283), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT49), .Z(new_n1087));
  AOI21_X1  g0887(.A(new_n307), .B1(new_n851), .B2(G326), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n538), .B2(new_n774), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1079), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1068), .B1(new_n1090), .B2(new_n752), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1056), .B1(new_n1057), .B2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1017), .A2(new_n701), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n736), .B2(new_n1016), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1092), .A2(new_n1094), .ZN(G393));
  NAND2_X1  g0895(.A1(new_n1021), .A2(new_n980), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1096), .A2(new_n1019), .A3(new_n979), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n243), .A2(new_n755), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n753), .B1(new_n466), .B2(new_n209), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n742), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n307), .B1(new_n768), .B2(G283), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n808), .A2(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n781), .A2(G303), .B1(G116), .B2(new_n777), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n797), .B2(new_n837), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT120), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1102), .B(new_n1105), .C1(G322), .C2(new_n851), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n790), .A2(G311), .B1(G317), .B2(new_n794), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT119), .ZN(new_n1108));
  OR2_X1    g0908(.A1(new_n1108), .A2(KEYINPUT52), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(KEYINPUT52), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1106), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n790), .A2(G159), .B1(G150), .B2(new_n794), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT118), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1113), .A2(KEYINPUT51), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(KEYINPUT51), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n849), .A2(new_n202), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n301), .B(new_n1116), .C1(G68), .C2(new_n768), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n781), .A2(G50), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n851), .A2(G143), .ZN(new_n1119));
  AND4_X1   g0919(.A1(new_n831), .A2(new_n1117), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1115), .B(new_n1120), .C1(new_n256), .C2(new_n797), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1111), .B1(new_n1114), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1100), .B1(new_n1122), .B2(new_n752), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n1048), .B2(new_n818), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1097), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1017), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1019), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n692), .B1(new_n1129), .B2(new_n1018), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1127), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n700), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1126), .B1(new_n1132), .B2(new_n1133), .ZN(G390));
  AND2_X1   g0934(.A1(new_n896), .A2(new_n909), .ZN(new_n1135));
  OR2_X1    g0935(.A1(new_n1135), .A2(new_n750), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n829), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n742), .B1(new_n257), .B2(new_n1137), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n790), .A2(G116), .B1(G283), .B2(new_n794), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1116), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n851), .A2(G294), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n307), .B1(new_n768), .B2(G87), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1140), .A2(new_n847), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G107), .B2(new_n781), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1139), .B(new_n1144), .C1(new_n466), .C2(new_n797), .ZN(new_n1145));
  INV_X1    g0945(.A(G137), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n782), .A2(new_n1146), .B1(new_n809), .B2(new_n849), .ZN(new_n1147));
  XOR2_X1   g0947(.A(KEYINPUT54), .B(G143), .Z(new_n1148));
  AOI21_X1  g0948(.A(new_n1147), .B1(new_n805), .B2(new_n1148), .ZN(new_n1149));
  XOR2_X1   g0949(.A(new_n1149), .B(KEYINPUT123), .Z(new_n1150));
  OAI21_X1  g0950(.A(new_n307), .B1(new_n774), .B2(new_n377), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G125), .B2(new_n851), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT124), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n768), .A2(new_n1070), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT53), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(new_n794), .B2(G128), .ZN(new_n1156));
  INV_X1    g0956(.A(G132), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1153), .B(new_n1156), .C1(new_n836), .C2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1145), .B1(new_n1150), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1138), .B1(new_n1159), .B2(new_n752), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1136), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n897), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n894), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n712), .A2(new_n677), .A3(new_n825), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n916), .B1(new_n1164), .B2(new_n919), .ZN(new_n1165));
  OR2_X1    g0965(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n729), .A2(KEYINPUT93), .A3(G330), .ZN(new_n1167));
  AOI21_X1  g0967(.A(KEYINPUT93), .B1(new_n729), .B2(G330), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n1167), .A2(new_n1168), .A3(new_n824), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n915), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n920), .A2(new_n897), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1166), .B(new_n1170), .C1(new_n1135), .C2(new_n1171), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n729), .A2(G330), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n927), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n917), .A2(new_n919), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n915), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n896), .A2(new_n909), .B1(new_n1177), .B2(new_n1162), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1175), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1172), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n979), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1161), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n456), .A2(new_n1173), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n924), .A2(new_n666), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(KEYINPUT121), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT121), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n924), .A2(new_n1188), .A3(new_n666), .A4(new_n1185), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(KEYINPUT122), .B1(new_n1169), .B2(new_n915), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n732), .A2(new_n733), .A3(new_n825), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT122), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1192), .A2(new_n1193), .A3(new_n916), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1191), .A2(new_n1174), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n1176), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1164), .A2(new_n919), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n915), .B1(new_n1173), .B2(new_n825), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1197), .B(new_n1198), .C1(new_n1169), .C2(new_n915), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1190), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1172), .A2(new_n1180), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n700), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1190), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1192), .A2(new_n916), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1175), .B1(new_n1205), .B2(KEYINPUT122), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1206), .A2(new_n1194), .B1(new_n917), .B2(new_n919), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1204), .B1(new_n1207), .B2(new_n1199), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1208), .A2(new_n1181), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1184), .B1(new_n1203), .B2(new_n1209), .ZN(G378));
  NOR3_X1   g1010(.A1(new_n929), .A2(new_n931), .A3(new_n668), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n923), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n418), .A2(new_n381), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n380), .A2(new_n866), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1213), .B(new_n1214), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1215), .B(new_n1216), .Z(new_n1217));
  NAND2_X1  g1017(.A1(new_n894), .A2(new_n928), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n927), .A2(new_n729), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n882), .B2(new_n908), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1218), .B(G330), .C1(new_n1220), .C2(KEYINPUT40), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1221), .A2(new_n910), .A3(new_n922), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1212), .A2(new_n1217), .A3(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1217), .B1(new_n1212), .B2(new_n1222), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n979), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n743), .B1(new_n377), .B2(new_n829), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n790), .A2(G128), .B1(G125), .B2(new_n794), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n768), .A2(new_n1148), .B1(new_n777), .B2(G150), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n782), .B2(new_n1157), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(G137), .B2(new_n805), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1231));
  XOR2_X1   g1031(.A(new_n1231), .B(KEYINPUT125), .Z(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  OR2_X1    g1033(.A1(new_n1233), .A2(KEYINPUT59), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(KEYINPUT59), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n295), .B(new_n273), .C1(new_n774), .C2(new_n809), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(G124), .B2(new_n851), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1234), .A2(new_n1235), .A3(new_n1237), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n790), .A2(G107), .B1(G116), .B2(new_n794), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n851), .A2(G283), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n775), .A2(G58), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n301), .A2(new_n273), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(new_n768), .B2(G77), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1240), .A2(new_n1241), .A3(new_n956), .A4(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G97), .B2(new_n781), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1239), .B(new_n1245), .C1(new_n391), .C2(new_n797), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT58), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  OR2_X1    g1048(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1242), .B(new_n377), .C1(G33), .C2(G41), .ZN(new_n1250));
  AND4_X1   g1050(.A1(new_n1238), .A2(new_n1248), .A3(new_n1249), .A4(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1217), .ZN(new_n1252));
  OAI221_X1 g1052(.A(new_n1226), .B1(new_n854), .B2(new_n1251), .C1(new_n1252), .C2(new_n750), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n1225), .A2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(KEYINPUT57), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1196), .A2(new_n1200), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1190), .B1(new_n1202), .B2(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n700), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1212), .A2(new_n1222), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1252), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1212), .A2(new_n1222), .A3(new_n1217), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1199), .B1(new_n1195), .B2(new_n1176), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1204), .B1(new_n1181), .B2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT57), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1254), .B1(new_n1258), .B2(new_n1265), .ZN(G375));
  NAND3_X1  g1066(.A1(new_n1196), .A2(new_n1190), .A3(new_n1200), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1208), .A2(new_n1025), .A3(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n916), .A2(new_n749), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n742), .B1(G68), .B2(new_n1137), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n805), .A2(G107), .B1(G294), .B2(new_n794), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n851), .A2(G303), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n777), .A2(new_n520), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n307), .B1(new_n768), .B2(G97), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n954), .A2(new_n1272), .A3(new_n1273), .A4(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(G116), .B2(new_n781), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1271), .B(new_n1276), .C1(new_n834), .C2(new_n836), .ZN(new_n1277));
  OR2_X1    g1077(.A1(new_n1277), .A2(KEYINPUT126), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n781), .A2(new_n1148), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n851), .A2(G128), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n307), .B1(new_n767), .B2(new_n809), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1281), .B1(G50), .B2(new_n777), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1279), .A2(new_n1241), .A3(new_n1280), .A4(new_n1282), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n797), .A2(new_n960), .ZN(new_n1284));
  AOI211_X1 g1084(.A(new_n1283), .B(new_n1284), .C1(G132), .C2(new_n794), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1285), .B1(new_n799), .B2(new_n1146), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1277), .A2(KEYINPUT126), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1278), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1270), .B1(new_n1288), .B2(new_n752), .ZN(new_n1289));
  AOI22_X1  g1089(.A1(new_n1256), .A2(new_n979), .B1(new_n1269), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1268), .A2(new_n1290), .ZN(G381));
  NAND3_X1  g1091(.A1(new_n1092), .A2(new_n820), .A3(new_n1094), .ZN(new_n1292));
  OR4_X1    g1092(.A1(G384), .A2(new_n1292), .A3(G390), .A4(G381), .ZN(new_n1293));
  OR4_X1    g1093(.A1(G387), .A2(new_n1293), .A3(G378), .A4(G375), .ZN(G407));
  NAND2_X1  g1094(.A1(new_n674), .A2(G213), .ZN(new_n1295));
  OR3_X1    g1095(.A1(G375), .A2(G378), .A3(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(G407), .A2(G213), .A3(new_n1296), .ZN(G409));
  OAI211_X1 g1097(.A(G378), .B(new_n1254), .C1(new_n1258), .C2(new_n1265), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n701), .B1(new_n1208), .B2(new_n1181), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1183), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1262), .A2(new_n1025), .A3(new_n1264), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1225), .A2(new_n1253), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1301), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1298), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1295), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT60), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1267), .A2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1263), .A2(KEYINPUT60), .A3(new_n1190), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1308), .A2(new_n700), .A3(new_n1208), .A4(new_n1309), .ZN(new_n1310));
  AND3_X1   g1110(.A1(new_n1310), .A2(G384), .A3(new_n1290), .ZN(new_n1311));
  AOI21_X1  g1111(.A(G384), .B1(new_n1310), .B2(new_n1290), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT127), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n674), .A2(G213), .A3(G2897), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1313), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1315), .ZN(new_n1317));
  INV_X1    g1117(.A(G384), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1263), .A2(KEYINPUT60), .A3(new_n1190), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n700), .B1(new_n1263), .B2(new_n1190), .ZN(new_n1320));
  AOI21_X1  g1120(.A(KEYINPUT60), .B1(new_n1263), .B2(new_n1190), .ZN(new_n1321));
  NOR3_X1   g1121(.A1(new_n1319), .A2(new_n1320), .A3(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1290), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1318), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1310), .A2(G384), .A3(new_n1290), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1317), .B1(new_n1326), .B2(KEYINPUT127), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1326), .A2(KEYINPUT127), .ZN(new_n1328));
  OAI211_X1 g1128(.A(new_n1306), .B(new_n1316), .C1(new_n1327), .C2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT61), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1305), .A2(new_n1295), .A3(new_n1313), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(KEYINPUT62), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT62), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1305), .A2(new_n1333), .A3(new_n1295), .A4(new_n1313), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1329), .A2(new_n1330), .A3(new_n1332), .A4(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(G393), .A2(G396), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(new_n1292), .ZN(new_n1337));
  AND3_X1   g1137(.A1(new_n1039), .A2(new_n1046), .A3(new_n1051), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1051), .B1(new_n1039), .B2(new_n1046), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT109), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1096), .A2(new_n1341), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1342), .A2(new_n1010), .A3(new_n1017), .A4(new_n1019), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1024), .B1(new_n1343), .B2(new_n736), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1340), .B1(new_n1344), .B2(new_n979), .ZN(new_n1345));
  AOI21_X1  g1145(.A(G390), .B1(new_n1345), .B2(new_n978), .ZN(new_n1346));
  OAI211_X1 g1146(.A(G390), .B(new_n978), .C1(new_n1026), .C2(new_n1053), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1347), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1337), .B1(new_n1346), .B2(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(G390), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(G387), .A2(new_n1350), .ZN(new_n1351));
  NAND4_X1  g1151(.A1(new_n1351), .A2(new_n1292), .A3(new_n1336), .A4(new_n1347), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1349), .A2(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1335), .A2(new_n1353), .ZN(new_n1354));
  NAND4_X1  g1154(.A1(new_n1305), .A2(KEYINPUT63), .A3(new_n1295), .A4(new_n1313), .ZN(new_n1355));
  AND3_X1   g1155(.A1(new_n1349), .A2(new_n1352), .A3(new_n1355), .ZN(new_n1356));
  INV_X1    g1156(.A(KEYINPUT63), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1331), .A2(new_n1357), .ZN(new_n1358));
  NAND4_X1  g1158(.A1(new_n1356), .A2(new_n1330), .A3(new_n1329), .A4(new_n1358), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1354), .A2(new_n1359), .ZN(G405));
  NAND2_X1  g1160(.A1(G375), .A2(new_n1301), .ZN(new_n1361));
  AND3_X1   g1161(.A1(new_n1361), .A2(new_n1298), .A3(new_n1326), .ZN(new_n1362));
  AOI21_X1  g1162(.A(new_n1326), .B1(new_n1361), .B2(new_n1298), .ZN(new_n1363));
  NOR2_X1   g1163(.A1(new_n1362), .A2(new_n1363), .ZN(new_n1364));
  XOR2_X1   g1164(.A(new_n1364), .B(new_n1353), .Z(G402));
endmodule


