//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 1 1 1 1 1 1 1 1 0 1 1 0 0 0 1 1 1 1 0 1 0 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 0 1 1 1 1 1 1 1 0 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1320, new_n1321,
    new_n1322, new_n1323, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1395,
    new_n1396, new_n1397;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(KEYINPUT65), .B(G68), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G58), .A2(G232), .ZN(new_n214));
  NAND4_X1  g0014(.A1(new_n211), .A2(new_n212), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n206), .B1(new_n210), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  OR3_X1    g0017(.A1(new_n206), .A2(KEYINPUT64), .A3(G13), .ZN(new_n218));
  OAI21_X1  g0018(.A(KEYINPUT64), .B1(new_n206), .B2(G13), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT0), .Z(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(new_n201), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G50), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  AOI211_X1 g0028(.A(new_n217), .B(new_n222), .C1(new_n225), .C2(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XOR2_X1   g0038(.A(G107), .B(G116), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G58), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  INV_X1    g0044(.A(KEYINPUT73), .ZN(new_n245));
  AND2_X1   g0045(.A1(KEYINPUT3), .A2(G33), .ZN(new_n246));
  NOR2_X1   g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  OAI21_X1  g0047(.A(KEYINPUT67), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT3), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT67), .ZN(new_n252));
  NAND2_X1  g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n248), .A2(new_n254), .A3(G222), .A4(new_n255), .ZN(new_n256));
  NAND4_X1  g0056(.A1(new_n248), .A2(new_n254), .A3(G223), .A4(G1698), .ZN(new_n257));
  NOR3_X1   g0057(.A1(new_n246), .A2(new_n247), .A3(KEYINPUT67), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n252), .B1(new_n251), .B2(new_n253), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G77), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n256), .B(new_n257), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  AND2_X1   g0062(.A1(G33), .A2(G41), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(new_n223), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT66), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(new_n263), .B2(new_n223), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n268), .B1(G41), .B2(G45), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n271), .A2(KEYINPUT66), .A3(G1), .A4(G13), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n267), .A2(new_n270), .A3(G274), .A4(new_n272), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n267), .A2(G226), .A3(new_n269), .A4(new_n272), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n265), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G179), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT68), .ZN(new_n279));
  INV_X1    g0079(.A(G58), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n279), .B1(new_n280), .B2(KEYINPUT8), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT8), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(KEYINPUT68), .A3(G58), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n281), .B(new_n283), .C1(new_n282), .C2(G58), .ZN(new_n284));
  OAI21_X1  g0084(.A(KEYINPUT69), .B1(new_n250), .B2(G20), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT69), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(new_n224), .A3(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n223), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n268), .A2(G13), .A3(G20), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(G50), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n293), .A2(new_n223), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n268), .A2(KEYINPUT70), .A3(G20), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT70), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(new_n224), .B2(G1), .ZN(new_n301));
  AND4_X1   g0101(.A1(new_n298), .A2(new_n296), .A3(new_n299), .A4(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n297), .B1(new_n302), .B2(G50), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n295), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n275), .B1(new_n262), .B2(new_n264), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n304), .B1(new_n305), .B2(G169), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n278), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n295), .A2(KEYINPUT9), .A3(new_n303), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT9), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n298), .B1(new_n289), .B2(new_n291), .ZN(new_n310));
  INV_X1    g0110(.A(new_n297), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n298), .A2(new_n296), .A3(new_n299), .A4(new_n301), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n311), .B1(new_n312), .B2(new_n202), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n309), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G200), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n308), .B(new_n314), .C1(new_n305), .C2(new_n315), .ZN(new_n316));
  AND2_X1   g0116(.A1(new_n305), .A2(G190), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT10), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n308), .A2(new_n314), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n277), .A2(G200), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT10), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n305), .A2(G190), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n319), .A2(new_n320), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n307), .B1(new_n318), .B2(new_n323), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n267), .A2(G244), .A3(new_n269), .A4(new_n272), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n273), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n248), .A2(new_n254), .A3(G238), .A4(G1698), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n248), .A2(new_n254), .A3(G232), .A4(new_n255), .ZN(new_n328));
  INV_X1    g0128(.A(G107), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n327), .B(new_n328), .C1(new_n260), .C2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n326), .B1(new_n330), .B2(new_n264), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n331), .A2(G190), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT15), .B(G87), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(new_n285), .B2(new_n287), .ZN(new_n334));
  XNOR2_X1  g0134(.A(KEYINPUT8), .B(G58), .ZN(new_n335));
  INV_X1    g0135(.A(new_n290), .ZN(new_n336));
  OAI22_X1  g0136(.A1(new_n335), .A2(new_n336), .B1(new_n224), .B2(new_n261), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n294), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n302), .A2(G77), .ZN(new_n339));
  INV_X1    g0139(.A(new_n296), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n261), .ZN(new_n341));
  AND3_X1   g0141(.A1(new_n338), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(new_n331), .B2(new_n315), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n332), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n338), .A2(new_n339), .A3(new_n341), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(new_n331), .B2(G169), .ZN(new_n346));
  INV_X1    g0146(.A(G179), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n346), .A2(KEYINPUT71), .B1(new_n347), .B2(new_n331), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT71), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n345), .B(new_n349), .C1(new_n331), .C2(G169), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n344), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT72), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n324), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n346), .A2(KEYINPUT71), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n331), .A2(new_n347), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(new_n350), .A3(new_n355), .ZN(new_n356));
  OR2_X1    g0156(.A1(new_n332), .A2(new_n343), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(KEYINPUT72), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n245), .B1(new_n353), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(KEYINPUT72), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n351), .A2(new_n352), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n361), .A2(new_n362), .A3(KEYINPUT73), .A4(new_n324), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n208), .A2(G20), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(G50), .B2(new_n290), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n288), .A2(G77), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n298), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT11), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT12), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n296), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G13), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n373), .A2(G1), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT12), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n370), .B(new_n372), .C1(new_n365), .C2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(G68), .B1(new_n302), .B2(new_n371), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n369), .B2(KEYINPUT11), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n248), .A2(new_n254), .A3(G232), .A4(G1698), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n248), .A2(new_n254), .A3(G226), .A4(new_n255), .ZN(new_n381));
  NAND2_X1  g0181(.A1(G33), .A2(G97), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n264), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n267), .A2(G238), .A3(new_n269), .A4(new_n272), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n273), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT13), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT13), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n384), .A2(new_n390), .A3(new_n387), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(G200), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n389), .A2(G190), .A3(new_n391), .ZN(new_n394));
  AND3_X1   g0194(.A1(new_n379), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT14), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(new_n392), .B2(G169), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n390), .B1(new_n384), .B2(new_n387), .ZN(new_n398));
  AOI211_X1 g0198(.A(KEYINPUT13), .B(new_n386), .C1(new_n383), .C2(new_n264), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n396), .B(G169), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n389), .A2(G179), .A3(new_n391), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(KEYINPUT74), .B1(new_n397), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(G169), .B1(new_n398), .B2(new_n399), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT14), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT74), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n405), .A2(new_n406), .A3(new_n401), .A4(new_n400), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n379), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n395), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n207), .A2(G58), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n226), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n412), .A2(G20), .B1(G159), .B2(new_n290), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n251), .A2(new_n224), .A3(new_n253), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT7), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NOR3_X1   g0216(.A1(new_n246), .A2(new_n247), .A3(G20), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT75), .B1(new_n417), .B2(KEYINPUT7), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT75), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n414), .A2(new_n419), .A3(new_n415), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n416), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(G68), .ZN(new_n422));
  OAI211_X1 g0222(.A(KEYINPUT16), .B(new_n413), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n201), .B1(new_n207), .B2(G58), .ZN(new_n424));
  INV_X1    g0224(.A(G159), .ZN(new_n425));
  OAI22_X1  g0225(.A1(new_n424), .A2(new_n224), .B1(new_n425), .B2(new_n336), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n417), .A2(KEYINPUT7), .ZN(new_n427));
  AOI21_X1  g0227(.A(G20), .B1(new_n248), .B2(new_n254), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n427), .B1(new_n428), .B2(KEYINPUT7), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n426), .B1(new_n429), .B2(new_n207), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n423), .B(new_n294), .C1(KEYINPUT16), .C2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(G223), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n255), .ZN(new_n433));
  INV_X1    g0233(.A(G226), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(G1698), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n433), .B(new_n435), .C1(new_n246), .C2(new_n247), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G33), .A2(G87), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT76), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n436), .A2(KEYINPUT76), .A3(new_n437), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n440), .A2(new_n264), .A3(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n267), .A2(G232), .A3(new_n269), .A4(new_n272), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n273), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n442), .A2(G190), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n315), .B1(new_n442), .B2(new_n445), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n284), .A2(new_n340), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n449), .B1(new_n312), .B2(new_n284), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n431), .A2(new_n448), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT17), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n431), .A2(new_n448), .A3(KEYINPUT17), .A4(new_n451), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n442), .ZN(new_n457));
  OAI21_X1  g0257(.A(G169), .B1(new_n457), .B2(new_n444), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n442), .A2(G179), .A3(new_n445), .ZN(new_n459));
  AOI221_X4 g0259(.A(KEYINPUT18), .B1(new_n458), .B2(new_n459), .C1(new_n431), .C2(new_n451), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT18), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n294), .B1(new_n430), .B2(KEYINPUT16), .ZN(new_n462));
  INV_X1    g0262(.A(new_n423), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n451), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n458), .A2(new_n459), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n460), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n456), .A2(new_n467), .A3(KEYINPUT77), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n224), .B1(new_n258), .B2(new_n259), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n416), .B1(new_n469), .B2(new_n415), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n413), .B1(new_n470), .B2(new_n208), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT16), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n298), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n450), .B1(new_n473), .B2(new_n423), .ZN(new_n474));
  INV_X1    g0274(.A(new_n465), .ZN(new_n475));
  OAI21_X1  g0275(.A(KEYINPUT18), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n464), .A2(new_n461), .A3(new_n465), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n476), .A2(new_n477), .A3(new_n454), .A4(new_n455), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT77), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n468), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n364), .A2(new_n410), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT78), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n481), .A2(new_n410), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n485), .A2(KEYINPUT78), .A3(new_n364), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(G116), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n340), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n268), .A2(G33), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n298), .A2(G116), .A3(new_n296), .A4(new_n490), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n293), .A2(new_n223), .B1(G20), .B2(new_n488), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G33), .A2(G283), .ZN(new_n493));
  INV_X1    g0293(.A(G97), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n493), .B(new_n224), .C1(G33), .C2(new_n494), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n492), .A2(KEYINPUT20), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT20), .B1(new_n492), .B2(new_n495), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n489), .B(new_n491), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n264), .ZN(new_n499));
  OAI21_X1  g0299(.A(G303), .B1(new_n258), .B2(new_n259), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n251), .A2(new_n253), .ZN(new_n501));
  OR2_X1    g0301(.A1(new_n255), .A2(G264), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n501), .B(new_n502), .C1(G257), .C2(G1698), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n499), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n268), .A2(G45), .ZN(new_n505));
  OR2_X1    g0305(.A1(KEYINPUT5), .A2(G41), .ZN(new_n506));
  NAND2_X1  g0306(.A1(KEYINPUT5), .A2(G41), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n508), .A2(G274), .A3(new_n267), .A4(new_n272), .ZN(new_n509));
  AND2_X1   g0309(.A1(KEYINPUT5), .A2(G41), .ZN(new_n510));
  NOR2_X1   g0310(.A1(KEYINPUT5), .A2(G41), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n268), .B(G45), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n512), .A2(new_n267), .A3(G270), .A4(new_n272), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n498), .B(G169), .C1(new_n504), .C2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT85), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(KEYINPUT21), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT21), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n515), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n503), .ZN(new_n521));
  INV_X1    g0321(.A(G303), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n522), .B1(new_n248), .B2(new_n254), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n264), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n509), .A2(new_n513), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n526), .A2(new_n347), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n498), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n524), .A2(new_n525), .A3(G190), .ZN(new_n529));
  INV_X1    g0329(.A(new_n498), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n504), .A2(new_n514), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n529), .B(new_n530), .C1(new_n531), .C2(new_n315), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n518), .A2(new_n520), .A3(new_n528), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT86), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n517), .A2(KEYINPUT21), .B1(new_n527), .B2(new_n498), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT86), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n535), .A2(new_n536), .A3(new_n520), .A4(new_n532), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n267), .A2(new_n272), .ZN(new_n539));
  INV_X1    g0339(.A(G45), .ZN(new_n540));
  OAI211_X1 g0340(.A(KEYINPUT80), .B(G250), .C1(new_n540), .C2(G1), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT80), .ZN(new_n542));
  AOI21_X1  g0342(.A(G274), .B1(new_n542), .B2(G250), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n541), .B1(new_n543), .B2(new_n505), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n209), .A2(new_n255), .ZN(new_n545));
  INV_X1    g0345(.A(G244), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G1698), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n545), .B(new_n547), .C1(new_n246), .C2(new_n247), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G116), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n539), .A2(new_n544), .B1(new_n550), .B2(new_n264), .ZN(new_n551));
  AOI21_X1  g0351(.A(KEYINPUT84), .B1(new_n551), .B2(G190), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n550), .A2(new_n264), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n544), .A2(new_n267), .A3(new_n272), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(G190), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n551), .B2(new_n315), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n552), .B1(KEYINPUT84), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n333), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n558), .A2(new_n296), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n296), .A2(new_n490), .A3(new_n223), .A4(new_n293), .ZN(new_n560));
  INV_X1    g0360(.A(G87), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n288), .A2(G97), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT82), .ZN(new_n564));
  OR2_X1    g0364(.A1(KEYINPUT81), .A2(KEYINPUT19), .ZN(new_n565));
  NAND2_X1  g0365(.A1(KEYINPUT81), .A2(KEYINPUT19), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n563), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n494), .B1(new_n285), .B2(new_n287), .ZN(new_n570));
  OAI21_X1  g0370(.A(KEYINPUT82), .B1(new_n570), .B2(new_n567), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n501), .A2(new_n224), .A3(G68), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n561), .A2(new_n494), .A3(new_n329), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n382), .B1(new_n565), .B2(new_n566), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n573), .B1(new_n574), .B2(G20), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n569), .A2(new_n571), .A3(new_n572), .A4(new_n575), .ZN(new_n576));
  AOI211_X1 g0376(.A(new_n559), .B(new_n562), .C1(new_n576), .C2(new_n294), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n557), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n512), .A2(new_n267), .A3(G264), .A4(new_n272), .ZN(new_n579));
  NOR2_X1   g0379(.A1(G250), .A2(G1698), .ZN(new_n580));
  INV_X1    g0380(.A(G257), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n580), .B1(new_n581), .B2(G1698), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n582), .A2(new_n501), .B1(G33), .B2(G294), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n509), .B(new_n579), .C1(new_n583), .C2(new_n499), .ZN(new_n584));
  INV_X1    g0384(.A(G169), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n581), .A2(G1698), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(G250), .B2(G1698), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n246), .A2(new_n247), .ZN(new_n589));
  INV_X1    g0389(.A(G294), .ZN(new_n590));
  OAI22_X1  g0390(.A1(new_n588), .A2(new_n589), .B1(new_n250), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n264), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n592), .A2(new_n347), .A3(new_n509), .A4(new_n579), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n586), .A2(new_n593), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n561), .A2(KEYINPUT22), .A3(G20), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n248), .A2(new_n254), .A3(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n224), .B(G87), .C1(new_n246), .C2(new_n247), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(KEYINPUT22), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(KEYINPUT88), .B(KEYINPUT23), .C1(new_n224), .C2(G107), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n224), .A2(G33), .A3(G116), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n329), .A2(G20), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n600), .B(new_n601), .C1(KEYINPUT23), .C2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(KEYINPUT88), .B1(new_n602), .B2(KEYINPUT23), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g0406(.A(KEYINPUT87), .B(KEYINPUT24), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n599), .A2(new_n605), .A3(new_n607), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n298), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n340), .A2(KEYINPUT25), .A3(new_n329), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT25), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n296), .B2(G107), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n329), .B2(new_n560), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n594), .B1(new_n611), .B2(new_n616), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n599), .A2(new_n605), .A3(new_n607), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n607), .B1(new_n599), .B2(new_n605), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n294), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n616), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n584), .A2(new_n315), .ZN(new_n622));
  INV_X1    g0422(.A(G190), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n592), .A2(new_n623), .A3(new_n509), .A4(new_n579), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n620), .A2(new_n621), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n576), .A2(new_n294), .ZN(new_n627));
  INV_X1    g0427(.A(new_n559), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT83), .ZN(new_n629));
  OR3_X1    g0429(.A1(new_n560), .A2(new_n629), .A3(new_n333), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n629), .B1(new_n560), .B2(new_n333), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n627), .A2(new_n628), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n551), .A2(G179), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n553), .A2(new_n554), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(G169), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n578), .A2(new_n617), .A3(new_n626), .A4(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n429), .A2(G107), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT6), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n642), .A2(new_n494), .A3(G107), .ZN(new_n643));
  XNOR2_X1  g0443(.A(G97), .B(G107), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n643), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  OAI22_X1  g0445(.A1(new_n645), .A2(new_n224), .B1(new_n261), .B2(new_n336), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n298), .B1(new_n641), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n340), .A2(new_n494), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n560), .B2(new_n494), .ZN(new_n650));
  OAI21_X1  g0450(.A(KEYINPUT79), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT79), .ZN(new_n652));
  INV_X1    g0452(.A(new_n650), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n646), .B1(new_n429), .B2(G107), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n652), .B(new_n653), .C1(new_n654), .C2(new_n298), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n512), .A2(new_n267), .A3(G257), .A4(new_n272), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n509), .A2(new_n656), .ZN(new_n657));
  OAI211_X1 g0457(.A(G244), .B(new_n255), .C1(new_n246), .C2(new_n247), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT4), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n658), .A2(new_n659), .B1(G33), .B2(G283), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n546), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n248), .A2(new_n254), .A3(new_n255), .A4(new_n661), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n248), .A2(new_n254), .A3(G250), .A4(G1698), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n660), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n657), .B1(new_n664), .B2(new_n264), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(G169), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(G179), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n651), .A2(new_n655), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n653), .B1(new_n654), .B2(new_n298), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n665), .A2(new_n315), .ZN(new_n671));
  AOI211_X1 g0471(.A(new_n623), .B(new_n657), .C1(new_n264), .C2(new_n664), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n640), .A2(new_n669), .A3(new_n673), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n487), .A2(new_n538), .A3(new_n674), .ZN(G372));
  INV_X1    g0475(.A(KEYINPUT89), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n651), .A2(new_n655), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n667), .A2(new_n668), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n673), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n315), .B1(new_n553), .B2(new_n554), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n680), .B1(G190), .B2(new_n551), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n559), .B1(new_n576), .B2(new_n294), .ZN(new_n682));
  INV_X1    g0482(.A(new_n562), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n639), .A2(new_n626), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n676), .B1(new_n679), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n639), .A2(new_n626), .A3(new_n684), .ZN(new_n687));
  NOR4_X1   g0487(.A1(new_n669), .A2(new_n687), .A3(new_n673), .A4(KEYINPUT89), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n617), .A2(new_n518), .A3(new_n520), .A4(new_n528), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT90), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n535), .A2(KEYINPUT90), .A3(new_n520), .A4(new_n617), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n686), .A2(new_n688), .A3(new_n693), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n557), .A2(new_n577), .B1(new_n634), .B2(new_n638), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n669), .A2(KEYINPUT26), .A3(new_n695), .ZN(new_n696));
  AOI22_X1  g0496(.A1(new_n577), .A2(new_n681), .B1(new_n634), .B2(new_n638), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n641), .A2(new_n647), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n294), .ZN(new_n699));
  AOI22_X1  g0499(.A1(new_n667), .A2(new_n668), .B1(new_n699), .B2(new_n653), .ZN(new_n700));
  AOI21_X1  g0500(.A(KEYINPUT26), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n696), .B1(new_n701), .B2(KEYINPUT91), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT26), .ZN(new_n703));
  AOI211_X1 g0503(.A(new_n559), .B(new_n632), .C1(new_n576), .C2(new_n294), .ZN(new_n704));
  INV_X1    g0504(.A(new_n638), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n627), .A2(new_n628), .A3(new_n683), .ZN(new_n706));
  OAI22_X1  g0506(.A1(new_n704), .A2(new_n705), .B1(new_n706), .B2(new_n556), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n665), .A2(G179), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n665), .A2(new_n585), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n670), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n703), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT91), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n639), .B1(new_n702), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n487), .B1(new_n694), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n318), .A2(new_n323), .ZN(new_n716));
  INV_X1    g0516(.A(new_n456), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n400), .A2(new_n401), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n406), .B1(new_n718), .B2(new_n405), .ZN(new_n719));
  AND4_X1   g0519(.A1(new_n406), .A2(new_n405), .A3(new_n401), .A4(new_n400), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n409), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n379), .A2(new_n393), .A3(new_n394), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(new_n350), .A3(new_n348), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n717), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n467), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n716), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n307), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n715), .A2(new_n729), .ZN(G369));
  AND2_X1   g0530(.A1(new_n617), .A2(new_n626), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n374), .A2(new_n224), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n732), .A2(KEYINPUT27), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(KEYINPUT27), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n733), .A2(new_n734), .A3(G213), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT92), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G343), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n738), .B1(new_n611), .B2(new_n616), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n731), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n617), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n738), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n535), .A2(new_n520), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n737), .A2(new_n530), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT93), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n746), .B(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n745), .B1(new_n534), .B2(new_n537), .ZN(new_n749));
  OAI211_X1 g0549(.A(G330), .B(new_n743), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n738), .B1(new_n535), .B2(new_n520), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n751), .A2(new_n731), .B1(new_n741), .B2(new_n737), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n750), .A2(new_n752), .ZN(G399));
  INV_X1    g0553(.A(new_n220), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G41), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n573), .A2(G116), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n755), .A2(new_n268), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(new_n228), .B2(new_n755), .ZN(new_n759));
  XNOR2_X1  g0559(.A(KEYINPUT94), .B(KEYINPUT28), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n677), .A2(new_n678), .ZN(new_n762));
  INV_X1    g0562(.A(new_n673), .ZN(new_n763));
  AND4_X1   g0563(.A1(new_n762), .A2(new_n685), .A3(new_n689), .A4(new_n763), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n695), .A2(new_n677), .A3(new_n703), .A4(new_n678), .ZN(new_n765));
  OAI21_X1  g0565(.A(KEYINPUT26), .B1(new_n707), .B2(new_n710), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n765), .A2(new_n766), .A3(new_n639), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT29), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n768), .A2(new_n769), .A3(new_n738), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n737), .B1(new_n694), .B2(new_n714), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n770), .B1(new_n771), .B2(new_n769), .ZN(new_n772));
  INV_X1    g0572(.A(G330), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n674), .A2(new_n538), .A3(new_n737), .ZN(new_n774));
  AND3_X1   g0574(.A1(new_n551), .A2(new_n579), .A3(new_n592), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n775), .A2(new_n531), .A3(new_n665), .A4(G179), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT30), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n527), .A2(KEYINPUT30), .A3(new_n665), .A4(new_n775), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n551), .A2(G179), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n666), .A2(new_n526), .A3(new_n584), .A4(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n778), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  AND3_X1   g0582(.A1(new_n782), .A2(KEYINPUT31), .A3(new_n738), .ZN(new_n783));
  AOI21_X1  g0583(.A(KEYINPUT31), .B1(new_n782), .B2(new_n738), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n773), .B1(new_n774), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n772), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n761), .B1(new_n787), .B2(G1), .ZN(G364));
  OAI21_X1  g0588(.A(G330), .B1(new_n748), .B2(new_n749), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n373), .A2(G20), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n268), .B1(new_n790), .B2(G45), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n755), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n789), .A2(new_n794), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n748), .A2(new_n749), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n795), .B1(G330), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n260), .A2(G355), .A3(new_n220), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n754), .A2(new_n501), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(G45), .B2(new_n227), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n243), .A2(new_n540), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n798), .B1(G116), .B2(new_n220), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(G13), .A2(G33), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT95), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(G20), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n223), .B1(G20), .B2(new_n585), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n794), .B1(new_n802), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(KEYINPUT96), .ZN(new_n809));
  INV_X1    g0609(.A(new_n806), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n224), .A2(G179), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n811), .A2(G190), .A3(G200), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n561), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n224), .A2(new_n347), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n814), .A2(G190), .A3(new_n315), .ZN(new_n815));
  NOR2_X1   g0615(.A1(G190), .A2(G200), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n260), .B1(new_n280), .B2(new_n815), .C1(new_n261), .C2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT32), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n811), .A2(new_n816), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(new_n425), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n813), .B(new_n818), .C1(new_n819), .C2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n814), .A2(G200), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(G190), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n823), .A2(new_n623), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n825), .A2(new_n422), .B1(new_n827), .B2(new_n202), .ZN(new_n828));
  NOR3_X1   g0628(.A1(new_n623), .A2(G179), .A3(G200), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n829), .A2(new_n224), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n821), .A2(new_n819), .B1(new_n830), .B2(new_n494), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n811), .A2(new_n623), .A3(G200), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT97), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n833), .A2(new_n834), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n822), .B(new_n832), .C1(new_n329), .C2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n826), .A2(G326), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n590), .B2(new_n830), .ZN(new_n840));
  XNOR2_X1  g0640(.A(KEYINPUT33), .B(G317), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n840), .B1(new_n824), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(G322), .ZN(new_n843));
  INV_X1    g0643(.A(G311), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n815), .A2(new_n843), .B1(new_n817), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n820), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n845), .B1(G329), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n837), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(G283), .ZN(new_n849));
  INV_X1    g0649(.A(new_n812), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n260), .B1(G303), .B2(new_n850), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n842), .A2(new_n847), .A3(new_n849), .A4(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n810), .B1(new_n838), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n808), .A2(KEYINPUT96), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n805), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n809), .B(new_n855), .C1(new_n796), .C2(new_n856), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n797), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(G396));
  NAND2_X1  g0659(.A1(new_n738), .A2(new_n345), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n356), .A2(new_n357), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(new_n356), .B2(new_n860), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n771), .A2(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n737), .B(new_n862), .C1(new_n694), .C2(new_n714), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n786), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n866), .A2(new_n793), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n864), .A2(new_n786), .A3(new_n865), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n848), .A2(G87), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n844), .B2(new_n820), .ZN(new_n871));
  XOR2_X1   g0671(.A(new_n871), .B(KEYINPUT99), .Z(new_n872));
  INV_X1    g0672(.A(new_n260), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n873), .B1(new_n488), .B2(new_n817), .C1(new_n590), .C2(new_n815), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n824), .A2(G283), .B1(new_n850), .B2(G107), .ZN(new_n875));
  OAI221_X1 g0675(.A(new_n875), .B1(new_n494), .B2(new_n830), .C1(new_n522), .C2(new_n827), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n872), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n848), .A2(G68), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n589), .B1(new_n846), .B2(G132), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n280), .B2(new_n830), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n880), .B1(G50), .B2(new_n850), .ZN(new_n881));
  INV_X1    g0681(.A(new_n815), .ZN(new_n882));
  INV_X1    g0682(.A(new_n817), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n882), .A2(G143), .B1(new_n883), .B2(G159), .ZN(new_n884));
  INV_X1    g0684(.A(G150), .ZN(new_n885));
  INV_X1    g0685(.A(G137), .ZN(new_n886));
  OAI221_X1 g0686(.A(new_n884), .B1(new_n825), .B2(new_n885), .C1(new_n886), .C2(new_n827), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT34), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n878), .B(new_n881), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(new_n888), .B2(new_n887), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n806), .B1(new_n877), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n803), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n810), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n793), .B1(G77), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT98), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n896), .B(KEYINPUT100), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n804), .B2(new_n862), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n869), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(G384));
  INV_X1    g0700(.A(new_n645), .ZN(new_n901));
  OR2_X1    g0701(.A1(new_n901), .A2(KEYINPUT35), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(KEYINPUT35), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n902), .A2(G116), .A3(new_n225), .A4(new_n903), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n904), .B(KEYINPUT36), .Z(new_n905));
  NAND3_X1  g0705(.A1(new_n228), .A2(new_n411), .A3(G77), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n202), .A2(G68), .ZN(new_n907));
  AOI211_X1 g0707(.A(new_n268), .B(G13), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n774), .A2(new_n785), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n862), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n379), .A2(new_n737), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n721), .A2(new_n722), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n379), .B1(new_n403), .B2(new_n407), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n912), .B1(new_n915), .B2(new_n395), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n911), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT38), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n464), .A2(new_n465), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n464), .A2(new_n736), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT37), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n919), .A2(new_n920), .A3(new_n921), .A4(new_n452), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n413), .B1(new_n421), .B2(new_n422), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n298), .B1(new_n924), .B2(new_n472), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n423), .B1(new_n925), .B2(KEYINPUT102), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n414), .A2(new_n419), .A3(new_n415), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n419), .B1(new_n414), .B2(new_n415), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n427), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n426), .B1(new_n929), .B2(G68), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n294), .B1(new_n930), .B2(KEYINPUT16), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT102), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n451), .B1(new_n926), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n465), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n736), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n935), .A2(new_n936), .A3(new_n452), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n923), .B1(new_n937), .B2(KEYINPUT37), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n936), .B1(new_n456), .B2(new_n467), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n918), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n463), .B1(new_n931), .B2(new_n932), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n925), .A2(KEYINPUT102), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n450), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n736), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n452), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n943), .A2(new_n475), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT37), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n922), .ZN(new_n948));
  INV_X1    g0748(.A(new_n939), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n948), .A2(KEYINPUT38), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n940), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n917), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT40), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n919), .A2(new_n920), .A3(new_n452), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(KEYINPUT37), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n922), .ZN(new_n956));
  INV_X1    g0756(.A(new_n920), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n478), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(KEYINPUT38), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n953), .B1(new_n950), .B2(new_n960), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n952), .A2(new_n953), .B1(new_n917), .B2(new_n961), .ZN(new_n962));
  AND3_X1   g0762(.A1(new_n962), .A2(new_n487), .A3(new_n910), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n962), .B1(new_n487), .B2(new_n910), .ZN(new_n964));
  OR3_X1    g0764(.A1(new_n963), .A2(new_n964), .A3(new_n773), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n950), .A2(new_n960), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT39), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n721), .A2(new_n738), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n940), .A2(new_n950), .A3(KEYINPUT39), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n348), .A2(new_n350), .A3(new_n737), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT101), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n865), .A2(new_n973), .B1(new_n914), .B2(new_n916), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n951), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n725), .A2(new_n944), .ZN(new_n976));
  AND3_X1   g0776(.A1(new_n971), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n728), .B1(new_n487), .B2(new_n772), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n977), .B(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n965), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n268), .B2(new_n790), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n965), .A2(new_n979), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n909), .B1(new_n981), .B2(new_n982), .ZN(G367));
  INV_X1    g0783(.A(new_n787), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n738), .A2(new_n670), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n762), .A2(new_n763), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n700), .A2(new_n738), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n752), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT45), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n989), .B(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT44), .ZN(new_n992));
  OR3_X1    g0792(.A1(new_n988), .A2(new_n752), .A3(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n992), .B1(new_n988), .B2(new_n752), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n991), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n750), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n991), .A2(new_n750), .A3(new_n995), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT105), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n751), .A2(new_n731), .ZN(new_n1002));
  OAI211_X1 g0802(.A(KEYINPUT104), .B(new_n1002), .C1(new_n743), .C2(new_n751), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(KEYINPUT104), .B2(new_n1002), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(new_n789), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1000), .A2(new_n1001), .A3(new_n787), .A4(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n787), .A2(new_n1005), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n998), .A2(new_n999), .ZN(new_n1008));
  OAI21_X1  g0808(.A(KEYINPUT105), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n984), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n755), .B(KEYINPUT41), .Z(new_n1011));
  OAI21_X1  g0811(.A(new_n791), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n988), .A2(new_n731), .A3(new_n751), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT42), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n988), .A2(new_n741), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n738), .B1(new_n1015), .B2(new_n762), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT43), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n737), .A2(new_n577), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n639), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n697), .B2(new_n1018), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT103), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n1014), .A2(new_n1016), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1017), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1022), .B(new_n1023), .Z(new_n1024));
  INV_X1    g0824(.A(new_n988), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n750), .A2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1024), .B(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1012), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1021), .A2(new_n805), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n799), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1030), .A2(new_n236), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n807), .B1(new_n220), .B2(new_n333), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n793), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n825), .A2(new_n590), .B1(new_n329), .B2(new_n830), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G311), .B2(new_n826), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n812), .A2(new_n488), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1036), .A2(KEYINPUT46), .ZN(new_n1037));
  INV_X1    g0837(.A(G283), .ZN(new_n1038));
  INV_X1    g0838(.A(G317), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n817), .A2(new_n1038), .B1(new_n820), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n589), .B1(new_n815), .B2(new_n522), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1040), .B(new_n1041), .C1(KEYINPUT46), .C2(new_n1036), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n848), .A2(G97), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1035), .A2(new_n1037), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n837), .A2(new_n261), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n812), .A2(new_n280), .B1(new_n820), .B2(new_n886), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1045), .B1(KEYINPUT106), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(KEYINPUT106), .B2(new_n1046), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(G143), .A2(new_n826), .B1(new_n824), .B2(G159), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n882), .A2(G150), .B1(new_n883), .B2(G50), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n830), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(G68), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1049), .A2(new_n260), .A3(new_n1050), .A4(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1044), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT47), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1033), .B1(new_n1055), .B2(new_n806), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n1029), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1028), .A2(new_n1058), .ZN(G387));
  NOR2_X1   g0859(.A1(new_n787), .A2(new_n1005), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(KEYINPUT109), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1061), .A2(new_n755), .A3(new_n1007), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1060), .A2(KEYINPUT109), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n740), .A2(new_n742), .A3(new_n805), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n260), .A2(new_n220), .A3(new_n757), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(G107), .B2(new_n220), .ZN(new_n1067));
  AOI211_X1 g0867(.A(G45), .B(new_n757), .C1(G68), .C2(G77), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT107), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n335), .A2(G50), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT50), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1070), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1030), .B1(new_n233), .B2(G45), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1067), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n807), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n793), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT108), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n815), .A2(new_n202), .B1(new_n820), .B2(new_n885), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n589), .B(new_n1080), .C1(G68), .C2(new_n883), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n812), .A2(new_n261), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n830), .A2(new_n333), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1082), .B(new_n1083), .C1(G159), .C2(new_n826), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n824), .A2(new_n284), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1081), .A2(new_n1084), .A3(new_n1043), .A4(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n501), .B1(new_n846), .B2(G326), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n830), .A2(new_n1038), .B1(new_n812), .B2(new_n590), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n882), .A2(G317), .B1(new_n883), .B2(G303), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1089), .B1(new_n825), .B2(new_n844), .C1(new_n843), .C2(new_n827), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT48), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1088), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n1091), .B2(new_n1090), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT49), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n1087), .B1(new_n488), .B2(new_n837), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1086), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1079), .B1(new_n806), .B2(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1005), .A2(new_n792), .B1(new_n1065), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1064), .A2(new_n1099), .ZN(G393));
  NAND2_X1  g0900(.A1(new_n1000), .A2(new_n792), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1025), .A2(new_n805), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT110), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n799), .A2(new_n240), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1105), .B(new_n807), .C1(new_n494), .C2(new_n220), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT111), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n794), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n1107), .B2(new_n1106), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(G317), .A2(new_n826), .B1(new_n882), .B2(G311), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n848), .A2(G107), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n824), .A2(G303), .B1(new_n850), .B2(G283), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G294), .A2(new_n883), .B1(new_n846), .B2(G322), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1051), .A2(G116), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1114), .A2(new_n1115), .A3(new_n873), .A4(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(G143), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n501), .B1(new_n820), .B2(new_n1118), .C1(new_n335), .C2(new_n817), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n824), .A2(G50), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n830), .A2(new_n261), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(new_n207), .B2(new_n850), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n870), .A2(new_n1120), .A3(new_n1121), .A4(new_n1123), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(G150), .A2(new_n826), .B1(new_n882), .B2(G159), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT51), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n1113), .A2(new_n1117), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1109), .B1(new_n806), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1104), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT113), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n755), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1130), .A2(new_n1131), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1131), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1101), .B(new_n1129), .C1(new_n1135), .C2(new_n1136), .ZN(G390));
  INV_X1    g0937(.A(KEYINPUT115), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT114), .ZN(new_n1139));
  AOI21_X1  g0939(.A(KEYINPUT78), .B1(new_n485), .B2(new_n364), .ZN(new_n1140));
  AND4_X1   g0940(.A1(KEYINPUT78), .A2(new_n364), .A3(new_n410), .A4(new_n481), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n772), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n786), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1142), .A2(new_n1143), .A3(new_n729), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n910), .A2(G330), .A3(new_n862), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1145), .A2(new_n914), .A3(new_n916), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n913), .B1(new_n721), .B2(new_n722), .ZN(new_n1147));
  NOR3_X1   g0947(.A1(new_n915), .A2(new_n395), .A3(new_n912), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n786), .B(new_n862), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n862), .B(new_n737), .C1(new_n764), .C2(new_n767), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1150), .A2(new_n972), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1146), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1146), .A2(new_n1149), .B1(new_n865), .B2(new_n973), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1139), .B1(new_n1144), .B2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1146), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1146), .A2(new_n1149), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n973), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n639), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n695), .A2(new_n678), .A3(new_n677), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n1160), .A2(KEYINPUT26), .B1(new_n711), .B2(new_n712), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n713), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1159), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n762), .A2(new_n685), .A3(new_n763), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(KEYINPUT89), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n679), .A2(new_n676), .A3(new_n685), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1165), .A2(new_n1166), .A3(new_n691), .A4(new_n692), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n738), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1158), .B1(new_n1168), .B2(new_n862), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1156), .B1(new_n1157), .B2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1170), .A2(new_n978), .A3(KEYINPUT114), .A4(new_n1143), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1155), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1149), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n939), .B1(new_n922), .B2(new_n947), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n959), .B1(new_n1174), .B2(KEYINPUT38), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n914), .A2(new_n916), .B1(new_n1150), .B2(new_n972), .ZN(new_n1176));
  NOR3_X1   g0976(.A1(new_n1175), .A2(new_n1176), .A3(new_n969), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n969), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1178), .B1(new_n1169), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n968), .A2(new_n970), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1173), .B(new_n1177), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1175), .A2(KEYINPUT39), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n940), .A2(new_n950), .A3(KEYINPUT39), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n1183), .A2(new_n1184), .B1(new_n974), .B2(new_n969), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1177), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1149), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1182), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1138), .B1(new_n1172), .B2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1132), .B1(new_n1172), .B2(new_n1188), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n865), .A2(new_n973), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1179), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1193), .A2(new_n1178), .B1(new_n968), .B2(new_n970), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1173), .B1(new_n1194), .B2(new_n1177), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1185), .A2(new_n1149), .A3(new_n1186), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1197), .A2(KEYINPUT115), .A3(new_n1155), .A4(new_n1171), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1189), .A2(new_n1190), .A3(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n804), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1181), .A2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n793), .B1(new_n284), .B2(new_n893), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n827), .A2(new_n1038), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1122), .B(new_n1203), .C1(G107), .C2(new_n824), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n815), .A2(new_n488), .B1(new_n820), .B2(new_n590), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(G97), .B2(new_n883), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n260), .A2(new_n813), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1204), .A2(new_n878), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n873), .B1(G159), .B2(new_n1051), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n846), .A2(G125), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(KEYINPUT54), .B(G143), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n882), .A2(G132), .B1(new_n883), .B2(new_n1212), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G128), .A2(new_n826), .B1(new_n824), .B2(G137), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1209), .A2(new_n1210), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n812), .A2(new_n885), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1216), .B(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n202), .B2(new_n837), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1208), .B1(new_n1215), .B2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1202), .B1(new_n1220), .B2(new_n806), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1188), .A2(new_n792), .B1(new_n1201), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1199), .A2(new_n1222), .ZN(G378));
  INV_X1    g1023(.A(KEYINPUT57), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1144), .B1(new_n1172), .B2(new_n1188), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n736), .A2(new_n304), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n324), .A2(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n324), .A2(new_n1226), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  OR3_X1    g1030(.A1(new_n1227), .A2(new_n1228), .A3(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1230), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n962), .A2(G330), .A3(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n961), .A2(new_n917), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n863), .B1(new_n774), .B2(new_n785), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n950), .B2(new_n940), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1235), .B(G330), .C1(new_n1238), .C2(KEYINPUT40), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1233), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1234), .A2(new_n1241), .A3(new_n977), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n977), .B1(new_n1234), .B2(new_n1241), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1224), .B1(new_n1225), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1234), .A2(new_n1241), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n977), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1234), .A2(new_n1241), .A3(new_n977), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1197), .B1(new_n1155), .B2(new_n1171), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1250), .B(KEYINPUT57), .C1(new_n1251), .C2(new_n1144), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1245), .A2(new_n1252), .A3(new_n755), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1240), .A2(new_n1200), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n793), .B1(G50), .B2(new_n893), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n825), .A2(new_n494), .B1(new_n827), .B2(new_n488), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1082), .B(new_n1256), .C1(G68), .C2(new_n1051), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n848), .A2(G58), .ZN(new_n1258));
  OR2_X1    g1058(.A1(new_n501), .A2(G41), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(G283), .B2(new_n846), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n882), .A2(G107), .B1(new_n883), .B2(new_n558), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1257), .A2(new_n1258), .A3(new_n1260), .A4(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT58), .ZN(new_n1263));
  INV_X1    g1063(.A(G41), .ZN(new_n1264));
  AOI21_X1  g1064(.A(G50), .B1(new_n250), .B2(new_n1264), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n1262), .A2(new_n1263), .B1(new_n1259), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(G128), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n815), .A2(new_n1267), .B1(new_n817), .B2(new_n886), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n824), .A2(G132), .B1(new_n850), .B2(new_n1212), .ZN(new_n1269));
  INV_X1    g1069(.A(G125), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1269), .B1(new_n1270), .B2(new_n827), .ZN(new_n1271));
  AOI211_X1 g1071(.A(new_n1268), .B(new_n1271), .C1(G150), .C2(new_n1051), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1273), .A2(KEYINPUT59), .ZN(new_n1274));
  AOI211_X1 g1074(.A(G33), .B(G41), .C1(new_n846), .C2(G124), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT59), .ZN(new_n1276));
  OAI221_X1 g1076(.A(new_n1275), .B1(new_n425), .B2(new_n837), .C1(new_n1272), .C2(new_n1276), .ZN(new_n1277));
  OAI221_X1 g1077(.A(new_n1266), .B1(new_n1263), .B2(new_n1262), .C1(new_n1274), .C2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1255), .B1(new_n1278), .B2(new_n806), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1254), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1281), .B1(new_n1250), .B2(new_n792), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1253), .A2(new_n1282), .ZN(G375));
  AOI211_X1 g1083(.A(new_n1011), .B(new_n1172), .C1(new_n1144), .C2(new_n1154), .ZN(new_n1284));
  XOR2_X1   g1084(.A(new_n1284), .B(KEYINPUT117), .Z(new_n1285));
  XOR2_X1   g1085(.A(new_n791), .B(KEYINPUT118), .Z(new_n1286));
  OR2_X1    g1086(.A1(new_n1154), .A2(new_n1286), .ZN(new_n1287));
  OR2_X1    g1087(.A1(new_n1287), .A2(KEYINPUT119), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n793), .B1(G68), .B2(new_n893), .ZN(new_n1289));
  OAI22_X1  g1089(.A1(new_n815), .A2(new_n886), .B1(new_n817), .B2(new_n885), .ZN(new_n1290));
  AOI211_X1 g1090(.A(new_n589), .B(new_n1290), .C1(G128), .C2(new_n846), .ZN(new_n1291));
  AOI22_X1  g1091(.A1(G50), .A2(new_n1051), .B1(new_n824), .B2(new_n1212), .ZN(new_n1292));
  AOI22_X1  g1092(.A1(new_n826), .A2(G132), .B1(new_n850), .B2(G159), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1291), .A2(new_n1258), .A3(new_n1292), .A4(new_n1293), .ZN(new_n1294));
  OAI22_X1  g1094(.A1(new_n825), .A2(new_n488), .B1(new_n827), .B2(new_n590), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1295), .B1(G97), .B2(new_n850), .ZN(new_n1296));
  OAI22_X1  g1096(.A1(new_n817), .A2(new_n329), .B1(new_n820), .B2(new_n522), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1297), .B1(G283), .B2(new_n882), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1083), .A2(new_n260), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1296), .A2(new_n1298), .A3(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1294), .B1(new_n1300), .B2(new_n1045), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1289), .B1(new_n1301), .B2(new_n806), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1302), .B1(new_n1192), .B2(new_n892), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1287), .A2(KEYINPUT119), .ZN(new_n1304));
  AND3_X1   g1104(.A1(new_n1288), .A2(new_n1303), .A3(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1285), .A2(new_n1305), .ZN(G381));
  INV_X1    g1106(.A(KEYINPUT120), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n1199), .A2(new_n1307), .A3(new_n1222), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1307), .B1(new_n1199), .B2(new_n1222), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1310), .A2(new_n1253), .A3(new_n1282), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1101), .A2(new_n1129), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1136), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1312), .B1(new_n1313), .B2(new_n1134), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1057), .B1(new_n1012), .B2(new_n1027), .ZN(new_n1315));
  OAI211_X1 g1115(.A(new_n858), .B(new_n1099), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1314), .A2(new_n1315), .A3(new_n899), .A4(new_n1317), .ZN(new_n1318));
  OR3_X1    g1118(.A1(new_n1311), .A2(G381), .A3(new_n1318), .ZN(G407));
  INV_X1    g1119(.A(G343), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(G213), .ZN(new_n1321));
  XNOR2_X1  g1121(.A(new_n1321), .B(KEYINPUT121), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  OAI211_X1 g1123(.A(G407), .B(G213), .C1(new_n1311), .C2(new_n1323), .ZN(G409));
  NAND2_X1  g1124(.A1(G387), .A2(new_n1314), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(G390), .A2(new_n1315), .ZN(new_n1326));
  AOI21_X1  g1126(.A(KEYINPUT122), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n858), .B1(new_n1064), .B2(new_n1099), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1328), .A2(new_n1317), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1329), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1327), .A2(new_n1330), .ZN(new_n1331));
  AOI211_X1 g1131(.A(KEYINPUT122), .B(new_n1329), .C1(new_n1325), .C2(new_n1326), .ZN(new_n1332));
  NOR3_X1   g1132(.A1(new_n1331), .A2(new_n1332), .A3(KEYINPUT61), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1286), .B1(new_n1225), .B2(new_n1011), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1334), .A2(new_n1250), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(new_n1280), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(G378), .A2(KEYINPUT120), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1199), .A2(new_n1307), .A3(new_n1222), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1336), .A2(new_n1337), .A3(new_n1338), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1253), .A2(G378), .A3(new_n1282), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1144), .A2(new_n1154), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT60), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1342), .B1(new_n1172), .B2(new_n1343), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1144), .A2(KEYINPUT60), .A3(new_n1154), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1344), .A2(new_n755), .A3(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1346), .A2(new_n1305), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1347), .A2(new_n899), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1346), .A2(G384), .A3(new_n1305), .ZN(new_n1349));
  AND2_X1   g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  NAND4_X1  g1150(.A1(new_n1341), .A2(KEYINPUT63), .A3(new_n1323), .A4(new_n1350), .ZN(new_n1351));
  AND2_X1   g1151(.A1(new_n1341), .A2(new_n1321), .ZN(new_n1352));
  INV_X1    g1152(.A(G2897), .ZN(new_n1353));
  NOR2_X1   g1153(.A1(new_n1323), .A2(new_n1353), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1354), .B1(new_n1348), .B2(new_n1349), .ZN(new_n1355));
  NOR2_X1   g1155(.A1(new_n1321), .A2(new_n1353), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1355), .B1(new_n1350), .B2(new_n1356), .ZN(new_n1357));
  OAI211_X1 g1157(.A(new_n1333), .B(new_n1351), .C1(new_n1352), .C2(new_n1357), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1281), .B1(new_n1334), .B2(new_n1250), .ZN(new_n1359));
  NOR3_X1   g1159(.A1(new_n1308), .A2(new_n1359), .A3(new_n1309), .ZN(new_n1360));
  AND3_X1   g1160(.A1(new_n1253), .A2(G378), .A3(new_n1282), .ZN(new_n1361));
  OAI211_X1 g1161(.A(new_n1321), .B(new_n1350), .C1(new_n1360), .C2(new_n1361), .ZN(new_n1362));
  INV_X1    g1162(.A(KEYINPUT63), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1362), .A2(new_n1363), .ZN(new_n1364));
  INV_X1    g1164(.A(new_n1364), .ZN(new_n1365));
  OAI21_X1  g1165(.A(KEYINPUT123), .B1(new_n1358), .B2(new_n1365), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1367));
  INV_X1    g1167(.A(KEYINPUT122), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1367), .A2(new_n1368), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1369), .A2(new_n1329), .ZN(new_n1370));
  INV_X1    g1170(.A(KEYINPUT61), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1327), .A2(new_n1330), .ZN(new_n1372));
  NAND3_X1  g1172(.A1(new_n1370), .A2(new_n1371), .A3(new_n1372), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1341), .A2(new_n1321), .ZN(new_n1374));
  INV_X1    g1174(.A(new_n1357), .ZN(new_n1375));
  AOI21_X1  g1175(.A(new_n1373), .B1(new_n1374), .B2(new_n1375), .ZN(new_n1376));
  INV_X1    g1176(.A(KEYINPUT123), .ZN(new_n1377));
  NAND4_X1  g1177(.A1(new_n1376), .A2(new_n1377), .A3(new_n1364), .A4(new_n1351), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1366), .A2(new_n1378), .ZN(new_n1379));
  XNOR2_X1  g1179(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1362), .A2(new_n1380), .ZN(new_n1381));
  AND3_X1   g1181(.A1(new_n1348), .A2(KEYINPUT62), .A3(new_n1349), .ZN(new_n1382));
  OAI211_X1 g1182(.A(new_n1323), .B(new_n1382), .C1(new_n1360), .C2(new_n1361), .ZN(new_n1383));
  INV_X1    g1183(.A(KEYINPUT125), .ZN(new_n1384));
  NAND2_X1  g1184(.A1(new_n1383), .A2(new_n1384), .ZN(new_n1385));
  NAND4_X1  g1185(.A1(new_n1341), .A2(KEYINPUT125), .A3(new_n1323), .A4(new_n1382), .ZN(new_n1386));
  NAND3_X1  g1186(.A1(new_n1381), .A2(new_n1385), .A3(new_n1386), .ZN(new_n1387));
  NAND2_X1  g1187(.A1(new_n1341), .A2(new_n1323), .ZN(new_n1388));
  AOI21_X1  g1188(.A(KEYINPUT61), .B1(new_n1375), .B2(new_n1388), .ZN(new_n1389));
  NAND3_X1  g1189(.A1(new_n1387), .A2(KEYINPUT126), .A3(new_n1389), .ZN(new_n1390));
  NAND2_X1  g1190(.A1(new_n1370), .A2(new_n1372), .ZN(new_n1391));
  NAND2_X1  g1191(.A1(new_n1390), .A2(new_n1391), .ZN(new_n1392));
  AOI21_X1  g1192(.A(KEYINPUT126), .B1(new_n1387), .B2(new_n1389), .ZN(new_n1393));
  OAI21_X1  g1193(.A(new_n1379), .B1(new_n1392), .B2(new_n1393), .ZN(G405));
  AND2_X1   g1194(.A1(new_n1350), .A2(KEYINPUT127), .ZN(new_n1395));
  XOR2_X1   g1195(.A(new_n1391), .B(new_n1395), .Z(new_n1396));
  AOI21_X1  g1196(.A(new_n1361), .B1(new_n1310), .B2(G375), .ZN(new_n1397));
  XNOR2_X1  g1197(.A(new_n1396), .B(new_n1397), .ZN(G402));
endmodule


