//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 0 1 1 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1238, new_n1239, new_n1240, new_n1242, new_n1243,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G13), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT65), .ZN(new_n209));
  INV_X1    g0009(.A(new_n201), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G50), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G1), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n207), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(G13), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT64), .Z(new_n219));
  INV_X1    g0019(.A(KEYINPUT0), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n213), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(new_n220), .B2(new_n219), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT66), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT68), .Z(new_n225));
  INV_X1    g0025(.A(G58), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  INV_X1    g0027(.A(G107), .ZN(new_n228));
  INV_X1    g0028(.A(G264), .ZN(new_n229));
  OAI22_X1  g0029(.A1(new_n226), .A2(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n225), .A2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(KEYINPUT69), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  AOI22_X1  g0034(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT67), .ZN(new_n236));
  AOI22_X1  g0036(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n237));
  OAI211_X1 g0037(.A(new_n236), .B(new_n237), .C1(new_n231), .C2(new_n232), .ZN(new_n238));
  OAI21_X1  g0038(.A(new_n216), .B1(new_n234), .B2(new_n238), .ZN(new_n239));
  NOR2_X1   g0039(.A1(new_n239), .A2(KEYINPUT1), .ZN(new_n240));
  AND2_X1   g0040(.A1(new_n239), .A2(KEYINPUT1), .ZN(new_n241));
  NOR3_X1   g0041(.A1(new_n223), .A2(new_n240), .A3(new_n241), .ZN(G361));
  XNOR2_X1  g0042(.A(G238), .B(G244), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G232), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT2), .B(G226), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G264), .B(G270), .Z(new_n247));
  XNOR2_X1  g0047(.A(G250), .B(G257), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G358));
  XNOR2_X1  g0050(.A(G50), .B(G68), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G58), .B(G77), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n251), .B(new_n252), .Z(new_n253));
  XOR2_X1   g0053(.A(G87), .B(G97), .Z(new_n254));
  XNOR2_X1  g0054(.A(G107), .B(G116), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n253), .B(new_n256), .ZN(G351));
  XNOR2_X1  g0057(.A(KEYINPUT8), .B(G58), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n214), .A2(G13), .A3(G20), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n263));
  AND2_X1   g0063(.A1(new_n263), .A2(new_n206), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n260), .ZN(new_n265));
  OR2_X1    g0065(.A1(new_n265), .A2(KEYINPUT71), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n214), .A2(G20), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(KEYINPUT71), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n262), .B1(new_n269), .B2(new_n259), .ZN(new_n270));
  INV_X1    g0070(.A(G68), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n226), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(G20), .B1(new_n272), .B2(new_n201), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G20), .A2(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G159), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT75), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n277), .B1(new_n278), .B2(KEYINPUT3), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(KEYINPUT3), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT3), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(KEYINPUT75), .A3(G33), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n279), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n207), .ZN(new_n284));
  AND2_X1   g0084(.A1(KEYINPUT76), .A2(KEYINPUT7), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n271), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(KEYINPUT76), .A2(KEYINPUT7), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n283), .A2(new_n288), .A3(new_n207), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n276), .B1(new_n286), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n264), .B1(new_n290), .B2(KEYINPUT16), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT16), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT7), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT3), .B(G33), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n293), .B1(new_n294), .B2(G20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n281), .A2(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n280), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n297), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n271), .B1(new_n295), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n292), .B1(new_n299), .B2(new_n276), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n270), .B1(new_n291), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G41), .ZN(new_n302));
  INV_X1    g0102(.A(G45), .ZN(new_n303));
  AOI21_X1  g0103(.A(G1), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(G33), .A2(G41), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n305), .A2(G1), .A3(G13), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n304), .A2(new_n306), .A3(G274), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n214), .B1(G41), .B2(G45), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n307), .B1(new_n227), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n306), .ZN(new_n311));
  NAND2_X1  g0111(.A1(G33), .A2(G87), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n312), .B(KEYINPUT77), .ZN(new_n313));
  OR2_X1    g0113(.A1(G223), .A2(G1698), .ZN(new_n314));
  INV_X1    g0114(.A(G1698), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n314), .B1(G226), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n313), .B1(new_n283), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n310), .B1(new_n311), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G169), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n320), .B1(G179), .B2(new_n318), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT18), .B1(new_n301), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n270), .ZN(new_n323));
  INV_X1    g0123(.A(G200), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n317), .A2(new_n311), .ZN(new_n325));
  INV_X1    g0125(.A(new_n310), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n327), .B1(G190), .B2(new_n318), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n284), .A2(new_n285), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n329), .A2(G68), .A3(new_n289), .ZN(new_n330));
  INV_X1    g0130(.A(new_n276), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n330), .A2(KEYINPUT16), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n263), .A2(new_n206), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n332), .A2(new_n300), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n323), .A2(new_n328), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT17), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n301), .A2(KEYINPUT17), .A3(new_n328), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n323), .A2(new_n334), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n318), .A2(G179), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(new_n319), .B2(new_n318), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT18), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n339), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n322), .A2(new_n337), .A3(new_n338), .A4(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n227), .A2(G1698), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n294), .B(new_n346), .C1(G226), .C2(G1698), .ZN(new_n347));
  NAND2_X1  g0147(.A1(G33), .A2(G97), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n306), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G238), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n307), .B1(new_n351), .B2(new_n309), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT13), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n350), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT13), .B1(new_n349), .B2(new_n352), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G169), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT14), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT14), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n357), .A2(new_n360), .A3(G169), .ZN(new_n361));
  INV_X1    g0161(.A(G179), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n359), .B(new_n361), .C1(new_n362), .C2(new_n357), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n274), .A2(G50), .B1(G20), .B2(new_n271), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n207), .A2(G33), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT70), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n365), .B(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G77), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n364), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n369), .A2(KEYINPUT11), .A3(new_n333), .ZN(new_n370));
  OR3_X1    g0170(.A1(new_n260), .A2(KEYINPUT12), .A3(G68), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT12), .B1(new_n260), .B2(G68), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n267), .A2(G68), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n370), .B(new_n373), .C1(new_n265), .C2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT11), .B1(new_n369), .B2(new_n333), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n363), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G190), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n377), .B1(new_n380), .B2(new_n357), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n357), .A2(G200), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT74), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n357), .A2(KEYINPUT74), .A3(G200), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n381), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n379), .A2(new_n386), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n274), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n367), .B2(new_n258), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n389), .A2(new_n333), .B1(new_n202), .B2(new_n261), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n202), .B2(new_n269), .ZN(new_n391));
  INV_X1    g0191(.A(new_n307), .ZN(new_n392));
  INV_X1    g0192(.A(new_n309), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n392), .B1(G226), .B2(new_n393), .ZN(new_n394));
  NOR2_X1   g0194(.A1(G222), .A2(G1698), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n315), .A2(G223), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n294), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n397), .B(new_n311), .C1(G77), .C2(new_n294), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n319), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n394), .A2(new_n362), .A3(new_n398), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n391), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n399), .A2(new_n380), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n404), .B1(G200), .B2(new_n399), .ZN(new_n405));
  AND2_X1   g0205(.A1(new_n391), .A2(KEYINPUT9), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n391), .A2(KEYINPUT9), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OR2_X1    g0208(.A1(new_n408), .A2(KEYINPUT10), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(KEYINPUT10), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n403), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n259), .A2(new_n274), .B1(G20), .B2(G77), .ZN(new_n412));
  XNOR2_X1  g0212(.A(KEYINPUT15), .B(G87), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n412), .B1(new_n365), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n333), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n264), .A2(G77), .A3(new_n260), .A4(new_n267), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT73), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n260), .A2(G77), .ZN(new_n418));
  XNOR2_X1  g0218(.A(new_n418), .B(KEYINPUT72), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n415), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(G244), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n307), .B1(new_n421), .B2(new_n309), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n294), .A2(G238), .A3(G1698), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n294), .A2(G232), .A3(new_n315), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n423), .B(new_n424), .C1(new_n228), .C2(new_n294), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n422), .B1(new_n425), .B2(new_n311), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n362), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n420), .B(new_n427), .C1(G169), .C2(new_n426), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  OR2_X1    g0229(.A1(new_n426), .A2(new_n324), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n420), .B1(G190), .B2(new_n426), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AND4_X1   g0232(.A1(new_n345), .A2(new_n387), .A3(new_n411), .A4(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT82), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n274), .A2(G77), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n228), .A2(KEYINPUT6), .A3(G97), .ZN(new_n437));
  XNOR2_X1  g0237(.A(G97), .B(G107), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT6), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n436), .B1(new_n440), .B2(new_n207), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n228), .B1(new_n295), .B2(new_n298), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n441), .B1(KEYINPUT78), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(KEYINPUT7), .B1(new_n297), .B2(new_n207), .ZN(new_n444));
  AOI211_X1 g0244(.A(new_n293), .B(G20), .C1(new_n280), .C2(new_n296), .ZN(new_n445));
  OAI21_X1  g0245(.A(G107), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT78), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n264), .B1(new_n443), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n260), .A2(G97), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n214), .A2(G33), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n264), .A2(new_n260), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n450), .B1(new_n452), .B2(G97), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(G283), .ZN(new_n456));
  OAI21_X1  g0256(.A(KEYINPUT80), .B1(new_n278), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT80), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n458), .A2(G33), .A3(G283), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n280), .A2(new_n296), .A3(G250), .A4(G1698), .ZN(new_n461));
  AND2_X1   g0261(.A1(KEYINPUT4), .A2(G244), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n280), .A2(new_n296), .A3(new_n462), .A4(new_n315), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n460), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT4), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n421), .A2(G1698), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n465), .B1(new_n283), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n306), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT5), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT81), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n470), .B1(new_n471), .B2(G41), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n302), .A2(KEYINPUT81), .A3(KEYINPUT5), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n303), .A2(G1), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n306), .A2(G274), .ZN(new_n476));
  OR2_X1    g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G257), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n475), .A2(new_n306), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n469), .A2(new_n480), .A3(new_n362), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n279), .A2(new_n280), .A3(new_n282), .ZN(new_n482));
  AOI21_X1  g0282(.A(KEYINPUT4), .B1(new_n482), .B2(new_n466), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n461), .A2(new_n460), .A3(new_n463), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n311), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n475), .A2(new_n476), .ZN(new_n486));
  INV_X1    g0286(.A(new_n479), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n486), .B1(new_n487), .B2(G257), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n319), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n481), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n435), .B1(new_n455), .B2(new_n490), .ZN(new_n491));
  OAI211_X1 g0291(.A(KEYINPUT78), .B(G107), .C1(new_n444), .C2(new_n445), .ZN(new_n492));
  INV_X1    g0292(.A(new_n436), .ZN(new_n493));
  INV_X1    g0293(.A(G97), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n494), .A2(new_n228), .ZN(new_n495));
  NOR2_X1   g0295(.A1(G97), .A2(G107), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n439), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n437), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n493), .B1(new_n499), .B2(G20), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n492), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n442), .A2(KEYINPUT78), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n333), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n453), .ZN(new_n504));
  OAI21_X1  g0304(.A(G169), .B1(new_n469), .B2(new_n480), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n485), .A2(new_n488), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n505), .B1(new_n506), .B2(new_n362), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n504), .A2(new_n507), .A3(KEYINPUT82), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n491), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n279), .A2(new_n282), .A3(new_n207), .A4(new_n280), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n365), .A2(new_n494), .ZN(new_n511));
  OAI22_X1  g0311(.A1(new_n510), .A2(new_n271), .B1(KEYINPUT19), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT83), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n513), .A2(new_n514), .A3(new_n207), .ZN(new_n515));
  INV_X1    g0315(.A(G87), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n496), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n514), .B1(new_n513), .B2(new_n207), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n333), .B1(new_n512), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n413), .A2(new_n261), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n421), .A2(G1698), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(G238), .B2(G1698), .ZN(new_n525));
  INV_X1    g0325(.A(G116), .ZN(new_n526));
  OAI22_X1  g0326(.A1(new_n283), .A2(new_n525), .B1(new_n278), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n311), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n214), .A2(G45), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n306), .A2(G250), .A3(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n476), .B2(new_n529), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(G200), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n452), .A2(G87), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n531), .B1(new_n527), .B2(new_n311), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G190), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n523), .A2(new_n534), .A3(new_n535), .A4(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n264), .A2(new_n260), .A3(new_n451), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n521), .B(new_n522), .C1(new_n413), .C2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n533), .A2(new_n319), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n536), .A2(new_n362), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n538), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(KEYINPUT22), .A2(G87), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n510), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT24), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT22), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n207), .A2(G87), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n549), .B1(new_n297), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT23), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n207), .B2(G107), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n228), .A2(KEYINPUT23), .A3(G20), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n278), .A2(new_n526), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n553), .A2(new_n554), .B1(new_n555), .B2(new_n207), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n547), .A2(new_n548), .A3(new_n551), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n551), .A2(new_n556), .ZN(new_n558));
  OAI21_X1  g0358(.A(KEYINPUT24), .B1(new_n558), .B2(new_n546), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n264), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT25), .ZN(new_n561));
  NOR3_X1   g0361(.A1(new_n260), .A2(new_n561), .A3(G107), .ZN(new_n562));
  AOI21_X1  g0362(.A(KEYINPUT25), .B1(new_n261), .B2(new_n228), .ZN(new_n563));
  OAI22_X1  g0363(.A1(new_n562), .A2(new_n563), .B1(new_n228), .B2(new_n539), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n478), .A2(G1698), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(G250), .B2(G1698), .ZN(new_n567));
  INV_X1    g0367(.A(G294), .ZN(new_n568));
  OAI22_X1  g0368(.A1(new_n283), .A2(new_n567), .B1(new_n278), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n311), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n570), .B(new_n477), .C1(new_n229), .C2(new_n479), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n324), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(G190), .B2(new_n571), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n544), .B1(new_n565), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(KEYINPUT79), .B1(new_n449), .B2(new_n454), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n506), .A2(new_n324), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(G190), .B2(new_n506), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT79), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n503), .A2(new_n578), .A3(new_n453), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n575), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n509), .A2(new_n574), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT86), .ZN(new_n582));
  AOI21_X1  g0382(.A(G20), .B1(new_n278), .B2(G97), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n460), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT85), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n526), .A2(G20), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n333), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n585), .B1(new_n333), .B2(new_n586), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n584), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT20), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n584), .B(KEYINPUT20), .C1(new_n587), .C2(new_n588), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n452), .A2(KEYINPUT84), .A3(G116), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT84), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n539), .B2(new_n526), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n594), .A2(new_n596), .B1(new_n526), .B2(new_n261), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(G257), .A2(G1698), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n229), .B2(G1698), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n482), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n297), .A2(G303), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n306), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(G270), .ZN(new_n604));
  OAI22_X1  g0404(.A1(new_n479), .A2(new_n604), .B1(new_n476), .B2(new_n475), .ZN(new_n605));
  OAI21_X1  g0405(.A(G200), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n582), .B1(new_n598), .B2(new_n606), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n606), .A2(new_n593), .A3(new_n597), .A4(new_n582), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n603), .A2(new_n605), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(G190), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT21), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n601), .A2(new_n602), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n311), .ZN(new_n615));
  INV_X1    g0415(.A(new_n605), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(G169), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n613), .B1(new_n598), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n593), .A2(new_n597), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n603), .A2(new_n605), .A3(new_n362), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n620), .A2(KEYINPUT21), .A3(G169), .A4(new_n617), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n571), .A2(new_n319), .ZN(new_n624));
  AOI22_X1  g0424(.A1(G264), .A2(new_n487), .B1(new_n569), .B2(new_n311), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n625), .A2(new_n362), .A3(new_n477), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n624), .B(new_n626), .C1(new_n560), .C2(new_n564), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n619), .A2(new_n622), .A3(new_n623), .A4(new_n627), .ZN(new_n628));
  NOR4_X1   g0428(.A1(new_n434), .A2(new_n581), .A3(new_n612), .A4(new_n628), .ZN(G372));
  NAND2_X1  g0429(.A1(new_n337), .A2(new_n338), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n386), .A2(new_n428), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n631), .B1(new_n632), .B2(new_n379), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT89), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n301), .A2(KEYINPUT18), .A3(new_n321), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n342), .B1(new_n339), .B2(new_n341), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n322), .A2(KEYINPUT89), .A3(new_n343), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n633), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n409), .A2(new_n410), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n403), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n503), .A2(new_n578), .A3(new_n453), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n578), .B1(new_n503), .B2(new_n453), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n507), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT88), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT26), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n538), .A2(new_n543), .ZN(new_n649));
  OAI211_X1 g0449(.A(KEYINPUT88), .B(new_n507), .C1(new_n643), .C2(new_n644), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n647), .A2(new_n648), .A3(new_n649), .A4(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n543), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n491), .A2(new_n508), .A3(new_n649), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n652), .B1(new_n653), .B2(KEYINPUT26), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n628), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(new_n581), .B2(KEYINPUT87), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT87), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n509), .A2(new_n574), .A3(new_n658), .A4(new_n580), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n655), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n642), .B1(new_n434), .B2(new_n660), .ZN(G369));
  INV_X1    g0461(.A(G13), .ZN(new_n662));
  NOR3_X1   g0462(.A1(new_n662), .A2(G1), .A3(G20), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT90), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT27), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(G213), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n664), .A2(new_n665), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(G343), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n620), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT91), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n623), .A2(new_n622), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n619), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n674), .A2(new_n612), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n677), .B1(new_n678), .B2(new_n676), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(G330), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n627), .ZN(new_n682));
  OAI211_X1 g0482(.A(G343), .B(new_n669), .C1(new_n560), .C2(new_n564), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n573), .A2(new_n565), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n682), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n627), .A2(new_n672), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n672), .B1(new_n675), .B2(new_n619), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n686), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(G399));
  INV_X1    g0491(.A(new_n217), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n517), .A2(G116), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G1), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n211), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  INV_X1    g0498(.A(new_n672), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n509), .A2(new_n574), .A3(new_n580), .A4(new_n628), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n491), .A2(new_n649), .A3(new_n648), .A4(new_n508), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(new_n543), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n544), .B1(new_n645), .B2(new_n646), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n648), .B1(new_n703), .B2(new_n650), .ZN(new_n704));
  OAI211_X1 g0504(.A(KEYINPUT29), .B(new_n699), .C1(new_n702), .C2(new_n704), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n651), .A2(new_n654), .ZN(new_n706));
  AND3_X1   g0506(.A1(new_n504), .A2(new_n507), .A3(KEYINPUT82), .ZN(new_n707));
  AOI21_X1  g0507(.A(KEYINPUT82), .B1(new_n504), .B2(new_n507), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n580), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n649), .A2(new_n684), .ZN(new_n710));
  OAI21_X1  g0510(.A(KEYINPUT87), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n711), .A2(new_n628), .A3(new_n659), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n672), .B1(new_n706), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n705), .B1(new_n713), .B2(KEYINPUT29), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n643), .A2(new_n644), .ZN(new_n715));
  AOI22_X1  g0515(.A1(new_n715), .A2(new_n577), .B1(new_n491), .B2(new_n508), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n628), .A2(new_n612), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n716), .A2(new_n717), .A3(new_n574), .A4(new_n699), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT31), .ZN(new_n719));
  INV_X1    g0519(.A(new_n621), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n625), .A2(new_n485), .A3(new_n488), .A4(new_n536), .ZN(new_n721));
  OAI21_X1  g0521(.A(KEYINPUT30), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n625), .A2(new_n536), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT30), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n469), .A2(new_n480), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n723), .A2(new_n724), .A3(new_n725), .A4(new_n621), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n609), .A2(G179), .A3(new_n536), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n506), .A2(new_n571), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n722), .A2(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT92), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n672), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n722), .A2(new_n726), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n728), .A2(new_n727), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n732), .A2(new_n730), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n719), .B1(new_n731), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n732), .A2(new_n733), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n736), .A2(KEYINPUT31), .A3(new_n672), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n718), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G330), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n714), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n698), .B1(new_n740), .B2(G1), .ZN(G364));
  NOR2_X1   g0541(.A1(new_n662), .A2(G20), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n214), .B1(new_n742), .B2(G45), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n693), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n681), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(G330), .B2(new_n679), .ZN(new_n747));
  INV_X1    g0547(.A(new_n745), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n206), .B1(G20), .B2(new_n319), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n380), .A2(G20), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT95), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n753), .A2(G179), .A3(G200), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n755), .A2(KEYINPUT96), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(KEYINPUT96), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G159), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT32), .ZN(new_n761));
  NAND2_X1  g0561(.A1(G20), .A2(G179), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n762), .A2(new_n380), .A3(G200), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n762), .A2(G190), .A3(G200), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n764), .A2(new_n226), .B1(new_n766), .B2(new_n368), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n762), .A2(new_n324), .A3(G190), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n767), .B1(G68), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n762), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(G190), .A3(G200), .ZN(new_n771));
  OAI21_X1  g0571(.A(G20), .B1(G179), .B2(G200), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n751), .A2(new_n772), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n773), .A2(KEYINPUT98), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(KEYINPUT98), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n769), .B1(new_n202), .B2(new_n771), .C1(new_n494), .C2(new_n776), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n753), .A2(G179), .A3(new_n324), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G107), .ZN(new_n779));
  NOR4_X1   g0579(.A1(new_n207), .A2(new_n380), .A3(new_n324), .A4(G179), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI211_X1 g0581(.A(new_n779), .B(new_n294), .C1(new_n516), .C2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n777), .B1(KEYINPUT97), .B2(new_n782), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n761), .B(new_n783), .C1(KEYINPUT97), .C2(new_n782), .ZN(new_n784));
  INV_X1    g0584(.A(new_n758), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G329), .ZN(new_n786));
  INV_X1    g0586(.A(new_n776), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G294), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n778), .A2(G283), .ZN(new_n789));
  INV_X1    g0589(.A(G303), .ZN(new_n790));
  INV_X1    g0590(.A(G311), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n781), .A2(new_n790), .B1(new_n791), .B2(new_n766), .ZN(new_n792));
  INV_X1    g0592(.A(G322), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n297), .B1(new_n764), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n768), .ZN(new_n795));
  XOR2_X1   g0595(.A(KEYINPUT33), .B(G317), .Z(new_n796));
  INV_X1    g0596(.A(G326), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n795), .A2(new_n796), .B1(new_n771), .B2(new_n797), .ZN(new_n798));
  NOR3_X1   g0598(.A1(new_n792), .A2(new_n794), .A3(new_n798), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n786), .A2(new_n788), .A3(new_n789), .A4(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n750), .B1(new_n784), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(G13), .A2(G33), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(G20), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n749), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n692), .A2(new_n297), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n806), .A2(G355), .B1(new_n526), .B2(new_n692), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n253), .A2(new_n303), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT93), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n692), .A2(new_n482), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(new_n303), .B2(new_n212), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(KEYINPUT94), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n812), .A2(KEYINPUT94), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n807), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n748), .B(new_n801), .C1(new_n805), .C2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n804), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n679), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n747), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(G396));
  NAND2_X1  g0621(.A1(new_n429), .A2(new_n699), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n431), .A2(new_n430), .B1(new_n672), .B2(new_n420), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n823), .B2(new_n429), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n713), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n432), .A2(new_n699), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(new_n706), .B2(new_n712), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n739), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n745), .B1(new_n829), .B2(new_n830), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n831), .B1(new_n832), .B2(KEYINPUT100), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(KEYINPUT100), .B2(new_n832), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n778), .A2(G68), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n835), .B(new_n482), .C1(new_n202), .C2(new_n781), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(G58), .B2(new_n787), .ZN(new_n837));
  INV_X1    g0637(.A(G132), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n837), .B1(new_n838), .B2(new_n758), .ZN(new_n839));
  AOI22_X1  g0639(.A1(G143), .A2(new_n763), .B1(new_n765), .B2(G159), .ZN(new_n840));
  INV_X1    g0640(.A(G137), .ZN(new_n841));
  INV_X1    g0641(.A(G150), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n840), .B1(new_n841), .B2(new_n771), .C1(new_n842), .C2(new_n795), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT34), .Z(new_n844));
  AOI22_X1  g0644(.A1(G116), .A2(new_n765), .B1(new_n763), .B2(G294), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n845), .B1(new_n456), .B2(new_n795), .C1(new_n790), .C2(new_n771), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(G97), .B2(new_n787), .ZN(new_n847));
  INV_X1    g0647(.A(new_n778), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n848), .A2(new_n516), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n297), .B1(new_n781), .B2(new_n228), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n849), .B1(KEYINPUT99), .B2(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n847), .B(new_n851), .C1(KEYINPUT99), .C2(new_n850), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n758), .A2(new_n791), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n839), .A2(new_n844), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n749), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n749), .A2(new_n802), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n748), .B1(new_n368), .B2(new_n856), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n855), .B(new_n857), .C1(new_n825), .C2(new_n803), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n834), .A2(new_n858), .ZN(G384));
  NOR2_X1   g0659(.A1(new_n742), .A2(new_n214), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n339), .A2(new_n341), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n339), .A2(new_n669), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n861), .A2(new_n862), .A3(new_n335), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT37), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT37), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n861), .A2(new_n862), .A3(new_n865), .A4(new_n335), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n630), .B1(new_n637), .B2(new_n638), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n867), .B1(new_n868), .B2(new_n862), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT38), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n330), .A2(new_n331), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n292), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n270), .B1(new_n291), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n335), .B1(new_n874), .B2(new_n321), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n874), .A2(new_n670), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT37), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n866), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n344), .A2(new_n876), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n878), .A2(new_n879), .A3(KEYINPUT38), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n871), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n736), .A2(KEYINPUT92), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n729), .A2(new_n730), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n882), .A2(KEYINPUT31), .A3(new_n672), .A4(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n718), .A2(new_n735), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n363), .A2(new_n378), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n384), .A2(new_n385), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n887), .B(new_n377), .C1(new_n380), .C2(new_n357), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n378), .A2(new_n672), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n886), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n378), .B(new_n672), .C1(new_n386), .C2(new_n363), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n824), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n885), .A2(new_n892), .A3(KEYINPUT40), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n878), .A2(new_n879), .A3(KEYINPUT38), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT38), .B1(new_n878), .B2(new_n879), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n885), .B(new_n892), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT40), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n881), .A2(new_n893), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n898), .B(KEYINPUT101), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n433), .A2(new_n885), .ZN(new_n900));
  OR2_X1    g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n900), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n901), .A2(G330), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n878), .A2(new_n879), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n870), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n880), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n890), .A2(new_n891), .ZN(new_n907));
  INV_X1    g0707(.A(new_n822), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n906), .B(new_n907), .C1(new_n828), .C2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n637), .A2(new_n638), .A3(new_n670), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n379), .A2(new_n699), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT39), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n880), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n871), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT39), .B1(new_n894), .B2(new_n895), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n912), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n911), .A2(new_n918), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n433), .B(new_n705), .C1(new_n713), .C2(KEYINPUT29), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n642), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n919), .B(new_n921), .Z(new_n922));
  AOI21_X1  g0722(.A(new_n860), .B1(new_n903), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n922), .B2(new_n903), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n499), .A2(KEYINPUT35), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n499), .A2(KEYINPUT35), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n925), .A2(G116), .A3(new_n209), .A4(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT36), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n211), .A2(new_n368), .A3(new_n272), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n271), .A2(G50), .ZN(new_n930));
  OAI211_X1 g0730(.A(G1), .B(new_n662), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n924), .A2(new_n928), .A3(new_n931), .ZN(G367));
  OAI221_X1 g0732(.A(new_n805), .B1(new_n217), .B2(new_n413), .C1(new_n811), .C2(new_n249), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n933), .A2(new_n745), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n523), .A2(new_n535), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n672), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n649), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n652), .A2(new_n935), .A3(new_n672), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT46), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n781), .A2(new_n940), .A3(new_n526), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n940), .B1(new_n781), .B2(new_n526), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n791), .B2(new_n771), .ZN(new_n943));
  AOI211_X1 g0743(.A(new_n941), .B(new_n943), .C1(G294), .C2(new_n768), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n848), .A2(new_n494), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n764), .A2(new_n790), .B1(new_n766), .B2(new_n456), .ZN(new_n946));
  NOR3_X1   g0746(.A1(new_n945), .A2(new_n482), .A3(new_n946), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n944), .B(new_n947), .C1(new_n228), .C2(new_n776), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(G317), .B2(new_n785), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n776), .A2(new_n271), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n778), .A2(G77), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n297), .B1(new_n780), .B2(G58), .ZN(new_n952));
  AOI22_X1  g0752(.A1(G50), .A2(new_n765), .B1(new_n763), .B2(G150), .ZN(new_n953));
  INV_X1    g0753(.A(new_n771), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n954), .A2(G143), .B1(G159), .B2(new_n768), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n951), .A2(new_n952), .A3(new_n953), .A4(new_n955), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n950), .B(new_n956), .C1(new_n785), .C2(G137), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n949), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT47), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n934), .B1(new_n818), .B2(new_n939), .C1(new_n959), .C2(new_n750), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n645), .A2(new_n699), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n672), .B1(new_n643), .B2(new_n644), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n961), .B1(new_n716), .B2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT103), .ZN(new_n965));
  AND3_X1   g0765(.A1(new_n964), .A2(new_n965), .A3(new_n690), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n965), .B1(new_n964), .B2(new_n690), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT45), .ZN(new_n968));
  OR3_X1    g0768(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n964), .A2(new_n690), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT44), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n968), .B1(new_n966), .B2(new_n967), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n969), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n688), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n687), .B(new_n689), .Z(new_n976));
  INV_X1    g0776(.A(KEYINPUT104), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n976), .B1(new_n681), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n680), .B(KEYINPUT104), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n978), .B1(new_n979), .B2(new_n976), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n969), .A2(new_n971), .A3(new_n688), .A4(new_n972), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n975), .A2(new_n980), .A3(new_n740), .A4(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n740), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n693), .B(KEYINPUT41), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n744), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n687), .A2(new_n689), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n964), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(KEYINPUT42), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT102), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n509), .B1(new_n963), .B2(new_n627), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n699), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n988), .A2(new_n989), .A3(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(KEYINPUT42), .B2(new_n987), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n989), .B1(new_n988), .B2(new_n991), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT43), .ZN(new_n996));
  INV_X1    g0796(.A(new_n939), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n996), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n999), .B(new_n1000), .C1(new_n993), .C2(new_n994), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n688), .A2(new_n963), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n998), .A2(new_n1003), .A3(new_n1001), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n960), .B1(new_n985), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT105), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g0810(.A(KEYINPUT105), .B(new_n960), .C1(new_n985), .C2(new_n1007), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(G387));
  OAI211_X1 g0812(.A(new_n695), .B(new_n303), .C1(new_n271), .C2(new_n368), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(KEYINPUT106), .ZN(new_n1014));
  OAI21_X1  g0814(.A(KEYINPUT50), .B1(new_n258), .B2(G50), .ZN(new_n1015));
  OR3_X1    g0815(.A1(new_n258), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1013), .A2(KEYINPUT106), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n810), .B1(new_n1017), .B2(new_n1018), .C1(new_n246), .C2(new_n303), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n806), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1019), .B1(G107), .B2(new_n217), .C1(new_n695), .C2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n748), .B1(new_n1021), .B2(new_n805), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n687), .B2(new_n818), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n785), .A2(G150), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n781), .A2(new_n368), .B1(new_n202), .B2(new_n764), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1025), .B(new_n945), .C1(G68), .C2(new_n765), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n413), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n787), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n482), .B1(new_n258), .B2(new_n795), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(G159), .B2(new_n954), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1024), .A2(new_n1026), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n787), .A2(G283), .B1(G294), .B2(new_n780), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT48), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(G303), .A2(new_n765), .B1(new_n763), .B2(G317), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n791), .B2(new_n795), .C1(new_n793), .C2(new_n771), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1032), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT107), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(new_n1033), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1037), .A2(KEYINPUT49), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n482), .B1(new_n778), .B2(G116), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(new_n797), .C2(new_n758), .ZN(new_n1041));
  AOI21_X1  g0841(.A(KEYINPUT49), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1031), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1023), .B1(new_n1043), .B2(new_n749), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n980), .B2(new_n744), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n980), .A2(new_n740), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n693), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n980), .A2(new_n740), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1045), .B1(new_n1047), .B2(new_n1048), .ZN(G393));
  NAND2_X1  g0849(.A1(new_n975), .A2(new_n981), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n963), .A2(new_n804), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n805), .B1(new_n494), .B2(new_n217), .C1(new_n811), .C2(new_n256), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G294), .A2(new_n765), .B1(new_n768), .B2(G303), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n776), .B2(new_n526), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT108), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n954), .A2(G317), .B1(G311), .B2(new_n763), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT52), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n779), .B(new_n297), .C1(new_n456), .C2(new_n781), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1058), .B(new_n1059), .C1(new_n785), .C2(G322), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n780), .A2(G68), .B1(new_n259), .B2(new_n765), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1061), .B(new_n482), .C1(new_n202), .C2(new_n795), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n849), .B(new_n1062), .C1(new_n785), .C2(G143), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n787), .A2(G77), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n764), .A2(new_n759), .B1(new_n771), .B2(new_n842), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT51), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1068));
  AND3_X1   g0868(.A1(new_n1064), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1056), .A2(new_n1060), .B1(new_n1063), .B2(new_n1069), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n745), .B(new_n1053), .C1(new_n1070), .C2(new_n750), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT109), .Z(new_n1072));
  AOI22_X1  g0872(.A1(new_n1051), .A2(new_n744), .B1(new_n1052), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1050), .A2(new_n1046), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1074), .A2(new_n982), .A3(new_n693), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1073), .A2(new_n1075), .ZN(G390));
  NAND3_X1  g0876(.A1(new_n433), .A2(G330), .A3(new_n885), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n920), .A2(new_n642), .A3(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n738), .A2(G330), .A3(new_n825), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n907), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n885), .A2(new_n892), .A3(G330), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n822), .B1(new_n660), .B2(new_n827), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n823), .A2(new_n429), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n699), .B(new_n1086), .C1(new_n702), .C2(new_n704), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n1087), .A2(new_n822), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n738), .A2(G330), .A3(new_n825), .A4(new_n907), .ZN(new_n1089));
  AND3_X1   g0889(.A1(new_n885), .A2(G330), .A3(new_n825), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1088), .B(new_n1089), .C1(new_n907), .C2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1078), .B1(new_n1085), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT111), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1092), .B(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1082), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n322), .A2(KEYINPUT89), .A3(new_n343), .ZN(new_n1096));
  AOI21_X1  g0896(.A(KEYINPUT89), .B1(new_n322), .B2(new_n343), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n631), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n862), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(KEYINPUT38), .B1(new_n1100), .B2(new_n867), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n917), .B1(new_n1101), .B2(new_n914), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n907), .B1(new_n828), .B2(new_n908), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1102), .B1(new_n912), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n881), .A2(new_n912), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1080), .B1(new_n1087), .B2(new_n822), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1095), .B1(new_n1104), .B2(new_n1107), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n912), .B(new_n881), .C1(new_n1088), .C2(new_n1080), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n912), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n1084), .B2(new_n907), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1109), .B(new_n1089), .C1(new_n1111), .C2(new_n1102), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1108), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1094), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1108), .A2(new_n1092), .A3(new_n1112), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT110), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1108), .A2(new_n1092), .A3(new_n1112), .A4(KEYINPUT110), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1114), .A2(new_n1119), .A3(new_n693), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT114), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1108), .A2(new_n744), .A3(new_n1112), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(KEYINPUT112), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT112), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1108), .A2(new_n1112), .A3(new_n1124), .A4(new_n744), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n780), .A2(G150), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT113), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT53), .ZN(new_n1129));
  INV_X1    g0929(.A(G125), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1129), .B1(new_n758), .B2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT54), .B(G143), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n294), .B1(new_n766), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(G128), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n795), .A2(new_n841), .B1(new_n771), .B2(new_n1134), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1133), .B(new_n1135), .C1(G132), .C2(new_n763), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n1136), .B1(new_n202), .B2(new_n848), .C1(new_n759), .C2(new_n776), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n758), .A2(new_n568), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n764), .A2(new_n526), .B1(new_n766), .B2(new_n494), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n294), .B(new_n1139), .C1(G87), .C2(new_n780), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n954), .A2(G283), .B1(G107), .B2(new_n768), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1140), .A2(new_n835), .A3(new_n1064), .A4(new_n1141), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n1131), .A2(new_n1137), .B1(new_n1138), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n749), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n748), .B1(new_n258), .B2(new_n856), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1144), .B(new_n1145), .C1(new_n1102), .C2(new_n803), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1121), .B1(new_n1126), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1146), .ZN(new_n1148));
  AOI211_X1 g0948(.A(KEYINPUT114), .B(new_n1148), .C1(new_n1123), .C2(new_n1125), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1120), .B1(new_n1147), .B2(new_n1149), .ZN(G378));
  NAND2_X1  g0950(.A1(new_n881), .A2(new_n893), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n896), .A2(new_n897), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1151), .A2(new_n1152), .A3(G330), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n391), .A2(new_n669), .ZN(new_n1154));
  OR2_X1    g0954(.A1(new_n411), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n411), .A2(new_n1154), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1155), .A2(new_n1156), .A3(new_n1158), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1153), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n898), .A2(G330), .A3(new_n1162), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1164), .A2(new_n919), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n919), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1078), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1168), .B1(new_n1119), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(KEYINPUT118), .B1(new_n1170), .B2(KEYINPUT57), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n694), .B1(new_n1170), .B2(KEYINPUT57), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT118), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT57), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1078), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1173), .B(new_n1174), .C1(new_n1175), .C2(new_n1168), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1171), .A2(new_n1172), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1163), .A2(new_n802), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n856), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n745), .B1(G50), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n778), .A2(G58), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT115), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n758), .B2(new_n456), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n1027), .A2(new_n765), .B1(new_n763), .B2(G107), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1184), .B(new_n302), .C1(new_n368), .C2(new_n781), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n283), .B1(new_n771), .B2(new_n526), .C1(new_n795), .C2(new_n494), .ZN(new_n1186));
  NOR4_X1   g0986(.A1(new_n1183), .A2(new_n950), .A3(new_n1185), .A4(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n302), .B1(new_n283), .B2(new_n278), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n1187), .A2(KEYINPUT58), .B1(new_n202), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1132), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n780), .A2(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT117), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n954), .A2(G125), .B1(G128), .B2(new_n763), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1192), .B(new_n1193), .C1(new_n842), .C2(new_n776), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(G132), .A2(new_n768), .B1(new_n765), .B2(G137), .ZN(new_n1195));
  XOR2_X1   g0995(.A(new_n1195), .B(KEYINPUT116), .Z(new_n1196));
  NOR2_X1   g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1198), .A2(KEYINPUT59), .ZN(new_n1199));
  AOI211_X1 g0999(.A(G33), .B(G41), .C1(new_n778), .C2(G159), .ZN(new_n1200));
  INV_X1    g1000(.A(G124), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT59), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1200), .B1(new_n1201), .B2(new_n758), .C1(new_n1197), .C2(new_n1202), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1189), .B1(KEYINPUT58), .B2(new_n1187), .C1(new_n1199), .C2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1180), .B1(new_n1204), .B2(new_n749), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1178), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n919), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1164), .A2(new_n919), .A3(new_n1165), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1207), .B1(new_n1212), .B2(new_n744), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1177), .A2(new_n1213), .ZN(G375));
  AND2_X1   g1014(.A1(new_n1085), .A2(new_n1091), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n1078), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1094), .A2(new_n984), .A3(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1215), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1080), .A2(new_n802), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n745), .B1(G68), .B2(new_n1179), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n297), .B1(new_n456), .B2(new_n764), .C1(new_n781), .C2(new_n494), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(G77), .B2(new_n778), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1222), .B(new_n1028), .C1(new_n758), .C2(new_n790), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n954), .A2(G294), .B1(G107), .B2(new_n765), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n526), .B2(new_n795), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1225), .B(KEYINPUT119), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1182), .B1(new_n758), .B2(new_n1134), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n781), .A2(new_n759), .B1(new_n841), .B2(new_n764), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G150), .B2(new_n765), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n787), .A2(G50), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n954), .A2(G132), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n283), .B1(new_n768), .B2(new_n1190), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n1223), .A2(new_n1226), .B1(new_n1227), .B2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1220), .B1(new_n1234), .B2(new_n749), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1218), .A2(new_n744), .B1(new_n1219), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1217), .A2(new_n1236), .ZN(G381));
  XNOR2_X1  g1037(.A(G375), .B(KEYINPUT120), .ZN(new_n1238));
  OR4_X1    g1038(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1239));
  OR4_X1    g1039(.A1(G387), .A2(new_n1239), .A3(G378), .A4(G381), .ZN(new_n1240));
  OR2_X1    g1040(.A1(new_n1238), .A2(new_n1240), .ZN(G407));
  NAND2_X1  g1041(.A1(new_n671), .A2(G213), .ZN(new_n1242));
  OR2_X1    g1042(.A1(G378), .A2(new_n1242), .ZN(new_n1243));
  OAI211_X1 g1043(.A(G407), .B(G213), .C1(new_n1238), .C2(new_n1243), .ZN(G409));
  OAI21_X1  g1044(.A(KEYINPUT60), .B1(new_n1215), .B2(new_n1078), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1245), .A2(new_n1216), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n693), .B1(new_n1245), .B2(new_n1216), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1236), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(G384), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  OAI211_X1 g1050(.A(G384), .B(new_n1236), .C1(new_n1246), .C2(new_n1247), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n1250), .A2(KEYINPUT123), .A3(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(KEYINPUT123), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1177), .A2(G378), .A3(new_n1213), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT122), .ZN(new_n1257));
  OAI21_X1  g1057(.A(KEYINPUT121), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT121), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1210), .A2(new_n1259), .A3(new_n1211), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(new_n1260), .A3(new_n744), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1206), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(new_n984), .B2(new_n1170), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1257), .B1(new_n1263), .B2(G378), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1119), .A2(new_n1169), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1265), .A2(new_n984), .A3(new_n1212), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n743), .B1(new_n1212), .B2(KEYINPUT121), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1207), .B1(new_n1267), .B2(new_n1260), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1126), .A2(new_n1146), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(KEYINPUT114), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1126), .A2(new_n1121), .A3(new_n1146), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1269), .A2(new_n1273), .A3(KEYINPUT122), .A4(new_n1120), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1264), .A2(new_n1274), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1242), .B(new_n1255), .C1(new_n1256), .C2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(KEYINPUT62), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1242), .B1(new_n1256), .B2(new_n1275), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n671), .A2(G213), .A3(G2897), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1279), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1280), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1278), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT61), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1177), .A2(G378), .A3(new_n1213), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1287), .A2(new_n1264), .A3(new_n1274), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT62), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1288), .A2(new_n1289), .A3(new_n1242), .A4(new_n1255), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1277), .A2(new_n1285), .A3(new_n1286), .A4(new_n1290), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(G393), .B(new_n820), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT125), .ZN(new_n1293));
  INV_X1    g1093(.A(G390), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1008), .A2(new_n1293), .A3(new_n1294), .ZN(new_n1295));
  OAI211_X1 g1095(.A(G390), .B(new_n960), .C1(new_n985), .C2(new_n1007), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1293), .B1(new_n1008), .B2(new_n1294), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1292), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1296), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1300), .A2(new_n1292), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT126), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(G390), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1294), .A2(KEYINPUT126), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1010), .A2(new_n1011), .A3(new_n1303), .A4(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1301), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1299), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1291), .A2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT127), .B1(new_n1307), .B2(new_n1286), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT127), .ZN(new_n1311));
  AOI211_X1 g1111(.A(new_n1311), .B(KEYINPUT61), .C1(new_n1299), .C2(new_n1306), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1280), .A2(new_n1283), .A3(KEYINPUT124), .ZN(new_n1314));
  AOI21_X1  g1114(.A(KEYINPUT124), .B1(new_n1280), .B2(new_n1283), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1278), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1288), .A2(KEYINPUT63), .A3(new_n1242), .A4(new_n1255), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT63), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1276), .A2(new_n1319), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1313), .A2(new_n1317), .A3(new_n1318), .A4(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1309), .A2(new_n1321), .ZN(G405));
  XNOR2_X1  g1122(.A(G375), .B(G378), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(new_n1281), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1324), .B1(new_n1254), .B2(new_n1323), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(new_n1308), .ZN(new_n1326));
  OAI211_X1 g1126(.A(new_n1324), .B(new_n1307), .C1(new_n1254), .C2(new_n1323), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(G402));
endmodule


