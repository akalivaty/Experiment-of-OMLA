//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 1 1 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 0 1 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  AOI21_X1  g004(.A(G128), .B1(new_n188), .B2(new_n190), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n189), .A2(KEYINPUT1), .A3(G146), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT66), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT66), .ZN(new_n195));
  XNOR2_X1  g009(.A(G143), .B(G146), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n192), .B(new_n195), .C1(new_n196), .C2(G128), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(new_n198), .A3(G128), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n194), .A2(new_n197), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT71), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n194), .A2(new_n197), .A3(KEYINPUT71), .A4(new_n199), .ZN(new_n203));
  INV_X1    g017(.A(G134), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G137), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n205), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  INV_X1    g024(.A(G137), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(G134), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(G134), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n209), .A2(new_n210), .A3(new_n213), .A4(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(G131), .B1(new_n212), .B2(new_n205), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT70), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n216), .A2(KEYINPUT70), .A3(new_n217), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n202), .A2(new_n203), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G119), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G116), .ZN(new_n224));
  INV_X1    g038(.A(G116), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G119), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT2), .A2(G113), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT2), .ZN(new_n230));
  INV_X1    g044(.A(G113), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n231), .A3(KEYINPUT67), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n233), .B1(KEYINPUT2), .B2(G113), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n229), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n227), .B1(new_n235), .B2(KEYINPUT68), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n237));
  AOI211_X1 g051(.A(new_n237), .B(new_n229), .C1(new_n232), .C2(new_n234), .ZN(new_n238));
  OAI21_X1  g052(.A(KEYINPUT69), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  NOR3_X1   g053(.A1(new_n233), .A2(KEYINPUT2), .A3(G113), .ZN(new_n240));
  AOI21_X1  g054(.A(KEYINPUT67), .B1(new_n230), .B2(new_n231), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n228), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n237), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n235), .A2(KEYINPUT68), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n243), .A2(new_n244), .A3(new_n245), .A4(new_n227), .ZN(new_n246));
  INV_X1    g060(.A(new_n227), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n235), .A2(new_n247), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n239), .A2(new_n246), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n188), .A2(new_n190), .ZN(new_n250));
  NOR2_X1   g064(.A1(KEYINPUT0), .A2(G128), .ZN(new_n251));
  AND2_X1   g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n253), .B1(new_n250), .B2(new_n252), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n212), .B1(new_n214), .B2(new_n206), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n255), .A2(new_n210), .A3(new_n209), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n210), .B1(new_n255), .B2(new_n209), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n254), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n222), .A2(new_n249), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT28), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G101), .ZN(new_n262));
  XOR2_X1   g076(.A(KEYINPUT73), .B(G237), .Z(new_n263));
  AND2_X1   g077(.A1(KEYINPUT74), .A2(G953), .ZN(new_n264));
  NOR2_X1   g078(.A1(KEYINPUT74), .A2(G953), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n263), .A2(G210), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT27), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT26), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT27), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n263), .A2(new_n270), .A3(G210), .A4(new_n266), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n268), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n269), .B1(new_n268), .B2(new_n271), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n262), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n274), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n276), .A2(G101), .A3(new_n272), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n222), .A2(new_n249), .A3(KEYINPUT28), .A4(new_n258), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT65), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n258), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n200), .A2(new_n217), .A3(new_n216), .ZN(new_n282));
  OAI211_X1 g096(.A(KEYINPUT65), .B(new_n254), .C1(new_n256), .C2(new_n257), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n239), .A2(new_n246), .A3(new_n248), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n261), .A2(new_n278), .A3(new_n279), .A4(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT76), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT29), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n291), .B1(new_n287), .B2(new_n288), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT30), .ZN(new_n293));
  INV_X1    g107(.A(new_n257), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n216), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n293), .B1(new_n295), .B2(new_n254), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n222), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT72), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n284), .A2(new_n293), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n222), .A2(new_n296), .A3(KEYINPUT72), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n299), .A2(new_n285), .A3(new_n300), .A4(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n278), .B1(new_n302), .B2(new_n259), .ZN(new_n303));
  NOR3_X1   g117(.A1(new_n290), .A2(new_n292), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n259), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n249), .B1(new_n222), .B2(new_n258), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT28), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT77), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT77), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n309), .B(KEYINPUT28), .C1(new_n305), .C2(new_n306), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n275), .A2(new_n277), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n311), .A2(new_n291), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n308), .A2(new_n261), .A3(new_n310), .A4(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G902), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(G472), .B1(new_n304), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT32), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n317), .A2(G472), .A3(G902), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n261), .A2(new_n279), .A3(new_n286), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n311), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n305), .A2(new_n311), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT31), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n302), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n322), .B1(new_n302), .B2(new_n321), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n320), .B(new_n323), .C1(new_n324), .C2(KEYINPUT75), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n324), .A2(KEYINPUT75), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n318), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n316), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n302), .A2(new_n321), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT31), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AND2_X1   g146(.A1(new_n323), .A2(new_n320), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n324), .A2(KEYINPUT75), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(G472), .A2(G902), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT32), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT78), .B1(new_n328), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n302), .A2(new_n259), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n311), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n289), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n314), .B(new_n313), .C1(new_n341), .C2(new_n292), .ZN(new_n342));
  AOI22_X1  g156(.A1(new_n342), .A2(G472), .B1(new_n335), .B2(new_n318), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT78), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n336), .B1(new_n325), .B2(new_n326), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n317), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n343), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n338), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G234), .ZN(new_n349));
  OAI21_X1  g163(.A(G217), .B1(new_n349), .B2(G902), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n266), .A2(G221), .A3(G234), .ZN(new_n351));
  XOR2_X1   g165(.A(new_n351), .B(KEYINPUT22), .Z(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(new_n211), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT16), .ZN(new_n354));
  INV_X1    g168(.A(G140), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n355), .A3(G125), .ZN(new_n356));
  XOR2_X1   g170(.A(G125), .B(G140), .Z(new_n357));
  OAI21_X1  g171(.A(new_n356), .B1(new_n357), .B2(new_n354), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n187), .ZN(new_n359));
  OAI211_X1 g173(.A(G146), .B(new_n356), .C1(new_n357), .C2(new_n354), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n223), .A2(G128), .ZN(new_n362));
  NAND2_X1  g176(.A1(KEYINPUT23), .A2(G119), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n223), .A2(G128), .ZN(new_n364));
  OAI221_X1 g178(.A(new_n362), .B1(G128), .B2(new_n363), .C1(new_n364), .C2(KEYINPUT23), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G110), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT24), .B(G110), .ZN(new_n367));
  OR2_X1    g181(.A1(new_n364), .A2(KEYINPUT79), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n364), .A2(KEYINPUT79), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n362), .A3(new_n369), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n361), .B(new_n366), .C1(new_n367), .C2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n367), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n372), .B1(G110), .B2(new_n365), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n373), .B(new_n360), .C1(G146), .C2(new_n357), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n353), .A2(new_n371), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n371), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n352), .B(G137), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n375), .A2(new_n378), .A3(new_n314), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n350), .B1(new_n379), .B2(KEYINPUT25), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n380), .B1(KEYINPUT25), .B2(new_n379), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n375), .A2(new_n378), .ZN(new_n382));
  AOI21_X1  g196(.A(G902), .B1(new_n349), .B2(G217), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(KEYINPUT9), .B(G234), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n386), .B(KEYINPUT80), .ZN(new_n387));
  OAI21_X1  g201(.A(G221), .B1(new_n387), .B2(G902), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G104), .ZN(new_n390));
  NOR3_X1   g204(.A1(new_n390), .A2(KEYINPUT3), .A3(G107), .ZN(new_n391));
  INV_X1    g205(.A(G107), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT81), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n393), .A2(G104), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n390), .A2(KEYINPUT81), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n392), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n391), .B1(new_n396), .B2(KEYINPUT3), .ZN(new_n397));
  XNOR2_X1  g211(.A(KEYINPUT81), .B(G104), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT82), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n398), .A2(new_n399), .A3(G107), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n399), .B1(new_n398), .B2(G107), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n397), .B(new_n262), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n396), .A2(KEYINPUT3), .ZN(new_n403));
  INV_X1    g217(.A(new_n391), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n403), .B(new_n404), .C1(new_n400), .C2(new_n401), .ZN(new_n405));
  AND2_X1   g219(.A1(KEYINPUT83), .A2(G101), .ZN(new_n406));
  AOI22_X1  g220(.A1(new_n402), .A2(KEYINPUT4), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n405), .A2(KEYINPUT4), .A3(new_n406), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n254), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n202), .A2(new_n203), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n396), .B1(G104), .B2(new_n392), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G101), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n402), .A2(KEYINPUT10), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n295), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n199), .B(new_n192), .C1(G128), .C2(new_n196), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n402), .A2(new_n412), .A3(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT10), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n409), .A2(new_n414), .A3(new_n415), .A4(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n266), .A2(G227), .ZN(new_n421));
  XOR2_X1   g235(.A(G110), .B(G140), .Z(new_n422));
  XNOR2_X1  g236(.A(new_n421), .B(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  AOI22_X1  g240(.A1(new_n410), .A2(new_n413), .B1(new_n418), .B2(new_n417), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n409), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n295), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n415), .A2(KEYINPUT84), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n402), .A2(new_n412), .A3(new_n416), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n200), .B1(new_n402), .B2(new_n412), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT12), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT12), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n430), .B(new_n435), .C1(new_n431), .C2(new_n432), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n420), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  AOI22_X1  g251(.A1(new_n426), .A2(new_n429), .B1(new_n437), .B2(new_n423), .ZN(new_n438));
  OAI21_X1  g252(.A(G469), .B1(new_n438), .B2(G902), .ZN(new_n439));
  INV_X1    g253(.A(G469), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n424), .B1(new_n429), .B2(new_n420), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n434), .A2(new_n436), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n425), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n440), .B(new_n314), .C1(new_n441), .C2(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n389), .B1(new_n439), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n285), .B1(new_n407), .B2(new_n408), .ZN(new_n446));
  XNOR2_X1  g260(.A(G110), .B(G122), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT85), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n247), .A2(KEYINPUT5), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n224), .A2(KEYINPUT5), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n450), .A2(new_n231), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n449), .A2(new_n451), .B1(new_n235), .B2(new_n247), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n402), .A2(new_n448), .A3(new_n412), .A4(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n402), .A2(new_n412), .A3(new_n452), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT85), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n446), .A2(new_n447), .A3(new_n453), .A4(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT87), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n402), .A2(new_n412), .ZN(new_n459));
  INV_X1    g273(.A(new_n452), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n402), .A2(KEYINPUT87), .A3(new_n412), .A4(new_n452), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n458), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n447), .B(KEYINPUT8), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G125), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n200), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n254), .A2(G125), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT7), .ZN(new_n471));
  XOR2_X1   g285(.A(KEYINPUT86), .B(G224), .Z(new_n472));
  NOR2_X1   g286(.A1(new_n472), .A2(G953), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n470), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n470), .A2(new_n474), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n469), .A2(new_n473), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n474), .A2(new_n471), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n456), .A2(new_n465), .A3(new_n475), .A4(new_n479), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n480), .A2(new_n314), .ZN(new_n481));
  OAI21_X1  g295(.A(G210), .B1(G237), .B2(G902), .ZN(new_n482));
  XOR2_X1   g296(.A(new_n482), .B(KEYINPUT88), .Z(new_n483));
  INV_X1    g297(.A(new_n447), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n402), .A2(KEYINPUT4), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n405), .A2(new_n406), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n405), .A2(KEYINPUT4), .A3(new_n406), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n249), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n455), .A2(new_n453), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n484), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(KEYINPUT6), .A3(new_n456), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT6), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n493), .B(new_n484), .C1(new_n489), .C2(new_n490), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n476), .A2(new_n477), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n492), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n481), .A2(new_n483), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n483), .B1(new_n481), .B2(new_n496), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(G214), .B1(G237), .B2(G902), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n263), .A2(G214), .A3(new_n266), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n189), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n263), .A2(G143), .A3(G214), .A4(new_n266), .ZN(new_n503));
  NAND2_X1  g317(.A1(KEYINPUT18), .A2(G131), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n357), .B(G146), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n504), .B1(new_n502), .B2(new_n503), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT90), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n508), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT90), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n510), .A2(new_n511), .A3(new_n506), .A4(new_n505), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n210), .B1(new_n502), .B2(new_n503), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n361), .B1(new_n514), .B2(KEYINPUT17), .ZN(new_n515));
  INV_X1    g329(.A(new_n514), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n502), .A2(new_n210), .A3(new_n503), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n515), .B1(new_n518), .B2(KEYINPUT17), .ZN(new_n519));
  XNOR2_X1  g333(.A(G113), .B(G122), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n520), .B(new_n390), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n513), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n521), .B1(new_n513), .B2(new_n519), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n314), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(G475), .ZN(new_n526));
  INV_X1    g340(.A(G217), .ZN(new_n527));
  NOR3_X1   g341(.A1(new_n387), .A2(new_n527), .A3(G953), .ZN(new_n528));
  XNOR2_X1  g342(.A(G128), .B(G143), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT13), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n189), .A2(G128), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n530), .B(G134), .C1(KEYINPUT13), .C2(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(G116), .B(G122), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(new_n392), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n529), .A2(new_n204), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n532), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n529), .B(new_n204), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n225), .A2(KEYINPUT14), .A3(G122), .ZN(new_n538));
  INV_X1    g352(.A(new_n533), .ZN(new_n539));
  OAI211_X1 g353(.A(G107), .B(new_n538), .C1(new_n539), .C2(KEYINPUT14), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n533), .A2(new_n392), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n537), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n528), .A2(new_n536), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n528), .B1(new_n536), .B2(new_n542), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n314), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(G478), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n546), .B1(KEYINPUT15), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT15), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n545), .A2(new_n549), .A3(G478), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G952), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(G953), .ZN(new_n553));
  NAND2_X1  g367(.A1(G234), .A2(G237), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(KEYINPUT21), .B(G898), .ZN(new_n556));
  XOR2_X1   g370(.A(new_n556), .B(KEYINPUT94), .Z(new_n557));
  INV_X1    g371(.A(new_n266), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n558), .A2(G902), .A3(new_n554), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n555), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n551), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT89), .B(KEYINPUT20), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n516), .A2(KEYINPUT91), .A3(new_n517), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT91), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n502), .A2(new_n210), .A3(new_n503), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n565), .B1(new_n566), .B2(new_n514), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n357), .B(KEYINPUT19), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n360), .B1(new_n569), .B2(G146), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(KEYINPUT92), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n568), .A2(new_n571), .B1(new_n512), .B2(new_n509), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n522), .B1(new_n572), .B2(new_n521), .ZN(new_n573));
  NOR2_X1   g387(.A1(G475), .A2(G902), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n563), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n574), .ZN(new_n576));
  OR2_X1    g390(.A1(new_n576), .A2(KEYINPUT93), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT20), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(KEYINPUT93), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n568), .A2(new_n571), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n513), .ZN(new_n583));
  INV_X1    g397(.A(new_n521), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n581), .B1(new_n585), .B2(new_n522), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n526), .B(new_n562), .C1(new_n575), .C2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n445), .A2(new_n499), .A3(new_n500), .A4(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n348), .A2(new_n385), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(G101), .ZN(G3));
  NAND2_X1  g406(.A1(G469), .A2(G902), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n437), .A2(new_n423), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n415), .B1(new_n427), .B2(new_n409), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n594), .B(G469), .C1(new_n595), .C2(new_n425), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n444), .A2(new_n593), .A3(new_n596), .ZN(new_n597));
  AND4_X1   g411(.A1(new_n345), .A2(new_n597), .A3(new_n385), .A4(new_n388), .ZN(new_n598));
  AOI21_X1  g412(.A(KEYINPUT75), .B1(new_n329), .B2(KEYINPUT31), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n323), .A2(new_n320), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(G902), .B1(new_n601), .B2(new_n334), .ZN(new_n602));
  INV_X1    g416(.A(G472), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT95), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n335), .A2(new_n314), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT95), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n605), .A2(new_n606), .A3(G472), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n598), .A2(new_n604), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT33), .ZN(new_n609));
  OR3_X1    g423(.A1(new_n543), .A2(new_n544), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n609), .B1(new_n543), .B2(new_n544), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n547), .A2(G902), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(KEYINPUT96), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT96), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n610), .A2(new_n615), .A3(new_n611), .A4(new_n612), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n545), .A2(KEYINPUT97), .A3(new_n547), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT97), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n618), .B1(new_n546), .B2(G478), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n614), .A2(new_n616), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n575), .A2(new_n586), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n525), .A2(G475), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n481), .A2(new_n496), .ZN(new_n625));
  INV_X1    g439(.A(new_n483), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n481), .A2(new_n483), .A3(new_n496), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n627), .A2(new_n500), .A3(new_n628), .A4(new_n560), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n608), .A2(new_n624), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT34), .B(G104), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT98), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n630), .B(new_n632), .ZN(G6));
  NAND3_X1  g447(.A1(new_n573), .A2(new_n574), .A3(new_n563), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n573), .A2(new_n574), .ZN(new_n635));
  INV_X1    g449(.A(new_n563), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n623), .B1(new_n634), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n551), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n608), .A2(new_n629), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT35), .B(G107), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G9));
  NAND3_X1  g456(.A1(new_n604), .A2(new_n607), .A3(new_n345), .ZN(new_n643));
  INV_X1    g457(.A(new_n500), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n497), .A2(new_n498), .A3(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n377), .A2(KEYINPUT36), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(new_n376), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n383), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n381), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n645), .A2(new_n445), .A3(new_n588), .A4(new_n649), .ZN(new_n650));
  OR2_X1    g464(.A1(new_n643), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT37), .B(G110), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G12));
  XNOR2_X1  g467(.A(new_n555), .B(KEYINPUT99), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n654), .B1(G900), .B2(new_n559), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n638), .A2(new_n551), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n597), .A2(new_n388), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n627), .A2(new_n500), .A3(new_n628), .ZN(new_n658));
  INV_X1    g472(.A(new_n649), .ZN(new_n659));
  NOR4_X1   g473(.A1(new_n656), .A2(new_n657), .A3(new_n658), .A4(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n348), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G128), .ZN(G30));
  AND2_X1   g476(.A1(new_n499), .A2(KEYINPUT38), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n499), .A2(KEYINPUT38), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n622), .A2(new_n623), .ZN(new_n666));
  INV_X1    g480(.A(new_n551), .ZN(new_n667));
  OR4_X1    g481(.A1(new_n644), .A2(new_n666), .A3(new_n667), .A4(new_n649), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n339), .A2(new_n278), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n305), .A2(new_n306), .ZN(new_n670));
  AOI21_X1  g484(.A(G902), .B1(new_n670), .B2(new_n311), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n603), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n672), .B1(new_n335), .B2(new_n318), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n346), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n665), .A2(new_n668), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n655), .B(KEYINPUT39), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n445), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(new_n678), .B(KEYINPUT40), .Z(new_n679));
  NAND2_X1  g493(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT100), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(new_n189), .ZN(G45));
  NOR3_X1   g496(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n621), .B(new_n655), .C1(new_n622), .C2(new_n623), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n348), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G146), .ZN(G48));
  INV_X1    g501(.A(new_n420), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n423), .B1(new_n688), .B2(new_n595), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n689), .B1(new_n425), .B2(new_n442), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n314), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(G469), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n692), .A2(new_n388), .A3(new_n444), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n693), .A2(new_n629), .A3(new_n624), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n348), .A2(new_n385), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(KEYINPUT101), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n381), .A2(new_n384), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n697), .B1(new_n338), .B2(new_n347), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT101), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n698), .A2(new_n699), .A3(new_n694), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT41), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G113), .ZN(G15));
  NOR3_X1   g517(.A1(new_n693), .A2(new_n639), .A3(new_n629), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n328), .A2(KEYINPUT78), .A3(new_n337), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n344), .B1(new_n343), .B2(new_n346), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n704), .B(new_n385), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G116), .ZN(G18));
  NOR4_X1   g522(.A1(new_n693), .A2(new_n658), .A3(new_n587), .A4(new_n659), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n709), .B1(new_n705), .B2(new_n706), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G119), .ZN(G21));
  NOR2_X1   g525(.A1(new_n602), .A2(new_n603), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n308), .A2(new_n261), .A3(new_n310), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n330), .B(new_n323), .C1(new_n713), .C2(new_n278), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n714), .A2(new_n336), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n693), .A2(new_n561), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n658), .A2(new_n666), .A3(new_n667), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n697), .B(KEYINPUT102), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n716), .A2(new_n717), .A3(new_n718), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G122), .ZN(G24));
  NOR3_X1   g535(.A1(new_n712), .A2(new_n715), .A3(new_n659), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n693), .A2(new_n658), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(new_n685), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G125), .ZN(G27));
  NAND2_X1  g539(.A1(new_n573), .A2(new_n580), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n637), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n620), .B1(new_n727), .B2(new_n526), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n445), .A2(new_n728), .A3(new_n655), .ZN(new_n729));
  NOR4_X1   g543(.A1(new_n729), .A2(KEYINPUT42), .A3(new_n644), .A4(new_n499), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n657), .A2(new_n684), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n346), .A2(new_n327), .A3(new_n316), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n499), .A2(new_n644), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n731), .A2(new_n732), .A3(new_n719), .A4(new_n733), .ZN(new_n734));
  AOI22_X1  g548(.A1(new_n698), .A2(new_n730), .B1(KEYINPUT42), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G131), .ZN(G33));
  NOR2_X1   g550(.A1(new_n656), .A2(new_n657), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n698), .A2(new_n733), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G134), .ZN(G36));
  NAND2_X1  g553(.A1(new_n666), .A2(new_n621), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n741), .B1(KEYINPUT105), .B2(KEYINPUT43), .ZN(new_n742));
  XNOR2_X1  g556(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n659), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT44), .B1(new_n745), .B2(new_n643), .ZN(new_n746));
  AOI211_X1 g560(.A(new_n644), .B(new_n746), .C1(new_n628), .C2(new_n627), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n438), .A2(KEYINPUT45), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n748), .A2(KEYINPUT103), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n748), .A2(KEYINPUT103), .ZN(new_n750));
  OAI21_X1  g564(.A(G469), .B1(new_n438), .B2(KEYINPUT45), .ZN(new_n751));
  OR3_X1    g565(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(KEYINPUT46), .A3(new_n593), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT104), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n753), .A2(new_n754), .A3(new_n444), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n754), .B1(new_n753), .B2(new_n444), .ZN(new_n756));
  AOI21_X1  g570(.A(KEYINPUT46), .B1(new_n752), .B2(new_n593), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n755), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n389), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n745), .A2(KEYINPUT44), .A3(new_n643), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n747), .A2(new_n677), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(KEYINPUT106), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(new_n211), .ZN(G39));
  INV_X1    g577(.A(KEYINPUT47), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(KEYINPUT47), .B1(new_n758), .B2(new_n389), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n733), .A2(new_n697), .A3(new_n685), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n348), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n765), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G140), .ZN(G42));
  NAND4_X1  g584(.A1(new_n741), .A2(new_n719), .A3(new_n500), .A4(new_n388), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n692), .A2(new_n444), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(KEYINPUT49), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n772), .A2(KEYINPUT49), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n771), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(new_n675), .A3(new_n665), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n654), .B1(new_n742), .B2(new_n744), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n732), .A2(new_n719), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n693), .A2(new_n644), .A3(new_n499), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n777), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT48), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n777), .A2(new_n716), .A3(new_n719), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n723), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n697), .A2(new_n555), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n780), .A2(new_n675), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n728), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n782), .A2(new_n553), .A3(new_n784), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n765), .A2(new_n766), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n789), .B1(new_n388), .B2(new_n772), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n790), .A2(new_n733), .A3(new_n783), .ZN(new_n791));
  NOR4_X1   g605(.A1(new_n663), .A2(new_n664), .A3(new_n500), .A4(new_n693), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n783), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT50), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n783), .A2(KEYINPUT50), .A3(new_n792), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n777), .A2(new_n722), .A3(new_n780), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n786), .A2(new_n666), .A3(new_n620), .ZN(new_n799));
  AND4_X1   g613(.A1(KEYINPUT51), .A2(new_n797), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n788), .B1(new_n791), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n798), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n802), .B1(new_n797), .B2(KEYINPUT111), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT111), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n795), .A2(new_n804), .A3(new_n796), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT112), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n803), .A2(KEYINPUT112), .A3(new_n805), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n791), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n801), .B1(new_n810), .B2(KEYINPUT51), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n707), .A2(new_n710), .A3(new_n720), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n813), .B1(new_n700), .B2(new_n696), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n499), .A2(new_n644), .A3(new_n659), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n445), .A2(new_n638), .A3(new_n667), .A4(new_n655), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n816), .B1(new_n338), .B2(new_n347), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n729), .A2(new_n712), .A3(new_n715), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n815), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n735), .A2(new_n819), .A3(new_n738), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT107), .ZN(new_n821));
  AOI211_X1 g635(.A(new_n697), .B(new_n589), .C1(new_n338), .C2(new_n347), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n727), .A2(new_n526), .A3(new_n551), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(new_n624), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n645), .A3(new_n560), .ZN(new_n825));
  OAI22_X1  g639(.A1(new_n608), .A2(new_n825), .B1(new_n643), .B2(new_n650), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n821), .B1(new_n822), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n629), .B1(new_n624), .B2(new_n823), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n828), .A2(new_n604), .A3(new_n607), .A4(new_n598), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n591), .A2(KEYINPUT107), .A3(new_n651), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n814), .A2(new_n820), .A3(new_n831), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n381), .A2(new_n648), .A3(new_n655), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(KEYINPUT109), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n834), .A2(new_n718), .A3(new_n445), .A4(new_n674), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n686), .A2(new_n661), .A3(new_n724), .A4(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT52), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n832), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT108), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n832), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n814), .A2(new_n820), .A3(new_n831), .A4(KEYINPUT108), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n836), .B(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n838), .B1(new_n841), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n839), .B1(new_n846), .B2(KEYINPUT110), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT110), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n848), .B(new_n838), .C1(new_n841), .C2(new_n845), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n812), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n832), .A2(new_n837), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT53), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n838), .B1(new_n832), .B2(new_n837), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n852), .A2(new_n812), .A3(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n811), .A2(new_n850), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(G952), .A2(G953), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n776), .B1(new_n855), .B2(new_n856), .ZN(G75));
  AOI21_X1  g671(.A(new_n314), .B1(new_n852), .B2(new_n853), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n483), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT113), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n860), .A2(KEYINPUT56), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT55), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n492), .A2(new_n494), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(new_n495), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT55), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n859), .A2(new_n866), .A3(new_n861), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n863), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n865), .B1(new_n863), .B2(new_n867), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n266), .A2(G952), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(G51));
  XOR2_X1   g685(.A(new_n593), .B(KEYINPUT57), .Z(new_n872));
  AOI21_X1  g686(.A(new_n812), .B1(new_n852), .B2(new_n853), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n872), .B1(new_n854), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n690), .ZN(new_n875));
  INV_X1    g689(.A(new_n752), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n858), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n870), .B1(new_n875), .B2(new_n877), .ZN(G54));
  NAND2_X1  g692(.A1(KEYINPUT58), .A2(G475), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT114), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n573), .B1(new_n858), .B2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT115), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n870), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n858), .A2(new_n573), .A3(new_n880), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n882), .B2(new_n881), .ZN(G60));
  INV_X1    g701(.A(KEYINPUT117), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n610), .A2(new_n611), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n846), .A2(KEYINPUT110), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n890), .A2(new_n849), .A3(new_n852), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n854), .B1(new_n891), .B2(KEYINPUT54), .ZN(new_n892));
  NAND2_X1  g706(.A1(G478), .A2(G902), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT59), .Z(new_n894));
  OAI211_X1 g708(.A(new_n888), .B(new_n889), .C1(new_n892), .C2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n894), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n897), .B1(new_n850), .B2(new_n854), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n888), .B1(new_n898), .B2(new_n889), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n889), .A2(new_n894), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n900), .B1(new_n854), .B2(new_n873), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT116), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n901), .A2(new_n902), .A3(new_n884), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n902), .B1(new_n901), .B2(new_n884), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n896), .A2(new_n899), .A3(new_n905), .ZN(G63));
  OAI21_X1  g720(.A(new_n884), .B1(KEYINPUT119), .B2(KEYINPUT61), .ZN(new_n907));
  NAND2_X1  g721(.A1(G217), .A2(G902), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT118), .Z(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT60), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n910), .B1(new_n852), .B2(new_n853), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n907), .B1(new_n911), .B2(new_n647), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n912), .B1(new_n382), .B2(new_n911), .ZN(new_n913));
  NAND2_X1  g727(.A1(KEYINPUT119), .A2(KEYINPUT61), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n913), .B(new_n914), .ZN(G66));
  INV_X1    g729(.A(new_n557), .ZN(new_n916));
  OAI21_X1  g730(.A(G953), .B1(new_n916), .B2(new_n472), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT121), .Z(new_n918));
  NAND2_X1  g732(.A1(new_n814), .A2(new_n831), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT120), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n918), .B1(new_n920), .B2(new_n558), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n864), .B1(G898), .B2(new_n266), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n921), .B(new_n922), .ZN(G69));
  AOI21_X1  g737(.A(new_n266), .B1(G227), .B2(G900), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT122), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT124), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n299), .A2(new_n301), .A3(new_n300), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(new_n569), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n686), .A2(new_n661), .A3(new_n724), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n680), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT62), .Z(new_n932));
  INV_X1    g746(.A(new_n678), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n698), .A2(new_n933), .A3(new_n733), .A4(new_n824), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n769), .A2(new_n761), .ZN(new_n936));
  AOI211_X1 g750(.A(new_n558), .B(new_n929), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n266), .A2(G900), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT123), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n929), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n759), .A2(new_n677), .A3(new_n718), .A4(new_n779), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n930), .A2(new_n735), .A3(new_n738), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n769), .A2(new_n761), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n940), .B1(new_n943), .B2(new_n266), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n926), .B(new_n927), .C1(new_n937), .C2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n935), .A2(new_n936), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n929), .A2(new_n558), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n943), .A2(new_n266), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n949), .B1(new_n950), .B2(new_n940), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n927), .B1(new_n951), .B2(new_n926), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n925), .B1(new_n946), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n937), .A2(new_n944), .ZN(new_n954));
  OAI21_X1  g768(.A(KEYINPUT124), .B1(new_n954), .B2(KEYINPUT122), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n955), .A2(new_n945), .A3(new_n924), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n953), .A2(new_n956), .ZN(G72));
  NAND4_X1  g771(.A1(new_n936), .A2(new_n920), .A3(new_n941), .A4(new_n942), .ZN(new_n958));
  NAND2_X1  g772(.A1(G472), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT63), .Z(new_n960));
  NAND2_X1  g774(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n339), .A2(new_n278), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n870), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n669), .ZN(new_n964));
  INV_X1    g778(.A(new_n960), .ZN(new_n965));
  INV_X1    g779(.A(new_n947), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n965), .B1(new_n966), .B2(new_n920), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT125), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI211_X1 g783(.A(KEYINPUT125), .B(new_n965), .C1(new_n966), .C2(new_n920), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n963), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n340), .A2(KEYINPUT126), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT126), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n329), .B1(new_n303), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n960), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT127), .Z(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(new_n847), .B2(new_n849), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n971), .A2(new_n977), .ZN(G57));
endmodule


