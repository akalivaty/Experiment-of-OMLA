//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 0 0 0 1 1 0 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 1 1 0 0 0 0 1 1 0 0 1 0 0 0 0 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n553, new_n555, new_n556, new_n557, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n600, new_n601, new_n602,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1180, new_n1181;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(G101), .A2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n470), .B1(new_n466), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  AND2_X1   g051(.A1(new_n466), .A2(KEYINPUT66), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n466), .A2(KEYINPUT66), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(new_n473), .ZN(new_n480));
  MUX2_X1   g055(.A(G100), .B(G112), .S(G2105), .Z(new_n481));
  AOI22_X1  g056(.A1(new_n480), .A2(G124), .B1(G2104), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n479), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n482), .A2(new_n484), .ZN(G162));
  NAND2_X1  g060(.A1(KEYINPUT4), .A2(G138), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT3), .ZN(new_n487));
  INV_X1    g062(.A(G2104), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n486), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AND2_X1   g066(.A1(G102), .A2(G2104), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n473), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G126), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n494), .B1(new_n489), .B2(new_n490), .ZN(new_n495));
  AND2_X1   g070(.A1(G114), .A2(G2104), .ZN(new_n496));
  OAI21_X1  g071(.A(G2105), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(G138), .B(new_n473), .C1(new_n464), .C2(new_n465), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n493), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT67), .A3(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n504), .A2(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  OAI21_X1  g087(.A(KEYINPUT68), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n505), .A2(new_n507), .B1(KEYINPUT5), .B2(new_n504), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT68), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n514), .A2(new_n515), .A3(new_n511), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT69), .B(G88), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(G75), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G62), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n520), .B1(new_n510), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n512), .A2(new_n504), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n522), .A2(G651), .B1(G50), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n519), .A2(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  NAND2_X1  g101(.A1(new_n523), .A2(G51), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  AND3_X1   g105(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n513), .A2(G89), .A3(new_n516), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n510), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n537), .A2(G651), .B1(G52), .B2(new_n523), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n513), .A2(G90), .A3(new_n516), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  NAND3_X1  g116(.A1(new_n513), .A2(G81), .A3(new_n516), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n523), .A2(G43), .ZN(new_n543));
  INV_X1    g118(.A(G68), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n504), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n545), .B1(new_n514), .B2(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(G651), .B1(new_n546), .B2(KEYINPUT70), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT70), .ZN(new_n548));
  AOI211_X1 g123(.A(new_n548), .B(new_n545), .C1(new_n514), .C2(G56), .ZN(new_n549));
  OAI211_X1 g124(.A(new_n542), .B(new_n543), .C1(new_n547), .C2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(G176));
  XOR2_X1   g129(.A(KEYINPUT71), .B(KEYINPUT8), .Z(new_n555));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n553), .A2(new_n557), .ZN(G188));
  NAND2_X1  g133(.A1(new_n517), .A2(G91), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n510), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G651), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n511), .A2(G53), .A3(G543), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT9), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n559), .A2(new_n563), .A3(new_n565), .ZN(G299));
  NAND2_X1  g141(.A1(new_n517), .A2(G87), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n523), .A2(G49), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(G288));
  NAND2_X1  g145(.A1(new_n517), .A2(G86), .ZN(new_n571));
  NAND2_X1  g146(.A1(G73), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(G61), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n510), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n574), .A2(G651), .B1(G48), .B2(new_n523), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n571), .A2(new_n575), .ZN(G305));
  NAND2_X1  g151(.A1(new_n517), .A2(G85), .ZN(new_n577));
  XOR2_X1   g152(.A(KEYINPUT72), .B(G47), .Z(new_n578));
  NAND2_X1  g153(.A1(new_n523), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(G651), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n577), .B(new_n579), .C1(new_n580), .C2(new_n581), .ZN(G290));
  NAND2_X1  g157(.A1(G301), .A2(G868), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n513), .A2(G92), .A3(new_n516), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT10), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n584), .B(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n514), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT73), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n580), .B1(new_n587), .B2(new_n588), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n589), .A2(new_n590), .B1(G54), .B2(new_n523), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n586), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(KEYINPUT74), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT74), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n586), .A2(new_n594), .A3(new_n591), .ZN(new_n595));
  AND2_X1   g170(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n583), .B1(new_n596), .B2(G868), .ZN(G284));
  OAI21_X1  g172(.A(new_n583), .B1(new_n596), .B2(G868), .ZN(G321));
  NAND2_X1  g173(.A1(new_n563), .A2(new_n565), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n599), .B1(G91), .B2(new_n517), .ZN(new_n600));
  OAI21_X1  g175(.A(KEYINPUT75), .B1(new_n600), .B2(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(G286), .A2(G868), .ZN(new_n602));
  MUX2_X1   g177(.A(KEYINPUT75), .B(new_n601), .S(new_n602), .Z(G297));
  MUX2_X1   g178(.A(KEYINPUT75), .B(new_n601), .S(new_n602), .Z(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n596), .B1(new_n605), .B2(G860), .ZN(G148));
  NAND3_X1  g181(.A1(new_n593), .A2(new_n605), .A3(new_n595), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT76), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n607), .A2(new_n608), .ZN(new_n611));
  OAI21_X1  g186(.A(G868), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n551), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  MUX2_X1   g189(.A(G99), .B(G111), .S(G2105), .Z(new_n615));
  AOI22_X1  g190(.A1(new_n480), .A2(G123), .B1(G2104), .B2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G135), .ZN(new_n617));
  INV_X1    g192(.A(new_n483), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(G2096), .Z(new_n620));
  NAND3_X1  g195(.A1(new_n473), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2100), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n620), .A2(new_n624), .ZN(G156));
  INV_X1    g200(.A(KEYINPUT14), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT15), .B(G2435), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2438), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2427), .ZN(new_n629));
  INV_X1    g204(.A(G2430), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n626), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n630), .B2(new_n629), .ZN(new_n632));
  XOR2_X1   g207(.A(G2451), .B(G2454), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT16), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT77), .ZN(new_n635));
  XOR2_X1   g210(.A(G2443), .B(G2446), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n632), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G1341), .B(G1348), .Z(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT78), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n641), .B(G14), .C1(new_n638), .C2(new_n639), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(G401));
  XNOR2_X1  g218(.A(G2072), .B(G2078), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(KEYINPUT17), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2084), .B(G2090), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n649), .B1(new_n646), .B2(new_n645), .ZN(new_n650));
  INV_X1    g225(.A(new_n646), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n651), .A2(new_n648), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n644), .B1(new_n652), .B2(KEYINPUT17), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n651), .A2(new_n644), .A3(new_n648), .ZN(new_n654));
  INV_X1    g229(.A(KEYINPUT18), .ZN(new_n655));
  AND2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  OAI22_X1  g232(.A1(new_n650), .A2(new_n653), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT79), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2096), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT80), .B(G2100), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(G227));
  XOR2_X1   g237(.A(G1961), .B(G1966), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT81), .ZN(new_n664));
  XOR2_X1   g239(.A(G1956), .B(G2474), .Z(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT82), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT20), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n664), .A2(new_n665), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n673), .A2(new_n669), .A3(new_n666), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n672), .B(new_n674), .C1(new_n669), .C2(new_n673), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1991), .B(G1996), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1981), .B(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n677), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(G229));
  MUX2_X1   g257(.A(G6), .B(G305), .S(G16), .Z(new_n683));
  XOR2_X1   g258(.A(KEYINPUT32), .B(G1981), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(G16), .A2(G22), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(G166), .B2(G16), .ZN(new_n687));
  INV_X1    g262(.A(G1971), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(G16), .A2(G23), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT85), .ZN(new_n691));
  INV_X1    g266(.A(G16), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n691), .B1(G288), .B2(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT33), .B(G1976), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n685), .A2(new_n689), .A3(new_n695), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n696), .A2(KEYINPUT34), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(KEYINPUT34), .ZN(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n699), .A2(KEYINPUT83), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(KEYINPUT83), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n703), .A2(G25), .ZN(new_n704));
  MUX2_X1   g279(.A(G95), .B(G107), .S(G2105), .Z(new_n705));
  AOI22_X1  g280(.A1(new_n480), .A2(G119), .B1(G2104), .B2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G131), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(new_n707), .B2(new_n618), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT84), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n704), .B1(new_n709), .B2(new_n703), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT35), .B(G1991), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  MUX2_X1   g287(.A(G24), .B(G290), .S(G16), .Z(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(G1986), .Z(new_n714));
  NAND4_X1  g289(.A1(new_n697), .A2(new_n698), .A3(new_n712), .A4(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT36), .Z(new_n716));
  NAND2_X1  g291(.A1(new_n483), .A2(G139), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT92), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT91), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT25), .Z(new_n721));
  NAND2_X1  g296(.A1(G115), .A2(G2104), .ZN(new_n722));
  INV_X1    g297(.A(G127), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n466), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n721), .B1(G2105), .B2(new_n724), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n718), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G29), .ZN(new_n727));
  NOR2_X1   g302(.A1(G29), .A2(G33), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT90), .Z(new_n729));
  NAND2_X1  g304(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G2072), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(G5), .A2(G16), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT97), .Z(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G301), .B2(new_n692), .ZN(new_n735));
  INV_X1    g310(.A(G1961), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT31), .B(G11), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT30), .B(G28), .Z(new_n739));
  OAI21_X1  g314(.A(new_n738), .B1(new_n739), .B2(G29), .ZN(new_n740));
  INV_X1    g315(.A(G2084), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT93), .ZN(new_n742));
  INV_X1    g317(.A(G34), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(KEYINPUT24), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n702), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(KEYINPUT24), .B2(new_n743), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n742), .B1(new_n702), .B2(new_n744), .ZN(new_n747));
  OAI22_X1  g322(.A1(new_n746), .A2(new_n747), .B1(new_n475), .B2(new_n699), .ZN(new_n748));
  OAI22_X1  g323(.A1(new_n619), .A2(new_n702), .B1(new_n741), .B2(new_n748), .ZN(new_n749));
  AOI211_X1 g324(.A(new_n740), .B(new_n749), .C1(new_n741), .C2(new_n748), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n735), .A2(new_n736), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n703), .A2(G27), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G164), .B2(new_n703), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(G2078), .Z(new_n754));
  NAND3_X1  g329(.A1(new_n750), .A2(new_n751), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n692), .A2(G20), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT23), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n600), .B2(new_n692), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G1956), .ZN(new_n759));
  NOR4_X1   g334(.A1(new_n732), .A2(new_n737), .A3(new_n755), .A4(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n703), .A2(G35), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G162), .B2(new_n703), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT29), .Z(new_n763));
  INV_X1    g338(.A(G2090), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT98), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(KEYINPUT95), .B1(G29), .B2(G32), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n483), .A2(G141), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n480), .A2(G129), .ZN(new_n770));
  NAND3_X1  g345(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT26), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  AND2_X1   g349(.A1(G105), .A2(G2104), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n773), .A2(new_n774), .B1(new_n473), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n769), .A2(new_n770), .A3(new_n776), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT94), .Z(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n768), .B1(new_n779), .B2(new_n699), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n778), .A2(KEYINPUT95), .A3(G29), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT27), .B(G1996), .Z(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(G1966), .ZN(new_n785));
  NAND2_X1  g360(.A1(G168), .A2(G16), .ZN(new_n786));
  NOR2_X1   g361(.A1(G16), .A2(G21), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(KEYINPUT96), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n786), .B2(KEYINPUT96), .ZN(new_n789));
  OAI22_X1  g364(.A1(new_n763), .A2(new_n764), .B1(new_n785), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n785), .B2(new_n789), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n760), .A2(new_n767), .A3(new_n784), .A4(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n692), .A2(G4), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n596), .B2(new_n692), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G1348), .ZN(new_n796));
  NOR2_X1   g371(.A1(G16), .A2(G19), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n551), .B2(G16), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G1341), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n702), .A2(G26), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT28), .Z(new_n801));
  NAND2_X1  g376(.A1(new_n480), .A2(G128), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT86), .ZN(new_n803));
  MUX2_X1   g378(.A(G104), .B(G116), .S(G2105), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(G2104), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT87), .Z(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n483), .B2(G140), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n803), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n801), .B1(new_n808), .B2(G29), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT88), .B(G2067), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n796), .A2(new_n799), .A3(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT89), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n793), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n812), .A2(new_n813), .ZN(new_n816));
  OAI21_X1  g391(.A(KEYINPUT99), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n816), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT99), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n793), .A2(new_n818), .A3(new_n819), .A4(new_n814), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n716), .B1(new_n817), .B2(new_n820), .ZN(G311));
  NAND2_X1  g396(.A1(new_n817), .A2(new_n820), .ZN(new_n822));
  INV_X1    g397(.A(new_n716), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(G150));
  NAND2_X1  g399(.A1(new_n596), .A2(G559), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT38), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n550), .A2(KEYINPUT101), .ZN(new_n827));
  INV_X1    g402(.A(G56), .ZN(new_n828));
  OAI22_X1  g403(.A1(new_n510), .A2(new_n828), .B1(new_n544), .B2(new_n504), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(new_n548), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n546), .A2(KEYINPUT70), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n830), .A2(G651), .A3(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT101), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n832), .A2(new_n833), .A3(new_n543), .A4(new_n542), .ZN(new_n834));
  NAND2_X1  g409(.A1(G80), .A2(G543), .ZN(new_n835));
  INV_X1    g410(.A(G67), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n835), .B1(new_n510), .B2(new_n836), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n837), .A2(G651), .B1(G55), .B2(new_n523), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT100), .B(G93), .Z(new_n839));
  NAND3_X1  g414(.A1(new_n513), .A2(new_n516), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n827), .A2(new_n834), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n550), .A2(KEYINPUT101), .A3(new_n841), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n826), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n847));
  AOI21_X1  g422(.A(G860), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n847), .B2(new_n846), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n841), .A2(G860), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT37), .Z(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(G145));
  INV_X1    g427(.A(KEYINPUT40), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n808), .B(new_n501), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n709), .B(KEYINPUT102), .ZN(new_n855));
  MUX2_X1   g430(.A(G106), .B(G118), .S(G2105), .Z(new_n856));
  AOI22_X1  g431(.A1(new_n480), .A2(G130), .B1(G2104), .B2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(G142), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n857), .B1(new_n858), .B2(new_n618), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n622), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT84), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n708), .B(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT102), .ZN(new_n864));
  INV_X1    g439(.A(new_n860), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n854), .B1(new_n861), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n861), .A2(new_n866), .A3(new_n854), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n726), .A2(new_n777), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n870), .B1(new_n726), .B2(new_n779), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n868), .A2(new_n869), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n869), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n871), .B1(new_n874), .B2(new_n867), .ZN(new_n875));
  XNOR2_X1  g450(.A(G162), .B(new_n475), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n876), .B(new_n619), .Z(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n873), .A2(new_n875), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(G37), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n878), .B1(new_n873), .B2(new_n875), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n853), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n882), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n884), .A2(KEYINPUT40), .A3(new_n880), .A4(new_n879), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n883), .A2(new_n885), .ZN(G395));
  NOR2_X1   g461(.A1(new_n841), .A2(G868), .ZN(new_n887));
  XNOR2_X1  g462(.A(G290), .B(G288), .ZN(new_n888));
  XNOR2_X1  g463(.A(G303), .B(G305), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n888), .B(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT103), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n891), .B1(new_n610), .B2(new_n611), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n596), .A2(KEYINPUT76), .A3(new_n605), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n893), .A2(KEYINPUT103), .A3(new_n609), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n845), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n845), .B1(new_n892), .B2(new_n894), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n586), .A2(new_n600), .A3(new_n591), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n600), .B1(new_n586), .B2(new_n591), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n896), .A2(new_n897), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n900), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(KEYINPUT41), .A3(new_n898), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(new_n899), .B2(new_n900), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n845), .ZN(new_n909));
  INV_X1    g484(.A(new_n894), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT103), .B1(new_n893), .B2(new_n609), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n908), .B1(new_n912), .B2(new_n895), .ZN(new_n913));
  NOR3_X1   g488(.A1(new_n903), .A2(new_n913), .A3(KEYINPUT42), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT42), .ZN(new_n915));
  INV_X1    g490(.A(new_n908), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(new_n896), .B2(new_n897), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n912), .A2(new_n895), .A3(new_n901), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n890), .B1(new_n914), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT42), .B1(new_n903), .B2(new_n913), .ZN(new_n921));
  INV_X1    g496(.A(new_n890), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n917), .A2(new_n915), .A3(new_n918), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n887), .B1(new_n925), .B2(G868), .ZN(G295));
  AOI21_X1  g501(.A(new_n887), .B1(new_n925), .B2(G868), .ZN(G331));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n928));
  NAND2_X1  g503(.A1(G168), .A2(G171), .ZN(new_n929));
  NAND2_X1  g504(.A1(G286), .A2(G301), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n845), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n843), .A2(new_n844), .A3(new_n930), .A4(new_n929), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n932), .A2(KEYINPUT105), .A3(new_n933), .ZN(new_n934));
  OR3_X1    g509(.A1(new_n845), .A2(KEYINPUT105), .A3(new_n931), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n933), .A2(KEYINPUT104), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n929), .A2(new_n930), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT104), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n938), .A2(new_n939), .A3(new_n843), .A4(new_n844), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n937), .A2(new_n940), .A3(new_n932), .ZN(new_n941));
  OAI22_X1  g516(.A1(new_n936), .A2(new_n908), .B1(new_n941), .B2(new_n902), .ZN(new_n942));
  AOI21_X1  g517(.A(G37), .B1(new_n942), .B2(new_n922), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n936), .A2(new_n901), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n916), .A2(new_n941), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(new_n890), .A3(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n946), .A2(KEYINPUT106), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n948));
  AOI22_X1  g523(.A1(new_n936), .A2(new_n901), .B1(new_n916), .B2(new_n941), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n948), .B1(new_n949), .B2(new_n890), .ZN(new_n950));
  OAI211_X1 g525(.A(KEYINPUT108), .B(new_n943), .C1(new_n947), .C2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n946), .A2(KEYINPUT106), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n949), .A2(new_n948), .A3(new_n890), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT108), .B1(new_n955), .B2(new_n943), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT43), .B1(new_n952), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n880), .B1(new_n949), .B2(new_n890), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n958), .B1(new_n953), .B2(new_n954), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n928), .B1(new_n957), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT107), .B1(new_n959), .B2(new_n960), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n944), .A2(new_n945), .ZN(new_n964));
  AOI21_X1  g539(.A(G37), .B1(new_n964), .B2(new_n922), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n965), .B1(new_n947), .B2(new_n950), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT107), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n966), .A2(new_n967), .A3(KEYINPUT43), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n955), .A2(new_n960), .A3(new_n943), .ZN(new_n969));
  AND4_X1   g544(.A1(new_n928), .A2(new_n963), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n962), .A2(new_n970), .ZN(G397));
  INV_X1    g546(.A(KEYINPUT50), .ZN(new_n972));
  INV_X1    g547(.A(G1384), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n501), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT111), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT111), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n501), .A2(new_n976), .A3(new_n972), .A4(new_n973), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT119), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n469), .A2(new_n474), .A3(G40), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n501), .A2(new_n973), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n980), .B1(new_n981), .B2(KEYINPUT50), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n978), .A2(new_n979), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n979), .B1(new_n978), .B2(new_n982), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n983), .A2(new_n984), .A3(G1961), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n981), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n973), .ZN(new_n988));
  INV_X1    g563(.A(new_n980), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n991));
  NOR3_X1   g566(.A1(new_n990), .A2(new_n991), .A3(G2078), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT124), .B1(new_n985), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT124), .ZN(new_n994));
  INV_X1    g569(.A(new_n992), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n978), .A2(new_n982), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT119), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n978), .A2(new_n979), .A3(new_n982), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n994), .B(new_n995), .C1(new_n999), .C2(G1961), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n991), .B1(new_n990), .B2(G2078), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n993), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n1002), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT125), .B1(new_n1002), .B2(G171), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n995), .B(new_n1001), .C1(new_n999), .C2(G1961), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1005), .A2(G171), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n1003), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT126), .B1(new_n1007), .B2(KEYINPUT54), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT126), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1002), .A2(G171), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT125), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1002), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1009), .B(new_n1010), .C1(new_n1015), .C2(new_n1006), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT118), .ZN(new_n1017));
  AND3_X1   g592(.A1(G299), .A2(new_n1017), .A3(KEYINPUT57), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT57), .B1(G299), .B2(new_n1017), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g595(.A(KEYINPUT56), .B(G2072), .Z(new_n1021));
  OR2_X1    g596(.A1(new_n990), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n974), .ZN(new_n1023));
  OR2_X1    g598(.A1(new_n982), .A2(KEYINPUT115), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n982), .A2(KEYINPUT115), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1023), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1020), .B(new_n1022), .C1(G1956), .C2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n592), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1348), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n997), .A2(new_n1030), .A3(new_n998), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n981), .A2(new_n980), .ZN(new_n1032));
  INV_X1    g607(.A(G2067), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AND3_X1   g609(.A1(new_n1031), .A2(KEYINPUT120), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT120), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1020), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1022), .B1(new_n1026), .B2(G1956), .ZN(new_n1039));
  AOI22_X1  g614(.A1(new_n1029), .A2(new_n1037), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1038), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n1027), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT61), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT122), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT122), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1041), .A2(new_n1027), .A3(new_n1045), .A4(KEYINPUT61), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT58), .B(G1341), .ZN(new_n1048));
  OAI22_X1  g623(.A1(new_n990), .A2(G1996), .B1(new_n1032), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n551), .ZN(new_n1050));
  XOR2_X1   g625(.A(new_n1050), .B(KEYINPUT59), .Z(new_n1051));
  XNOR2_X1  g626(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1051), .B1(new_n1042), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1047), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT60), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n1028), .ZN(new_n1056));
  OAI211_X1 g631(.A(KEYINPUT60), .B(new_n592), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT60), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1056), .A2(new_n1057), .B1(new_n1058), .B2(new_n1037), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1040), .B1(new_n1054), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n1061));
  INV_X1    g636(.A(G8), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1061), .B1(G166), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n982), .A2(KEYINPUT115), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n982), .A2(KEYINPUT115), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n764), .B(new_n974), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n990), .A2(new_n688), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1065), .B1(new_n1070), .B2(G8), .ZN(new_n1071));
  NAND2_X1  g646(.A1(G305), .A2(G1981), .ZN(new_n1072));
  INV_X1    g647(.A(G1981), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n571), .A2(new_n1073), .A3(new_n575), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1072), .B(new_n1074), .C1(KEYINPUT114), .C2(KEYINPUT49), .ZN(new_n1075));
  NOR2_X1   g650(.A1(KEYINPUT114), .A2(KEYINPUT49), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1074), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1073), .B1(new_n571), .B2(new_n575), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1032), .A2(new_n1062), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1075), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(G1976), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1080), .B1(G288), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT52), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT52), .B1(G288), .B2(new_n1082), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1085), .B(new_n1080), .C1(new_n1082), .C2(G288), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1081), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n978), .A2(new_n764), .A3(new_n982), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT112), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n978), .A2(KEYINPUT112), .A3(new_n764), .A4(new_n982), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1090), .A2(new_n1069), .A3(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1092), .A2(G8), .A3(new_n1065), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT113), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1092), .A2(KEYINPUT113), .A3(G8), .A4(new_n1065), .ZN(new_n1096));
  AOI211_X1 g671(.A(new_n1071), .B(new_n1087), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n978), .A2(new_n741), .A3(new_n982), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n990), .A2(new_n785), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1062), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(G168), .A2(new_n1062), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1100), .A2(KEYINPUT51), .A3(new_n1101), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1102), .A2(KEYINPUT123), .ZN(new_n1103));
  OAI21_X1  g678(.A(KEYINPUT51), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n1102), .B2(KEYINPUT123), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1100), .ZN(new_n1106));
  OAI22_X1  g681(.A1(new_n1103), .A2(new_n1105), .B1(G168), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1097), .A2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT127), .B1(new_n1002), .B2(G171), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1002), .A2(KEYINPUT127), .A3(G171), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1005), .A2(G171), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(KEYINPUT54), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1108), .B1(new_n1109), .B2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1008), .A2(new_n1016), .A3(new_n1060), .A4(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1087), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1071), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1106), .A2(G286), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT63), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1117), .B1(new_n1097), .B2(new_n1119), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT117), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1116), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT116), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT117), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1126), .A2(new_n1127), .A3(new_n1121), .A4(new_n1120), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1092), .A2(G8), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1129), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1116), .A2(KEYINPUT63), .A3(new_n1119), .A4(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1124), .A2(new_n1128), .A3(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(G288), .A2(G1976), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1081), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1080), .B1(new_n1134), .B2(new_n1077), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1135), .B1(new_n1136), .B2(new_n1087), .ZN(new_n1137));
  XOR2_X1   g712(.A(new_n1107), .B(KEYINPUT62), .Z(new_n1138));
  AND2_X1   g713(.A1(new_n1015), .A2(new_n1097), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1137), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1115), .A2(new_n1132), .A3(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n808), .B(new_n1033), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1142), .B(KEYINPUT110), .ZN(new_n1143));
  INV_X1    g718(.A(new_n987), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n989), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(KEYINPUT109), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n777), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1145), .A2(G1996), .ZN(new_n1150));
  AOI22_X1  g725(.A1(new_n1149), .A2(G1996), .B1(new_n778), .B2(new_n1150), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n1147), .A2(new_n1151), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n709), .A2(new_n711), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n709), .A2(new_n711), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1146), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1145), .ZN(new_n1157));
  XNOR2_X1  g732(.A(G290), .B(G1986), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1156), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1141), .A2(new_n1159), .ZN(new_n1160));
  OR2_X1    g735(.A1(new_n1150), .A2(KEYINPUT46), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1150), .A2(KEYINPUT46), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1147), .A2(new_n1148), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  XOR2_X1   g738(.A(new_n1163), .B(KEYINPUT47), .Z(new_n1164));
  INV_X1    g739(.A(new_n1146), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n803), .A2(new_n1033), .A3(new_n807), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1165), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NOR3_X1   g743(.A1(new_n1145), .A2(G290), .A3(G1986), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1169), .B(KEYINPUT48), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1156), .A2(new_n1170), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n1164), .A2(new_n1168), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1160), .A2(new_n1172), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g748(.A1(G227), .A2(new_n461), .ZN(new_n1175));
  NOR3_X1   g749(.A1(G229), .A2(G401), .A3(new_n1175), .ZN(new_n1176));
  OAI21_X1  g750(.A(new_n1176), .B1(new_n881), .B2(new_n882), .ZN(new_n1177));
  AND2_X1   g751(.A1(new_n968), .A2(new_n969), .ZN(new_n1178));
  AOI21_X1  g752(.A(new_n1177), .B1(new_n963), .B2(new_n1178), .ZN(G308));
  NAND2_X1  g753(.A1(new_n1178), .A2(new_n963), .ZN(new_n1180));
  NAND3_X1  g754(.A1(new_n884), .A2(new_n880), .A3(new_n879), .ZN(new_n1181));
  NAND3_X1  g755(.A1(new_n1180), .A2(new_n1181), .A3(new_n1176), .ZN(G225));
endmodule


