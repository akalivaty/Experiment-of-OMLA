//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n627, new_n628, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1230;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n455), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(G125), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI211_X1 g041(.A(G137), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n461), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n466), .A2(new_n470), .ZN(G160));
  OR2_X1    g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n461), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  XOR2_X1   g049(.A(new_n474), .B(KEYINPUT66), .Z(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  XOR2_X1   g051(.A(new_n476), .B(KEYINPUT67), .Z(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G112), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  AOI21_X1  g055(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(G136), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  OAI211_X1 g059(.A(G126), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n461), .A2(G114), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI211_X1 g063(.A(G138), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n481), .A2(new_n491), .A3(G138), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n488), .B1(new_n490), .B2(new_n492), .ZN(G164));
  INV_X1    g068(.A(KEYINPUT5), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(G543), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n496));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(KEYINPUT5), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n494), .A2(KEYINPUT70), .A3(G543), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n495), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(KEYINPUT68), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(KEYINPUT6), .A3(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  AND2_X1   g081(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G88), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n506), .A2(G50), .A3(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n509), .A2(KEYINPUT69), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(KEYINPUT69), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n508), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n500), .A2(G62), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n502), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n512), .A2(new_n515), .ZN(G166));
  NAND2_X1  g091(.A1(new_n507), .A2(G89), .ZN(new_n517));
  AND2_X1   g092(.A1(G63), .A2(G651), .ZN(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n519), .A2(KEYINPUT7), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(KEYINPUT7), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n500), .A2(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n497), .B1(new_n506), .B2(KEYINPUT71), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT71), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n503), .A2(new_n525), .A3(new_n505), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n523), .A2(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  NAND2_X1  g105(.A1(new_n524), .A2(new_n526), .ZN(new_n531));
  INV_X1    g106(.A(G52), .ZN(new_n532));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n500), .A2(new_n506), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n531), .A2(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n500), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n502), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n535), .A2(new_n537), .ZN(G171));
  AND3_X1   g113(.A1(new_n504), .A2(KEYINPUT6), .A3(G651), .ZN(new_n539));
  AOI21_X1  g114(.A(KEYINPUT6), .B1(new_n504), .B2(G651), .ZN(new_n540));
  OAI21_X1  g115(.A(KEYINPUT71), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  XOR2_X1   g116(.A(KEYINPUT72), .B(G43), .Z(new_n542));
  NAND4_X1  g117(.A1(new_n541), .A2(G543), .A3(new_n526), .A4(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n500), .A2(G81), .A3(new_n506), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n500), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n543), .B(new_n544), .C1(new_n545), .C2(new_n502), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT73), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n498), .A2(new_n499), .ZN(new_n549));
  INV_X1    g124(.A(new_n495), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n549), .A2(G56), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G651), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n554), .A2(KEYINPUT73), .A3(new_n543), .A4(new_n544), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n548), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n549), .A2(new_n550), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT74), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n566), .A2(new_n567), .A3(G651), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n500), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT74), .B1(new_n569), .B2(new_n502), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n524), .A2(G53), .A3(new_n526), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(KEYINPUT9), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n524), .A2(new_n574), .A3(G53), .A4(new_n526), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n507), .A2(G91), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n571), .A2(new_n576), .A3(new_n577), .ZN(G299));
  INV_X1    g153(.A(G171), .ZN(G301));
  XNOR2_X1  g154(.A(new_n509), .B(KEYINPUT69), .ZN(new_n580));
  INV_X1    g155(.A(new_n515), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n580), .A2(new_n581), .A3(new_n508), .ZN(G303));
  OAI21_X1  g157(.A(G651), .B1(new_n500), .B2(G74), .ZN(new_n583));
  INV_X1    g158(.A(G87), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n584), .B2(new_n534), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n541), .A2(G49), .A3(G543), .A4(new_n526), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(KEYINPUT75), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT75), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n524), .A2(new_n588), .A3(G49), .A4(new_n526), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n585), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G288));
  AOI22_X1  g166(.A1(new_n500), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n502), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n506), .A2(G48), .A3(G543), .ZN(new_n594));
  INV_X1    g169(.A(G86), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n534), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(new_n507), .A2(G85), .ZN(new_n599));
  INV_X1    g174(.A(G47), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(new_n531), .ZN(new_n601));
  NAND2_X1  g176(.A1(G72), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G60), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n564), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G651), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(KEYINPUT76), .B1(new_n601), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n527), .A2(G47), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT76), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n608), .A2(new_n609), .A3(new_n605), .A4(new_n599), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n607), .A2(new_n610), .ZN(G290));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n564), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n527), .A2(G54), .B1(new_n614), .B2(G651), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n500), .A2(G92), .A3(new_n506), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT10), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(G868), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(new_n620), .B2(G171), .ZN(G284));
  OAI21_X1  g197(.A(new_n621), .B1(new_n620), .B2(G171), .ZN(G321));
  NAND2_X1  g198(.A1(G299), .A2(new_n620), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(new_n620), .B2(G168), .ZN(G297));
  XNOR2_X1  g200(.A(G297), .B(KEYINPUT77), .ZN(G280));
  INV_X1    g201(.A(new_n619), .ZN(new_n627));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(G860), .ZN(G148));
  NAND2_X1  g204(.A1(new_n556), .A2(new_n620), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n619), .A2(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(new_n620), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g208(.A1(new_n472), .A2(new_n473), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(new_n468), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n638), .A2(G2100), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n475), .A2(G123), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n461), .A2(G111), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(KEYINPUT78), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(new_n641), .B2(KEYINPUT78), .ZN(new_n644));
  AOI22_X1  g219(.A1(new_n642), .A2(new_n644), .B1(new_n481), .B2(G135), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n640), .A2(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n646), .A2(G2096), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n638), .A2(G2100), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(G2096), .ZN(new_n649));
  NAND4_X1  g224(.A1(new_n639), .A2(new_n647), .A3(new_n648), .A4(new_n649), .ZN(G156));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT79), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2427), .B(G2430), .Z(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(KEYINPUT14), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2443), .B(G2446), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2451), .B(G2454), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT80), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n659), .A2(new_n662), .ZN(new_n664));
  AND2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1341), .B(G1348), .ZN(new_n666));
  OAI21_X1  g241(.A(G14), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n663), .A2(new_n666), .A3(new_n664), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(KEYINPUT81), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(KEYINPUT81), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n667), .B1(new_n669), .B2(new_n670), .ZN(G401));
  XNOR2_X1  g246(.A(G2072), .B(G2078), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT17), .Z(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2084), .B(G2090), .Z(new_n677));
  INV_X1    g252(.A(new_n672), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n677), .B1(new_n675), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n676), .B1(KEYINPUT82), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(KEYINPUT82), .B2(new_n679), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n677), .A2(new_n674), .A3(new_n672), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT18), .Z(new_n683));
  NAND3_X1  g258(.A1(new_n673), .A2(new_n677), .A3(new_n675), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n681), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G2096), .B(G2100), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT83), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n685), .B(new_n687), .ZN(G227));
  XOR2_X1   g263(.A(G1971), .B(G1976), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  XOR2_X1   g265(.A(G1956), .B(G2474), .Z(new_n691));
  XOR2_X1   g266(.A(G1961), .B(G1966), .Z(new_n692));
  AND2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT84), .B(KEYINPUT20), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n691), .A2(new_n692), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  MUX2_X1   g273(.A(new_n698), .B(new_n697), .S(new_n690), .Z(new_n699));
  NOR2_X1   g274(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT85), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n700), .B(new_n702), .Z(new_n703));
  XNOR2_X1  g278(.A(G1991), .B(G1996), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1981), .B(G1986), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(G229));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G21), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G168), .B2(new_n709), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT92), .ZN(new_n712));
  INV_X1    g287(.A(G1966), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT94), .Z(new_n715));
  NOR2_X1   g290(.A1(new_n712), .A2(new_n713), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT93), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n709), .A2(G19), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT88), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(new_n557), .B2(new_n709), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT89), .B(G1341), .Z(new_n722));
  OR2_X1    g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n709), .A2(G20), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT23), .Z(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G299), .B2(G16), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT95), .B(G1956), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n721), .A2(new_n722), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n723), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G29), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G32), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n475), .A2(G129), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n468), .A2(G105), .ZN(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT26), .ZN(new_n737));
  AOI211_X1 g312(.A(new_n735), .B(new_n737), .C1(G141), .C2(new_n481), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n733), .B1(new_n740), .B2(new_n732), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT91), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT27), .B(G1996), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n742), .B(new_n743), .Z(new_n744));
  NAND2_X1  g319(.A1(new_n732), .A2(G26), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT28), .Z(new_n746));
  NAND2_X1  g321(.A1(new_n475), .A2(G128), .ZN(new_n747));
  OAI21_X1  g322(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n748));
  INV_X1    g323(.A(G116), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(G2105), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G140), .B2(new_n481), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n746), .B1(new_n752), .B2(G29), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G2067), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT31), .B(G11), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT30), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n756), .A2(G28), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n732), .B1(new_n756), .B2(G28), .ZN(new_n758));
  OAI221_X1 g333(.A(new_n755), .B1(new_n757), .B2(new_n758), .C1(new_n646), .C2(new_n732), .ZN(new_n759));
  OAI21_X1  g334(.A(G29), .B1(new_n466), .B2(new_n470), .ZN(new_n760));
  INV_X1    g335(.A(G2084), .ZN(new_n761));
  INV_X1    g336(.A(G34), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n762), .A2(KEYINPUT24), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n762), .A2(KEYINPUT24), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n732), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AND3_X1   g340(.A1(new_n760), .A2(new_n761), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n761), .B1(new_n760), .B2(new_n765), .ZN(new_n767));
  NOR3_X1   g342(.A1(new_n759), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(G27), .A2(G29), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G164), .B2(G29), .ZN(new_n770));
  INV_X1    g345(.A(G2078), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n732), .A2(G33), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n481), .A2(G139), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT90), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT25), .Z(new_n777));
  AOI22_X1  g352(.A1(new_n634), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(new_n778), .B2(new_n461), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n773), .B1(new_n780), .B2(new_n732), .ZN(new_n781));
  INV_X1    g356(.A(G2072), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n754), .A2(new_n768), .A3(new_n772), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n709), .A2(G4), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n627), .B2(new_n709), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G1348), .ZN(new_n787));
  NOR3_X1   g362(.A1(new_n744), .A2(new_n784), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(G29), .A2(G35), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G162), .B2(G29), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT29), .B(G2090), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n726), .A2(new_n727), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n709), .A2(G5), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G171), .B2(new_n709), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G1961), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n792), .A2(new_n793), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n718), .A2(new_n731), .A3(new_n788), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n732), .A2(G25), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n475), .A2(G119), .ZN(new_n800));
  OAI21_X1  g375(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n801));
  INV_X1    g376(.A(G107), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(G2105), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G131), .B2(new_n481), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n799), .B1(new_n806), .B2(new_n732), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT35), .B(G1991), .Z(new_n808));
  XOR2_X1   g383(.A(new_n807), .B(new_n808), .Z(new_n809));
  MUX2_X1   g384(.A(G24), .B(G290), .S(G16), .Z(new_n810));
  AOI21_X1  g385(.A(new_n809), .B1(G1986), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G1986), .B2(new_n810), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n709), .A2(G22), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G166), .B2(new_n709), .ZN(new_n814));
  INV_X1    g389(.A(G1971), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n709), .A2(G23), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n590), .B2(new_n709), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT33), .B(G1976), .Z(new_n819));
  OR2_X1    g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n709), .A2(G6), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n597), .B2(new_n709), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT32), .B(G1981), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT86), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n823), .B(new_n825), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n816), .A2(new_n820), .A3(new_n821), .A4(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n827), .A2(KEYINPUT34), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n812), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(KEYINPUT34), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT87), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(KEYINPUT36), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT36), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n829), .A2(new_n834), .A3(new_n831), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n798), .B1(new_n833), .B2(new_n835), .ZN(G311));
  INV_X1    g411(.A(new_n798), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n833), .A2(new_n835), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(G150));
  NAND2_X1  g414(.A1(new_n627), .A2(G559), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT99), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT38), .ZN(new_n842));
  INV_X1    g417(.A(G55), .ZN(new_n843));
  INV_X1    g418(.A(G93), .ZN(new_n844));
  OAI22_X1  g419(.A1(new_n531), .A2(new_n843), .B1(new_n844), .B2(new_n534), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n549), .A2(G67), .A3(new_n550), .ZN(new_n846));
  NAND2_X1  g421(.A1(G80), .A2(G543), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT96), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n847), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(new_n500), .B2(G67), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(KEYINPUT96), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n850), .A2(G651), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n845), .B1(new_n854), .B2(KEYINPUT97), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT97), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n850), .A2(new_n853), .A3(new_n856), .A4(G651), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n556), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(G651), .B1(new_n852), .B2(KEYINPUT96), .ZN(new_n859));
  AOI211_X1 g434(.A(new_n849), .B(new_n851), .C1(new_n500), .C2(G67), .ZN(new_n860));
  OAI21_X1  g435(.A(KEYINPUT97), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AOI22_X1  g436(.A1(new_n527), .A2(G55), .B1(G93), .B2(new_n507), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n861), .A2(new_n857), .A3(new_n862), .A4(new_n546), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(KEYINPUT98), .B1(new_n858), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT98), .ZN(new_n866));
  AND3_X1   g441(.A1(new_n861), .A2(new_n857), .A3(new_n862), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n866), .B(new_n863), .C1(new_n867), .C2(new_n556), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n842), .A2(new_n869), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n841), .A2(KEYINPUT38), .ZN(new_n871));
  INV_X1    g446(.A(new_n869), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n841), .A2(KEYINPUT38), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n870), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(G860), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n875), .B1(new_n870), .B2(new_n874), .ZN(new_n879));
  OAI21_X1  g454(.A(KEYINPUT100), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n879), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT100), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n881), .A2(new_n882), .A3(new_n877), .A4(new_n876), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n861), .A2(new_n857), .A3(new_n862), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(G860), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n886), .B(KEYINPUT37), .Z(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n887), .ZN(G145));
  XNOR2_X1  g463(.A(new_n805), .B(new_n636), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n475), .A2(G130), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT102), .ZN(new_n892));
  OAI21_X1  g467(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n893));
  INV_X1    g468(.A(G118), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n893), .B1(new_n894), .B2(G2105), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n895), .B1(G142), .B2(new_n481), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n890), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n889), .A2(new_n892), .A3(new_n896), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n752), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n740), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n739), .A2(new_n752), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(G164), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n492), .A2(new_n490), .ZN(new_n907));
  INV_X1    g482(.A(new_n488), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n903), .A2(new_n909), .A3(new_n904), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n780), .B(KEYINPUT101), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n906), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n780), .A2(KEYINPUT101), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n914), .B1(new_n906), .B2(new_n910), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n901), .B(KEYINPUT103), .C1(new_n913), .C2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n898), .A2(new_n899), .A3(KEYINPUT103), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n906), .A2(new_n910), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n917), .B(new_n912), .C1(new_n918), .C2(new_n914), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n646), .B(G160), .ZN(new_n920));
  XOR2_X1   g495(.A(new_n483), .B(new_n920), .Z(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n916), .A2(new_n919), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(G37), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n913), .A2(new_n915), .A3(new_n900), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n900), .B1(new_n913), .B2(new_n915), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(new_n921), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n923), .B(new_n924), .C1(new_n925), .C2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n928), .B(new_n929), .ZN(G395));
  OR2_X1    g505(.A1(new_n869), .A2(new_n631), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n869), .A2(new_n631), .ZN(new_n932));
  NAND2_X1  g507(.A1(G299), .A2(new_n619), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT41), .ZN(new_n934));
  AOI22_X1  g509(.A1(new_n573), .A2(new_n575), .B1(G91), .B2(new_n507), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n935), .A2(new_n571), .A3(new_n618), .A4(new_n615), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n933), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT105), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT105), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n933), .A2(new_n939), .A3(new_n936), .A4(new_n934), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n933), .A2(new_n936), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n938), .B(new_n940), .C1(new_n942), .C2(new_n943), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n931), .A2(new_n932), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n941), .B1(new_n931), .B2(new_n932), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(new_n512), .B2(new_n515), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n580), .A2(new_n581), .A3(KEYINPUT107), .A4(new_n508), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(G288), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(G288), .B1(new_n949), .B2(new_n950), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n607), .A2(G305), .A3(new_n610), .ZN(new_n954));
  AOI21_X1  g529(.A(G305), .B1(new_n607), .B2(new_n610), .ZN(new_n955));
  OAI22_X1  g530(.A1(new_n952), .A2(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(G290), .A2(new_n597), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n949), .A2(new_n950), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n590), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n607), .A2(G305), .A3(new_n610), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n957), .A2(new_n959), .A3(new_n960), .A4(new_n951), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n956), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g537(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n963));
  XNOR2_X1  g538(.A(new_n962), .B(new_n963), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n947), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n947), .A2(new_n964), .ZN(new_n966));
  OAI21_X1  g541(.A(G868), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(G868), .B2(new_n867), .ZN(G295));
  OAI21_X1  g543(.A(new_n967), .B1(G868), .B2(new_n867), .ZN(G331));
  INV_X1    g544(.A(new_n868), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n885), .A2(new_n548), .A3(new_n555), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n866), .B1(new_n971), .B2(new_n863), .ZN(new_n972));
  XNOR2_X1  g547(.A(G286), .B(G171), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n970), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n973), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n975), .B1(new_n865), .B2(new_n868), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n944), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n973), .B1(new_n970), .B2(new_n972), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n865), .A2(new_n868), .A3(new_n975), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(new_n942), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n977), .A2(new_n962), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n924), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n962), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n956), .A2(new_n961), .A3(KEYINPUT109), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n941), .A2(new_n934), .ZN(new_n987));
  INV_X1    g562(.A(new_n943), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n942), .A2(new_n988), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n987), .B(new_n989), .C1(new_n974), .C2(new_n976), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n986), .B1(new_n980), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT110), .B1(new_n982), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n985), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT109), .B1(new_n956), .B2(new_n961), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n980), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n989), .A2(new_n987), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n997), .B1(new_n978), .B2(new_n979), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n995), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT110), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n999), .A2(new_n1000), .A3(new_n981), .A4(new_n924), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n992), .A2(KEYINPUT43), .A3(new_n1001), .ZN(new_n1002));
  AOI22_X1  g577(.A1(new_n937), .A2(KEYINPUT105), .B1(new_n941), .B2(new_n988), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n978), .A2(new_n979), .B1(new_n940), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n995), .B1(new_n996), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT43), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1005), .A2(new_n1006), .A3(new_n924), .A4(new_n981), .ZN(new_n1007));
  AND2_X1   g582(.A1(new_n1007), .A2(KEYINPUT44), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1002), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n986), .B1(new_n977), .B2(new_n980), .ZN(new_n1010));
  OAI21_X1  g585(.A(KEYINPUT43), .B1(new_n982), .B2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n999), .A2(new_n1006), .A3(new_n981), .A4(new_n924), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT44), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1009), .A2(new_n1015), .ZN(G397));
  OR2_X1    g591(.A1(G290), .A2(G1986), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n467), .A2(new_n469), .ZN(new_n1018));
  INV_X1    g593(.A(G125), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1019), .B1(new_n472), .B2(new_n473), .ZN(new_n1020));
  INV_X1    g595(.A(new_n465), .ZN(new_n1021));
  OAI21_X1  g596(.A(G2105), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1018), .A2(new_n1022), .A3(G40), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT111), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(G160), .A2(KEYINPUT111), .A3(G40), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT45), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(G164), .B2(G1384), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  OR2_X1    g606(.A1(new_n1017), .A2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1033));
  INV_X1    g608(.A(G2067), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n752), .B(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1996), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n739), .B(new_n1036), .ZN(new_n1037));
  OR2_X1    g612(.A1(new_n806), .A2(new_n808), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n806), .A2(new_n808), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1035), .A2(new_n1037), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n1032), .A2(new_n1033), .B1(new_n1040), .B2(new_n1030), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1042));
  AND4_X1   g617(.A1(new_n808), .A2(new_n1035), .A3(new_n1037), .A4(new_n806), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1043), .B1(new_n1034), .B2(new_n902), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1042), .B1(new_n1031), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1030), .A2(new_n1036), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n1046), .B(KEYINPUT46), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n1035), .A2(new_n740), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1047), .B1(new_n1048), .B2(new_n1031), .ZN(new_n1049));
  XOR2_X1   g624(.A(new_n1049), .B(KEYINPUT125), .Z(new_n1050));
  INV_X1    g625(.A(KEYINPUT47), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1045), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n587), .A2(new_n589), .ZN(new_n1055));
  INV_X1    g630(.A(new_n585), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .A4(G1976), .ZN(new_n1058));
  AOI21_X1  g633(.A(G1384), .B1(new_n907), .B2(new_n908), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1025), .A2(new_n1059), .A3(new_n1026), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1058), .A2(G8), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1057), .B1(new_n590), .B2(G1976), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G1976), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT52), .B1(G288), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1061), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT115), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1061), .A2(new_n1063), .A3(new_n1065), .A4(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g644(.A(KEYINPUT117), .B(G86), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n594), .B1(new_n534), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(G1981), .B1(new_n593), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G1981), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT116), .B1(new_n597), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n1075));
  NOR4_X1   g650(.A1(new_n593), .A2(new_n596), .A3(new_n1075), .A4(G1981), .ZN(new_n1076));
  OAI211_X1 g651(.A(KEYINPUT49), .B(new_n1072), .C1(new_n1074), .C2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1060), .A2(G8), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1072), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT49), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1078), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1067), .A2(new_n1069), .B1(new_n1077), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G1384), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n909), .A2(KEYINPUT45), .A3(new_n1083), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1029), .A2(new_n1084), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT50), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n909), .A2(new_n1088), .A3(new_n1083), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1087), .A2(new_n1089), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1090));
  XOR2_X1   g665(.A(KEYINPUT112), .B(G2090), .Z(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  OAI22_X1  g667(.A1(new_n1086), .A2(G1971), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT55), .ZN(new_n1094));
  INV_X1    g669(.A(G8), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1094), .B1(G166), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1093), .A2(new_n1098), .A3(KEYINPUT119), .A4(G8), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n1095), .A2(KEYINPUT119), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1096), .A2(new_n1097), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1090), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1102), .A2(new_n1091), .B1(new_n815), .B2(new_n1085), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1101), .B1(new_n1103), .B2(new_n1095), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1099), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1058), .A2(G8), .A3(new_n1060), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT52), .B1(new_n1106), .B2(new_n1062), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT114), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT114), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1109), .B(KEYINPUT52), .C1(new_n1106), .C2(new_n1062), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(G168), .A2(G8), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1087), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1113), .A2(KEYINPUT120), .A3(new_n761), .A4(new_n1089), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1085), .A2(new_n713), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT120), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(new_n1090), .B2(G2084), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1112), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1082), .A2(new_n1105), .A3(new_n1111), .A4(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT63), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT121), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1098), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1124), .A2(G8), .A3(new_n1093), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1098), .B(new_n1123), .C1(new_n1103), .C2(new_n1095), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1119), .A2(new_n1125), .A3(KEYINPUT63), .A4(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1082), .A2(new_n1111), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1103), .A2(new_n1098), .A3(new_n1095), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1081), .A2(new_n1077), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1130), .A2(new_n1131), .A3(new_n1111), .A4(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n590), .A2(new_n1064), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1134), .B1(new_n1081), .B2(new_n1077), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1136));
  OAI211_X1 g711(.A(G8), .B(new_n1060), .C1(new_n1135), .C2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT118), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1133), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1138), .B1(new_n1133), .B2(new_n1137), .ZN(new_n1140));
  OAI22_X1  g715(.A1(new_n1122), .A2(new_n1129), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(KEYINPUT122), .B(KEYINPUT57), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n935), .A2(new_n571), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1142), .B1(new_n935), .B2(new_n571), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(G1956), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1090), .A2(new_n1147), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1149));
  XNOR2_X1  g724(.A(KEYINPUT123), .B(KEYINPUT56), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1150), .B(new_n782), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1149), .A2(new_n1029), .A3(new_n1084), .A4(new_n1151), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1146), .A2(KEYINPUT124), .A3(new_n1148), .A4(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1142), .ZN(new_n1154));
  NAND2_X1  g729(.A1(G299), .A2(new_n1154), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1148), .A2(new_n1155), .A3(new_n1152), .A4(new_n1143), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1153), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1148), .A2(new_n1152), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1155), .A2(new_n1143), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(KEYINPUT61), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(G1348), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1090), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1060), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(new_n1034), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1165), .A2(new_n619), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n619), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1169));
  OAI21_X1  g744(.A(KEYINPUT60), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1162), .A2(KEYINPUT61), .A3(new_n1156), .ZN(new_n1171));
  XOR2_X1   g746(.A(KEYINPUT58), .B(G1341), .Z(new_n1172));
  NAND2_X1  g747(.A1(new_n1060), .A2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1173), .B1(new_n1085), .B2(G1996), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(new_n557), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT59), .ZN(new_n1176));
  AOI22_X1  g751(.A1(new_n1090), .A2(new_n1164), .B1(new_n1166), .B2(new_n1034), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n619), .A2(KEYINPUT60), .ZN(new_n1178));
  AOI22_X1  g753(.A1(new_n1175), .A2(new_n1176), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1174), .A2(KEYINPUT59), .A3(new_n557), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1170), .A2(new_n1171), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1159), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1169), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1183));
  OAI22_X1  g758(.A1(new_n1163), .A2(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(G168), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1114), .A2(new_n1118), .A3(G168), .A4(new_n1115), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(G8), .ZN(new_n1187));
  OAI21_X1  g762(.A(KEYINPUT51), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1188));
  AND2_X1   g763(.A1(new_n1186), .A2(G8), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT51), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1188), .A2(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g767(.A(G171), .B(KEYINPUT54), .ZN(new_n1193));
  AOI21_X1  g768(.A(KEYINPUT53), .B1(new_n1086), .B2(new_n771), .ZN(new_n1194));
  INV_X1    g769(.A(G1961), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1194), .B1(new_n1195), .B2(new_n1090), .ZN(new_n1196));
  AND2_X1   g771(.A1(new_n771), .A2(KEYINPUT53), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1086), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1193), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1023), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1029), .A2(new_n1084), .A3(new_n1200), .A4(new_n1197), .ZN(new_n1201));
  AND2_X1   g776(.A1(new_n1193), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1199), .B1(new_n1196), .B2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1184), .A2(new_n1192), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1205));
  INV_X1    g780(.A(new_n1118), .ZN(new_n1206));
  OAI21_X1  g781(.A(G286), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1190), .B1(new_n1189), .B2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g783(.A1(new_n1187), .A2(KEYINPUT51), .ZN(new_n1209));
  OAI21_X1  g784(.A(KEYINPUT62), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT62), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1188), .A2(new_n1211), .A3(new_n1191), .ZN(new_n1212));
  AOI21_X1  g787(.A(G301), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1210), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1204), .A2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1128), .B1(new_n1104), .B2(new_n1099), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1141), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1040), .B1(G1986), .B2(G290), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1031), .B1(new_n1218), .B2(new_n1017), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1054), .B1(new_n1217), .B2(new_n1219), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g795(.A1(G227), .A2(new_n459), .ZN(new_n1222));
  INV_X1    g796(.A(new_n1222), .ZN(new_n1223));
  OAI21_X1  g797(.A(KEYINPUT127), .B1(G401), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g798(.A(KEYINPUT127), .ZN(new_n1225));
  AND2_X1   g799(.A1(new_n670), .A2(new_n669), .ZN(new_n1226));
  OAI211_X1 g800(.A(new_n1225), .B(new_n1222), .C1(new_n1226), .C2(new_n667), .ZN(new_n1227));
  NAND4_X1  g801(.A1(new_n928), .A2(new_n1224), .A3(new_n1227), .A4(new_n707), .ZN(new_n1228));
  AOI21_X1  g802(.A(new_n1228), .B1(new_n1011), .B2(new_n1012), .ZN(G308));
  AND2_X1   g803(.A1(new_n1224), .A2(new_n707), .ZN(new_n1230));
  NAND4_X1  g804(.A1(new_n1230), .A2(new_n1013), .A3(new_n928), .A4(new_n1227), .ZN(G225));
endmodule


