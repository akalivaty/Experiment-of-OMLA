

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748;

  NOR2_X1 U371 ( .A1(n586), .A2(n585), .ZN(n643) );
  AND2_X2 U372 ( .A1(n359), .A2(n620), .ZN(n621) );
  NOR2_X2 U373 ( .A1(n404), .A2(n438), .ZN(n379) );
  NOR2_X1 U374 ( .A1(n411), .A2(n668), .ZN(n390) );
  XNOR2_X2 U375 ( .A(n420), .B(n419), .ZN(n554) );
  NOR2_X1 U376 ( .A1(n686), .A2(n608), .ZN(n609) );
  XNOR2_X2 U377 ( .A(n509), .B(n412), .ZN(n544) );
  INV_X1 U378 ( .A(KEYINPUT4), .ZN(n444) );
  XOR2_X1 U379 ( .A(G143), .B(G128), .Z(n529) );
  OR2_X1 U380 ( .A1(n613), .A2(n440), .ZN(n437) );
  NOR2_X1 U381 ( .A1(n600), .A2(n599), .ZN(n613) );
  OR2_X1 U382 ( .A1(n612), .A2(n440), .ZN(n434) );
  NAND2_X1 U383 ( .A1(n361), .A2(n360), .ZN(n747) );
  XNOR2_X1 U384 ( .A(n606), .B(n605), .ZN(n380) );
  XNOR2_X1 U385 ( .A(n390), .B(KEYINPUT31), .ZN(n649) );
  XNOR2_X1 U386 ( .A(n601), .B(n405), .ZN(n672) );
  XNOR2_X1 U387 ( .A(n588), .B(KEYINPUT19), .ZN(n570) );
  BUF_X1 U388 ( .A(n558), .Z(n601) );
  XNOR2_X1 U389 ( .A(n394), .B(KEYINPUT69), .ZN(n656) );
  NOR2_X1 U390 ( .A1(n658), .A2(n659), .ZN(n394) );
  NOR2_X2 U391 ( .A1(G902), .A2(n699), .ZN(n455) );
  XNOR2_X1 U392 ( .A(n732), .B(n448), .ZN(n385) );
  XNOR2_X1 U393 ( .A(n446), .B(n529), .ZN(n732) );
  XNOR2_X1 U394 ( .A(n479), .B(n395), .ZN(n495) );
  XNOR2_X1 U395 ( .A(n445), .B(n444), .ZN(n446) );
  NOR2_X2 U396 ( .A1(n678), .A2(n411), .ZN(n512) );
  XNOR2_X2 U397 ( .A(n484), .B(n483), .ZN(n678) );
  XNOR2_X1 U398 ( .A(n366), .B(n611), .ZN(n612) );
  NOR2_X1 U399 ( .A1(n380), .A2(n746), .ZN(n366) );
  INV_X1 U400 ( .A(KEYINPUT78), .ZN(n419) );
  AND2_X1 U401 ( .A1(n613), .A2(n439), .ZN(n438) );
  AND2_X1 U402 ( .A1(n406), .A2(n631), .ZN(n357) );
  NAND2_X1 U403 ( .A1(n372), .A2(n376), .ZN(n371) );
  AND2_X1 U404 ( .A1(n349), .A2(n747), .ZN(n356) );
  XNOR2_X1 U405 ( .A(n381), .B(n350), .ZN(n546) );
  OR2_X1 U406 ( .A1(n624), .A2(G902), .ZN(n381) );
  INV_X1 U407 ( .A(KEYINPUT0), .ZN(n412) );
  NAND2_X1 U408 ( .A1(n570), .A2(n508), .ZN(n509) );
  XOR2_X1 U409 ( .A(G478), .B(n538), .Z(n552) );
  AND2_X1 U410 ( .A1(n375), .A2(n417), .ZN(n374) );
  NAND2_X1 U411 ( .A1(n377), .A2(n376), .ZN(n375) );
  INV_X1 U412 ( .A(n634), .ZN(n377) );
  XNOR2_X1 U413 ( .A(G131), .B(G137), .ZN(n449) );
  NAND2_X1 U414 ( .A1(n672), .A2(n671), .ZN(n369) );
  NOR2_X1 U415 ( .A1(n438), .A2(n431), .ZN(n615) );
  AND2_X1 U416 ( .A1(n434), .A2(n433), .ZN(n435) );
  NOR2_X1 U417 ( .A1(n654), .A2(n436), .ZN(n433) );
  INV_X1 U418 ( .A(KEYINPUT28), .ZN(n364) );
  XNOR2_X1 U419 ( .A(n482), .B(n476), .ZN(n382) );
  XNOR2_X1 U420 ( .A(n495), .B(n481), .ZN(n482) );
  XNOR2_X1 U421 ( .A(G953), .B(KEYINPUT64), .ZN(n561) );
  AND2_X1 U422 ( .A1(n434), .A2(n432), .ZN(n362) );
  INV_X1 U423 ( .A(n654), .ZN(n432) );
  NAND2_X1 U424 ( .A1(n400), .A2(n407), .ZN(n408) );
  AND2_X1 U425 ( .A1(n358), .A2(n357), .ZN(n400) );
  XOR2_X1 U426 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n531) );
  XNOR2_X1 U427 ( .A(G116), .B(G134), .ZN(n530) );
  XNOR2_X1 U428 ( .A(n529), .B(n392), .ZN(n533) );
  XNOR2_X1 U429 ( .A(G107), .B(G122), .ZN(n392) );
  XNOR2_X1 U430 ( .A(n527), .B(n526), .ZN(n706) );
  XNOR2_X1 U431 ( .A(n383), .B(n604), .ZN(n614) );
  NOR2_X1 U432 ( .A1(n602), .A2(n603), .ZN(n383) );
  XNOR2_X1 U433 ( .A(n422), .B(KEYINPUT109), .ZN(n587) );
  NAND2_X1 U434 ( .A1(n348), .A2(n355), .ZN(n388) );
  BUF_X1 U435 ( .A(n546), .Z(n663) );
  AND2_X1 U436 ( .A1(n607), .A2(n542), .ZN(n543) );
  XNOR2_X1 U437 ( .A(n663), .B(n424), .ZN(n568) );
  INV_X1 U438 ( .A(KEYINPUT6), .ZN(n424) );
  XNOR2_X1 U439 ( .A(n472), .B(n471), .ZN(n473) );
  INV_X1 U440 ( .A(KEYINPUT1), .ZN(n401) );
  NOR2_X1 U441 ( .A1(n741), .A2(G952), .ZN(n719) );
  INV_X1 U442 ( .A(KEYINPUT48), .ZN(n440) );
  INV_X1 U443 ( .A(KEYINPUT98), .ZN(n376) );
  INV_X1 U444 ( .A(n738), .ZN(n436) );
  XNOR2_X1 U445 ( .A(n459), .B(n488), .ZN(n516) );
  XOR2_X1 U446 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n521) );
  XNOR2_X1 U447 ( .A(G143), .B(G140), .ZN(n520) );
  XNOR2_X1 U448 ( .A(KEYINPUT12), .B(KEYINPUT102), .ZN(n522) );
  XOR2_X1 U449 ( .A(KEYINPUT11), .B(KEYINPUT99), .Z(n523) );
  XNOR2_X1 U450 ( .A(n385), .B(n450), .ZN(n477) );
  XOR2_X1 U451 ( .A(KEYINPUT72), .B(G140), .Z(n460) );
  INV_X1 U452 ( .A(KEYINPUT38), .ZN(n405) );
  XNOR2_X1 U453 ( .A(n426), .B(n425), .ZN(n551) );
  XNOR2_X1 U454 ( .A(n528), .B(G475), .ZN(n425) );
  OR2_X1 U455 ( .A1(n706), .A2(G902), .ZN(n426) );
  XOR2_X1 U456 ( .A(KEYINPUT76), .B(KEYINPUT16), .Z(n493) );
  XNOR2_X1 U457 ( .A(G122), .B(KEYINPUT77), .ZN(n492) );
  INV_X1 U458 ( .A(KEYINPUT73), .ZN(n395) );
  INV_X1 U459 ( .A(G953), .ZN(n723) );
  XNOR2_X1 U460 ( .A(G137), .B(KEYINPUT81), .ZN(n463) );
  XNOR2_X1 U461 ( .A(G119), .B(G128), .ZN(n461) );
  XNOR2_X1 U462 ( .A(n516), .B(n460), .ZN(n733) );
  XNOR2_X1 U463 ( .A(G146), .B(G125), .ZN(n488) );
  XOR2_X1 U464 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n487) );
  NAND2_X1 U465 ( .A1(n621), .A2(n379), .ZN(n370) );
  NAND2_X1 U466 ( .A1(n617), .A2(n618), .ZN(n430) );
  XNOR2_X1 U467 ( .A(n393), .B(KEYINPUT41), .ZN(n686) );
  AND2_X1 U468 ( .A1(n672), .A2(n367), .ZN(n393) );
  NOR2_X1 U469 ( .A1(n674), .A2(n368), .ZN(n367) );
  XNOR2_X1 U470 ( .A(n575), .B(KEYINPUT112), .ZN(n608) );
  XNOR2_X1 U471 ( .A(n365), .B(n364), .ZN(n574) );
  XNOR2_X1 U472 ( .A(n536), .B(n391), .ZN(n713) );
  XNOR2_X1 U473 ( .A(n535), .B(n537), .ZN(n391) );
  XNOR2_X1 U474 ( .A(n706), .B(n705), .ZN(n707) );
  AND2_X1 U475 ( .A1(n427), .A2(n583), .ZN(n654) );
  XNOR2_X1 U476 ( .A(n428), .B(KEYINPUT43), .ZN(n427) );
  NOR2_X1 U477 ( .A1(n591), .A2(n368), .ZN(n429) );
  XNOR2_X1 U478 ( .A(KEYINPUT113), .B(KEYINPUT40), .ZN(n605) );
  XNOR2_X1 U479 ( .A(KEYINPUT36), .B(KEYINPUT90), .ZN(n589) );
  NAND2_X1 U480 ( .A1(n387), .A2(n386), .ZN(n360) );
  AND2_X1 U481 ( .A1(n389), .A2(n388), .ZN(n361) );
  NOR2_X1 U482 ( .A1(n348), .A2(n355), .ZN(n386) );
  INV_X1 U483 ( .A(n663), .ZN(n410) );
  NAND2_X1 U484 ( .A1(n556), .A2(n414), .ZN(n413) );
  INV_X1 U485 ( .A(n568), .ZN(n414) );
  XNOR2_X1 U486 ( .A(n695), .B(n694), .ZN(n696) );
  OR2_X1 U487 ( .A1(n353), .A2(n568), .ZN(n348) );
  AND2_X1 U488 ( .A1(n639), .A2(n550), .ZN(n349) );
  INV_X1 U489 ( .A(n675), .ZN(n417) );
  XOR2_X1 U490 ( .A(G472), .B(KEYINPUT75), .Z(n350) );
  XOR2_X1 U491 ( .A(KEYINPUT3), .B(G119), .Z(n351) );
  AND2_X1 U492 ( .A1(n634), .A2(KEYINPUT98), .ZN(n352) );
  OR2_X1 U493 ( .A1(n655), .A2(n567), .ZN(n353) );
  NOR2_X1 U494 ( .A1(n656), .A2(n572), .ZN(n354) );
  INV_X1 U495 ( .A(n671), .ZN(n368) );
  INV_X1 U496 ( .A(n423), .ZN(n644) );
  OR2_X1 U497 ( .A1(n553), .A2(n552), .ZN(n423) );
  XOR2_X1 U498 ( .A(KEYINPUT83), .B(KEYINPUT32), .Z(n355) );
  XNOR2_X1 U499 ( .A(n477), .B(n382), .ZN(n624) );
  INV_X1 U500 ( .A(KEYINPUT44), .ZN(n550) );
  AND2_X1 U501 ( .A1(n568), .A2(n398), .ZN(n422) );
  NAND2_X1 U502 ( .A1(n363), .A2(n598), .ZN(n599) );
  INV_X1 U503 ( .A(n653), .ZN(n397) );
  INV_X1 U504 ( .A(n571), .ZN(n399) );
  NAND2_X1 U505 ( .A1(n416), .A2(n356), .ZN(n358) );
  AND2_X1 U506 ( .A1(n359), .A2(n557), .ZN(n616) );
  NAND2_X1 U507 ( .A1(n359), .A2(n723), .ZN(n724) );
  XNOR2_X2 U508 ( .A(n408), .B(KEYINPUT45), .ZN(n359) );
  NAND2_X1 U509 ( .A1(n747), .A2(n639), .ZN(n418) );
  NAND2_X1 U510 ( .A1(n437), .A2(n362), .ZN(n404) );
  NAND2_X1 U511 ( .A1(n715), .A2(G472), .ZN(n626) );
  AND2_X4 U512 ( .A1(n430), .A2(n623), .ZN(n715) );
  NAND2_X1 U513 ( .A1(n597), .A2(n417), .ZN(n363) );
  NOR2_X1 U514 ( .A1(n608), .A2(n576), .ZN(n577) );
  NAND2_X1 U515 ( .A1(n571), .A2(n580), .ZN(n365) );
  XNOR2_X1 U516 ( .A(n385), .B(KEYINPUT92), .ZN(n491) );
  XNOR2_X1 U517 ( .A(n609), .B(n610), .ZN(n746) );
  NOR2_X1 U518 ( .A1(n675), .A2(n369), .ZN(n676) );
  AND2_X2 U519 ( .A1(n370), .A2(n622), .ZN(n623) );
  NAND2_X1 U520 ( .A1(n430), .A2(n370), .ZN(n690) );
  NAND2_X1 U521 ( .A1(n373), .A2(n371), .ZN(n406) );
  INV_X1 U522 ( .A(n649), .ZN(n372) );
  AND2_X1 U523 ( .A1(n378), .A2(n374), .ZN(n373) );
  NAND2_X1 U524 ( .A1(n649), .A2(n352), .ZN(n378) );
  NAND2_X1 U525 ( .A1(n379), .A2(n738), .ZN(n739) );
  XNOR2_X1 U526 ( .A(n380), .B(n748), .ZN(G33) );
  NAND2_X1 U527 ( .A1(n441), .A2(n384), .ZN(n602) );
  AND2_X1 U528 ( .A1(n354), .A2(n582), .ZN(n384) );
  INV_X1 U529 ( .A(n548), .ZN(n387) );
  NAND2_X1 U530 ( .A1(n548), .A2(n355), .ZN(n389) );
  XNOR2_X2 U531 ( .A(n545), .B(KEYINPUT22), .ZN(n548) );
  NOR2_X1 U532 ( .A1(n423), .A2(n399), .ZN(n398) );
  XNOR2_X1 U533 ( .A(n590), .B(n589), .ZN(n592) );
  NOR2_X1 U534 ( .A1(n717), .A2(G902), .ZN(n474) );
  AND2_X1 U535 ( .A1(n396), .A2(n593), .ZN(n598) );
  NOR2_X1 U536 ( .A1(n397), .A2(n594), .ZN(n396) );
  NOR2_X2 U537 ( .A1(n709), .A2(n719), .ZN(n711) );
  XNOR2_X2 U538 ( .A(n572), .B(n401), .ZN(n591) );
  XNOR2_X2 U539 ( .A(n455), .B(G469), .ZN(n572) );
  XNOR2_X1 U540 ( .A(n402), .B(n630), .ZN(G57) );
  NOR2_X2 U541 ( .A1(n627), .A2(n719), .ZN(n402) );
  XNOR2_X1 U542 ( .A(n403), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U543 ( .A1(n698), .A2(n719), .ZN(n403) );
  AND2_X1 U544 ( .A1(n415), .A2(n409), .ZN(n407) );
  NAND2_X1 U545 ( .A1(n418), .A2(KEYINPUT44), .ZN(n409) );
  AND2_X1 U546 ( .A1(n544), .A2(n410), .ZN(n555) );
  INV_X1 U547 ( .A(n544), .ZN(n411) );
  OR2_X1 U548 ( .A1(n548), .A2(n413), .ZN(n631) );
  NAND2_X1 U549 ( .A1(n745), .A2(KEYINPUT44), .ZN(n415) );
  INV_X1 U550 ( .A(n745), .ZN(n416) );
  XNOR2_X2 U551 ( .A(n541), .B(KEYINPUT35), .ZN(n745) );
  INV_X1 U552 ( .A(n591), .ZN(n655) );
  NAND2_X1 U553 ( .A1(n554), .A2(n568), .ZN(n484) );
  NAND2_X1 U554 ( .A1(n421), .A2(n591), .ZN(n420) );
  INV_X1 U555 ( .A(n656), .ZN(n421) );
  NAND2_X1 U556 ( .A1(n569), .A2(n429), .ZN(n428) );
  NAND2_X1 U557 ( .A1(n435), .A2(n437), .ZN(n431) );
  AND2_X1 U558 ( .A1(n612), .A2(n440), .ZN(n439) );
  XNOR2_X1 U559 ( .A(n442), .B(n581), .ZN(n441) );
  NAND2_X1 U560 ( .A1(n580), .A2(n671), .ZN(n442) );
  XNOR2_X1 U561 ( .A(n546), .B(n443), .ZN(n580) );
  INV_X1 U562 ( .A(KEYINPUT107), .ZN(n443) );
  INV_X1 U563 ( .A(n659), .ZN(n542) );
  XNOR2_X1 U564 ( .A(KEYINPUT46), .B(KEYINPUT88), .ZN(n611) );
  XNOR2_X1 U565 ( .A(n475), .B(KEYINPUT97), .ZN(n476) );
  XNOR2_X1 U566 ( .A(n731), .B(G146), .ZN(n450) );
  XNOR2_X1 U567 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U568 ( .A(n510), .B(KEYINPUT74), .ZN(n511) );
  INV_X1 U569 ( .A(n601), .ZN(n583) );
  XNOR2_X1 U570 ( .A(n498), .B(n497), .ZN(n720) );
  XNOR2_X1 U571 ( .A(n708), .B(n707), .ZN(n709) );
  XNOR2_X1 U572 ( .A(n629), .B(n628), .ZN(n630) );
  INV_X1 U573 ( .A(n561), .ZN(n741) );
  XNOR2_X2 U574 ( .A(KEYINPUT65), .B(KEYINPUT70), .ZN(n445) );
  XOR2_X1 U575 ( .A(G101), .B(KEYINPUT68), .Z(n447) );
  XNOR2_X1 U576 ( .A(KEYINPUT67), .B(n447), .ZN(n448) );
  XNOR2_X1 U577 ( .A(n449), .B(G134), .ZN(n731) );
  XOR2_X1 U578 ( .A(G104), .B(G110), .Z(n451) );
  XOR2_X1 U579 ( .A(G107), .B(n451), .Z(n496) );
  XOR2_X1 U580 ( .A(n460), .B(n496), .Z(n453) );
  NAND2_X1 U581 ( .A1(G227), .A2(n741), .ZN(n452) );
  XNOR2_X1 U582 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U583 ( .A(n477), .B(n454), .ZN(n699) );
  XNOR2_X1 U584 ( .A(G902), .B(KEYINPUT15), .ZN(n485) );
  NAND2_X1 U585 ( .A1(G234), .A2(n485), .ZN(n456) );
  XNOR2_X1 U586 ( .A(KEYINPUT20), .B(n456), .ZN(n470) );
  NAND2_X1 U587 ( .A1(n470), .A2(G221), .ZN(n457) );
  XNOR2_X1 U588 ( .A(KEYINPUT21), .B(n457), .ZN(n659) );
  NAND2_X1 U589 ( .A1(n741), .A2(G234), .ZN(n458) );
  XOR2_X1 U590 ( .A(KEYINPUT8), .B(n458), .Z(n534) );
  NAND2_X1 U591 ( .A1(n534), .A2(G221), .ZN(n469) );
  XNOR2_X1 U592 ( .A(KEYINPUT10), .B(KEYINPUT71), .ZN(n459) );
  XOR2_X1 U593 ( .A(KEYINPUT23), .B(G110), .Z(n462) );
  XNOR2_X1 U594 ( .A(n462), .B(n461), .ZN(n466) );
  XOR2_X1 U595 ( .A(KEYINPUT24), .B(KEYINPUT95), .Z(n464) );
  XNOR2_X1 U596 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U597 ( .A(n733), .B(n467), .ZN(n468) );
  XNOR2_X1 U598 ( .A(n468), .B(n469), .ZN(n717) );
  NAND2_X1 U599 ( .A1(G217), .A2(n470), .ZN(n472) );
  XOR2_X1 U600 ( .A(KEYINPUT80), .B(KEYINPUT25), .Z(n471) );
  XNOR2_X2 U601 ( .A(n474), .B(n473), .ZN(n658) );
  XOR2_X1 U602 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n475) );
  XNOR2_X1 U603 ( .A(G116), .B(G113), .ZN(n478) );
  XNOR2_X1 U604 ( .A(n351), .B(n478), .ZN(n479) );
  NOR2_X1 U605 ( .A1(G953), .A2(G237), .ZN(n480) );
  XOR2_X1 U606 ( .A(KEYINPUT79), .B(n480), .Z(n517) );
  NAND2_X1 U607 ( .A1(n517), .A2(G210), .ZN(n481) );
  INV_X1 U608 ( .A(KEYINPUT33), .ZN(n483) );
  INV_X1 U609 ( .A(n485), .ZN(n622) );
  NAND2_X1 U610 ( .A1(G224), .A2(n741), .ZN(n486) );
  XNOR2_X1 U611 ( .A(n487), .B(n486), .ZN(n489) );
  XNOR2_X1 U612 ( .A(n488), .B(n489), .ZN(n490) );
  XNOR2_X1 U613 ( .A(n491), .B(n490), .ZN(n499) );
  XNOR2_X1 U614 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U615 ( .A(n495), .B(n494), .ZN(n498) );
  INV_X1 U616 ( .A(n496), .ZN(n497) );
  XNOR2_X1 U617 ( .A(n499), .B(n720), .ZN(n695) );
  NOR2_X1 U618 ( .A1(n622), .A2(n695), .ZN(n501) );
  OR2_X1 U619 ( .A1(G237), .A2(G902), .ZN(n502) );
  NAND2_X1 U620 ( .A1(G210), .A2(n502), .ZN(n500) );
  XNOR2_X1 U621 ( .A(n501), .B(n500), .ZN(n558) );
  NAND2_X1 U622 ( .A1(G214), .A2(n502), .ZN(n671) );
  NAND2_X1 U623 ( .A1(n558), .A2(n671), .ZN(n588) );
  NAND2_X1 U624 ( .A1(G234), .A2(G237), .ZN(n503) );
  XNOR2_X1 U625 ( .A(n503), .B(KEYINPUT14), .ZN(n505) );
  NAND2_X1 U626 ( .A1(n505), .A2(G902), .ZN(n504) );
  XOR2_X1 U627 ( .A(n504), .B(KEYINPUT94), .Z(n559) );
  NOR2_X1 U628 ( .A1(G898), .A2(n723), .ZN(n722) );
  NAND2_X1 U629 ( .A1(n559), .A2(n722), .ZN(n507) );
  NAND2_X1 U630 ( .A1(G952), .A2(n505), .ZN(n685) );
  NOR2_X1 U631 ( .A1(n685), .A2(G953), .ZN(n506) );
  XNOR2_X1 U632 ( .A(n506), .B(KEYINPUT93), .ZN(n564) );
  NAND2_X1 U633 ( .A1(n507), .A2(n564), .ZN(n508) );
  XNOR2_X1 U634 ( .A(KEYINPUT34), .B(KEYINPUT82), .ZN(n510) );
  XNOR2_X1 U635 ( .A(n512), .B(n511), .ZN(n540) );
  XOR2_X1 U636 ( .A(G122), .B(G104), .Z(n514) );
  XNOR2_X1 U637 ( .A(G113), .B(G131), .ZN(n513) );
  XNOR2_X1 U638 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U639 ( .A(n516), .B(n515), .ZN(n519) );
  NAND2_X1 U640 ( .A1(G214), .A2(n517), .ZN(n518) );
  XNOR2_X1 U641 ( .A(n519), .B(n518), .ZN(n527) );
  XNOR2_X1 U642 ( .A(n521), .B(n520), .ZN(n525) );
  XNOR2_X1 U643 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U644 ( .A(n525), .B(n524), .Z(n526) );
  XNOR2_X1 U645 ( .A(KEYINPUT13), .B(KEYINPUT103), .ZN(n528) );
  XNOR2_X1 U646 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n537) );
  XNOR2_X1 U647 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U648 ( .A(n533), .B(n532), .Z(n536) );
  NAND2_X1 U649 ( .A1(G217), .A2(n534), .ZN(n535) );
  NOR2_X1 U650 ( .A1(G902), .A2(n713), .ZN(n538) );
  NAND2_X1 U651 ( .A1(n551), .A2(n552), .ZN(n586) );
  INV_X1 U652 ( .A(n586), .ZN(n539) );
  NAND2_X1 U653 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U654 ( .A1(n551), .A2(n552), .ZN(n607) );
  NAND2_X1 U655 ( .A1(n544), .A2(n543), .ZN(n545) );
  INV_X1 U656 ( .A(n658), .ZN(n567) );
  OR2_X1 U657 ( .A1(n567), .A2(n580), .ZN(n547) );
  NOR2_X1 U658 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U659 ( .A1(n655), .A2(n549), .ZN(n639) );
  XOR2_X1 U660 ( .A(KEYINPUT104), .B(n551), .Z(n553) );
  NAND2_X1 U661 ( .A1(n553), .A2(n552), .ZN(n650) );
  INV_X1 U662 ( .A(n650), .ZN(n640) );
  NOR2_X1 U663 ( .A1(n644), .A2(n640), .ZN(n675) );
  NAND2_X1 U664 ( .A1(n663), .A2(n554), .ZN(n668) );
  NAND2_X1 U665 ( .A1(n354), .A2(n555), .ZN(n634) );
  NOR2_X1 U666 ( .A1(n591), .A2(n658), .ZN(n556) );
  INV_X1 U667 ( .A(KEYINPUT85), .ZN(n557) );
  INV_X1 U668 ( .A(n559), .ZN(n560) );
  NOR2_X1 U669 ( .A1(n560), .A2(G900), .ZN(n562) );
  NAND2_X1 U670 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U671 ( .A(n563), .B(KEYINPUT108), .ZN(n565) );
  NAND2_X1 U672 ( .A1(n565), .A2(n564), .ZN(n582) );
  NAND2_X1 U673 ( .A1(n542), .A2(n582), .ZN(n566) );
  NOR2_X1 U674 ( .A1(n567), .A2(n566), .ZN(n571) );
  INV_X1 U675 ( .A(n587), .ZN(n569) );
  NAND2_X1 U676 ( .A1(n675), .A2(KEYINPUT86), .ZN(n578) );
  INV_X1 U677 ( .A(n570), .ZN(n576) );
  XNOR2_X1 U678 ( .A(n572), .B(KEYINPUT111), .ZN(n573) );
  NAND2_X1 U679 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U680 ( .A(n577), .B(KEYINPUT84), .ZN(n645) );
  NAND2_X1 U681 ( .A1(n578), .A2(n645), .ZN(n579) );
  AND2_X1 U682 ( .A1(n579), .A2(KEYINPUT47), .ZN(n600) );
  INV_X1 U683 ( .A(KEYINPUT30), .ZN(n581) );
  NOR2_X1 U684 ( .A1(n583), .A2(n602), .ZN(n584) );
  XOR2_X1 U685 ( .A(KEYINPUT110), .B(n584), .Z(n585) );
  XNOR2_X1 U686 ( .A(n643), .B(KEYINPUT87), .ZN(n593) );
  NOR2_X1 U687 ( .A1(n588), .A2(n587), .ZN(n590) );
  NAND2_X1 U688 ( .A1(n592), .A2(n591), .ZN(n653) );
  NOR2_X1 U689 ( .A1(KEYINPUT86), .A2(KEYINPUT47), .ZN(n594) );
  INV_X1 U690 ( .A(KEYINPUT47), .ZN(n595) );
  NAND2_X1 U691 ( .A1(n595), .A2(n645), .ZN(n596) );
  NAND2_X1 U692 ( .A1(n596), .A2(KEYINPUT86), .ZN(n597) );
  INV_X1 U693 ( .A(n672), .ZN(n603) );
  XNOR2_X1 U694 ( .A(KEYINPUT89), .B(KEYINPUT39), .ZN(n604) );
  NAND2_X1 U695 ( .A1(n614), .A2(n644), .ZN(n606) );
  XNOR2_X1 U696 ( .A(KEYINPUT114), .B(KEYINPUT42), .ZN(n610) );
  INV_X1 U697 ( .A(n607), .ZN(n674) );
  NAND2_X1 U698 ( .A1(n614), .A2(n640), .ZN(n738) );
  NAND2_X1 U699 ( .A1(n616), .A2(n615), .ZN(n617) );
  INV_X1 U700 ( .A(KEYINPUT2), .ZN(n618) );
  XOR2_X1 U701 ( .A(n738), .B(KEYINPUT85), .Z(n619) );
  AND2_X1 U702 ( .A1(n619), .A2(KEYINPUT2), .ZN(n620) );
  XNOR2_X1 U703 ( .A(n624), .B(KEYINPUT62), .ZN(n625) );
  XNOR2_X1 U704 ( .A(n626), .B(n625), .ZN(n627) );
  XNOR2_X1 U705 ( .A(KEYINPUT115), .B(KEYINPUT63), .ZN(n629) );
  INV_X1 U706 ( .A(KEYINPUT91), .ZN(n628) );
  XNOR2_X1 U707 ( .A(G101), .B(n631), .ZN(G3) );
  NOR2_X1 U708 ( .A1(n423), .A2(n634), .ZN(n632) );
  XOR2_X1 U709 ( .A(KEYINPUT116), .B(n632), .Z(n633) );
  XNOR2_X1 U710 ( .A(G104), .B(n633), .ZN(G6) );
  NOR2_X1 U711 ( .A1(n650), .A2(n634), .ZN(n636) );
  XNOR2_X1 U712 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n635) );
  XNOR2_X1 U713 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U714 ( .A(G107), .B(n637), .ZN(G9) );
  XOR2_X1 U715 ( .A(G110), .B(KEYINPUT117), .Z(n638) );
  XNOR2_X1 U716 ( .A(n639), .B(n638), .ZN(G12) );
  XOR2_X1 U717 ( .A(G128), .B(KEYINPUT29), .Z(n642) );
  NAND2_X1 U718 ( .A1(n640), .A2(n645), .ZN(n641) );
  XNOR2_X1 U719 ( .A(n642), .B(n641), .ZN(G30) );
  XOR2_X1 U720 ( .A(G143), .B(n643), .Z(G45) );
  NAND2_X1 U721 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U722 ( .A(n646), .B(G146), .ZN(G48) );
  NOR2_X1 U723 ( .A1(n423), .A2(n649), .ZN(n647) );
  XOR2_X1 U724 ( .A(KEYINPUT118), .B(n647), .Z(n648) );
  XNOR2_X1 U725 ( .A(G113), .B(n648), .ZN(G15) );
  NOR2_X1 U726 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U727 ( .A(G116), .B(n651), .Z(G18) );
  XOR2_X1 U728 ( .A(G125), .B(KEYINPUT37), .Z(n652) );
  XNOR2_X1 U729 ( .A(n653), .B(n652), .ZN(G27) );
  XNOR2_X1 U730 ( .A(G134), .B(n738), .ZN(G36) );
  XOR2_X1 U731 ( .A(G140), .B(n654), .Z(G42) );
  AND2_X1 U732 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U733 ( .A(KEYINPUT50), .B(n657), .Z(n666) );
  XOR2_X1 U734 ( .A(KEYINPUT119), .B(KEYINPUT49), .Z(n661) );
  NAND2_X1 U735 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U736 ( .A(n661), .B(n660), .ZN(n662) );
  NOR2_X1 U737 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U738 ( .A(KEYINPUT120), .B(n664), .ZN(n665) );
  NAND2_X1 U739 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U740 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U741 ( .A(KEYINPUT51), .B(n669), .ZN(n670) );
  NOR2_X1 U742 ( .A1(n686), .A2(n670), .ZN(n681) );
  NOR2_X1 U743 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U744 ( .A1(n674), .A2(n673), .ZN(n677) );
  NOR2_X1 U745 ( .A1(n677), .A2(n676), .ZN(n679) );
  NOR2_X1 U746 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U747 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U748 ( .A(n682), .B(KEYINPUT52), .Z(n683) );
  XNOR2_X1 U749 ( .A(KEYINPUT121), .B(n683), .ZN(n684) );
  NOR2_X1 U750 ( .A1(n685), .A2(n684), .ZN(n689) );
  OR2_X1 U751 ( .A1(n686), .A2(n678), .ZN(n687) );
  XOR2_X1 U752 ( .A(KEYINPUT122), .B(n687), .Z(n688) );
  NOR2_X1 U753 ( .A1(n689), .A2(n688), .ZN(n691) );
  NAND2_X1 U754 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U755 ( .A1(n692), .A2(G953), .ZN(n693) );
  XNOR2_X1 U756 ( .A(n693), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U757 ( .A1(n715), .A2(G210), .ZN(n697) );
  XOR2_X1 U758 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n694) );
  XNOR2_X1 U759 ( .A(n697), .B(n696), .ZN(n698) );
  XNOR2_X1 U760 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n701) );
  XNOR2_X1 U761 ( .A(n699), .B(KEYINPUT57), .ZN(n700) );
  XNOR2_X1 U762 ( .A(n701), .B(n700), .ZN(n703) );
  NAND2_X1 U763 ( .A1(n715), .A2(G469), .ZN(n702) );
  XNOR2_X1 U764 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U765 ( .A1(n719), .A2(n704), .ZN(G54) );
  NAND2_X1 U766 ( .A1(n715), .A2(G475), .ZN(n708) );
  XOR2_X1 U767 ( .A(KEYINPUT59), .B(KEYINPUT124), .Z(n705) );
  XNOR2_X1 U768 ( .A(KEYINPUT66), .B(KEYINPUT60), .ZN(n710) );
  XNOR2_X1 U769 ( .A(n711), .B(n710), .ZN(G60) );
  NAND2_X1 U770 ( .A1(G478), .A2(n715), .ZN(n712) );
  XNOR2_X1 U771 ( .A(n713), .B(n712), .ZN(n714) );
  NOR2_X1 U772 ( .A1(n719), .A2(n714), .ZN(G63) );
  NAND2_X1 U773 ( .A1(G217), .A2(n715), .ZN(n716) );
  XNOR2_X1 U774 ( .A(n717), .B(n716), .ZN(n718) );
  NOR2_X1 U775 ( .A1(n719), .A2(n718), .ZN(G66) );
  XNOR2_X1 U776 ( .A(G101), .B(n720), .ZN(n721) );
  NOR2_X1 U777 ( .A1(n722), .A2(n721), .ZN(n730) );
  XOR2_X1 U778 ( .A(KEYINPUT125), .B(n724), .Z(n728) );
  NAND2_X1 U779 ( .A1(G953), .A2(G224), .ZN(n725) );
  XNOR2_X1 U780 ( .A(KEYINPUT61), .B(n725), .ZN(n726) );
  NAND2_X1 U781 ( .A1(n726), .A2(G898), .ZN(n727) );
  NAND2_X1 U782 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U783 ( .A(n730), .B(n729), .ZN(G69) );
  XNOR2_X1 U784 ( .A(n732), .B(n731), .ZN(n734) );
  XNOR2_X1 U785 ( .A(n733), .B(n734), .ZN(n740) );
  XNOR2_X1 U786 ( .A(G227), .B(n740), .ZN(n735) );
  NAND2_X1 U787 ( .A1(n735), .A2(G900), .ZN(n736) );
  XNOR2_X1 U788 ( .A(KEYINPUT126), .B(n736), .ZN(n737) );
  NAND2_X1 U789 ( .A1(n737), .A2(G953), .ZN(n744) );
  XNOR2_X1 U790 ( .A(n740), .B(n739), .ZN(n742) );
  NAND2_X1 U791 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U792 ( .A1(n744), .A2(n743), .ZN(G72) );
  XOR2_X1 U793 ( .A(n745), .B(G122), .Z(G24) );
  XOR2_X1 U794 ( .A(n746), .B(G137), .Z(G39) );
  XNOR2_X1 U795 ( .A(n747), .B(G119), .ZN(G21) );
  XNOR2_X1 U796 ( .A(G131), .B(KEYINPUT127), .ZN(n748) );
endmodule

