//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 1 1 0 0 0 0 1 1 0 0 0 0 0 0 0 0 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n623, new_n624, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190,
    new_n1191;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT65), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  INV_X1    g031(.A(G2105), .ZN(new_n457));
  INV_X1    g032(.A(G2104), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  AND3_X1   g036(.A1(new_n459), .A2(new_n461), .A3(KEYINPUT66), .ZN(new_n462));
  AOI21_X1  g037(.A(KEYINPUT66), .B1(new_n459), .B2(new_n461), .ZN(new_n463));
  OAI21_X1  g038(.A(G125), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n457), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n459), .A2(new_n461), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G137), .ZN(new_n468));
  NAND2_X1  g043(.A1(G101), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n466), .A2(new_n470), .ZN(G160));
  NAND2_X1  g046(.A1(new_n459), .A2(new_n461), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(new_n457), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G124), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n472), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G136), .ZN(new_n476));
  OR2_X1    g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n477), .B(G2104), .C1(G112), .C2(new_n457), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n474), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  INV_X1    g055(.A(G138), .ZN(new_n481));
  NOR3_X1   g056(.A1(new_n481), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n482), .B1(new_n462), .B2(new_n463), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n467), .A2(new_n457), .ZN(new_n486));
  OAI21_X1  g061(.A(KEYINPUT4), .B1(new_n486), .B2(new_n481), .ZN(new_n487));
  OAI211_X1 g062(.A(KEYINPUT69), .B(new_n482), .C1(new_n462), .C2(new_n463), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n485), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AND2_X1   g064(.A1(KEYINPUT67), .A2(G114), .ZN(new_n490));
  NOR2_X1   g065(.A1(KEYINPUT67), .A2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(G2105), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  OAI211_X1 g070(.A(KEYINPUT68), .B(G2105), .C1(new_n490), .C2(new_n491), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n494), .A2(G2104), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n473), .A2(G126), .ZN(new_n498));
  AND2_X1   g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n489), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  NAND2_X1  g076(.A1(G62), .A2(G651), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT70), .B1(new_n503), .B2(G651), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT6), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n503), .A2(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n502), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(G75), .A2(G651), .ZN(new_n520));
  INV_X1    g095(.A(G50), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n520), .B1(new_n510), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT71), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT71), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n519), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(new_n527), .ZN(G166));
  AOI22_X1  g103(.A1(new_n504), .A2(new_n507), .B1(new_n503), .B2(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(new_n518), .ZN(new_n530));
  INV_X1    g105(.A(G89), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n530), .B1(KEYINPUT72), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n532), .B1(KEYINPUT72), .B2(new_n531), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n510), .A2(new_n513), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G51), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n533), .A2(new_n535), .A3(new_n537), .A4(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  AOI22_X1  g115(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n541), .A2(new_n506), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n510), .A2(new_n517), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G90), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n536), .A2(G52), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n542), .A2(new_n544), .A3(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G56), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n517), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n536), .A2(G43), .B1(G651), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n543), .A2(G81), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT74), .ZN(new_n559));
  XOR2_X1   g134(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n560));
  XNOR2_X1  g135(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n556), .A2(new_n561), .ZN(G188));
  NAND3_X1  g137(.A1(new_n529), .A2(G91), .A3(new_n518), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT76), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT76), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n529), .A2(new_n565), .A3(new_n518), .A4(G91), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT77), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n514), .A2(new_n516), .A3(G65), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n567), .B1(new_n570), .B2(G651), .ZN(new_n571));
  AOI211_X1 g146(.A(KEYINPUT77), .B(new_n506), .C1(new_n568), .C2(new_n569), .ZN(new_n572));
  OAI211_X1 g147(.A(new_n564), .B(new_n566), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  XOR2_X1   g148(.A(KEYINPUT75), .B(KEYINPUT9), .Z(new_n574));
  NAND4_X1  g149(.A1(new_n529), .A2(G53), .A3(G543), .A4(new_n574), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n529), .A2(G53), .A3(G543), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT9), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(KEYINPUT75), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n573), .B1(new_n575), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G299));
  INV_X1    g156(.A(G166), .ZN(G303));
  NAND3_X1  g157(.A1(new_n529), .A2(G49), .A3(G543), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n529), .A2(G87), .A3(new_n518), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G288));
  AOI22_X1  g161(.A1(new_n529), .A2(G48), .B1(G73), .B2(G651), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(new_n513), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n529), .A2(G86), .B1(G61), .B2(G651), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(new_n517), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G305));
  NAND2_X1  g167(.A1(G72), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G60), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n517), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n536), .A2(G47), .B1(G651), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n543), .A2(G85), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT78), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n543), .A2(new_n600), .A3(G92), .ZN(new_n601));
  INV_X1    g176(.A(G92), .ZN(new_n602));
  OAI21_X1  g177(.A(KEYINPUT78), .B1(new_n530), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g178(.A(KEYINPUT10), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n518), .A2(G66), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT80), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n506), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n601), .A2(KEYINPUT10), .A3(new_n603), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n529), .A2(G543), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n612), .A2(KEYINPUT79), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(KEYINPUT79), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n613), .A2(G54), .A3(new_n614), .ZN(new_n615));
  NAND4_X1  g190(.A1(new_n605), .A2(new_n610), .A3(new_n611), .A4(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT81), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n599), .B1(new_n617), .B2(G868), .ZN(G284));
  OAI21_X1  g193(.A(new_n599), .B1(new_n617), .B2(G868), .ZN(G321));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G868), .B2(new_n580), .ZN(G297));
  OAI21_X1  g196(.A(new_n620), .B1(G868), .B2(new_n580), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n617), .B1(new_n623), .B2(G860), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT82), .ZN(G148));
  NAND2_X1  g200(.A1(new_n617), .A2(new_n623), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g204(.A1(new_n462), .A2(new_n463), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n458), .A2(G2105), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(KEYINPUT12), .ZN(new_n633));
  INV_X1    g208(.A(KEYINPUT12), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n630), .A2(new_n634), .A3(new_n631), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT83), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n638), .A2(G2100), .ZN(new_n639));
  AND2_X1   g214(.A1(new_n638), .A2(G2100), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n473), .A2(G123), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n475), .A2(G135), .ZN(new_n643));
  NOR2_X1   g218(.A1(G99), .A2(G2105), .ZN(new_n644));
  OAI21_X1  g219(.A(G2104), .B1(new_n457), .B2(G111), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n642), .B(new_n643), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(G2096), .Z(new_n647));
  OAI211_X1 g222(.A(new_n641), .B(new_n647), .C1(new_n637), .C2(new_n639), .ZN(G156));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XOR2_X1   g225(.A(G2443), .B(G2446), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2427), .B(G2438), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2430), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT15), .B(G2435), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT14), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n654), .B(new_n659), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n660), .A2(G14), .ZN(G401));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT17), .ZN(new_n663));
  XOR2_X1   g238(.A(G2067), .B(G2678), .Z(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  NAND3_X1  g240(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT84), .Z(new_n667));
  INV_X1    g242(.A(new_n665), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n664), .A2(new_n662), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n668), .B(new_n669), .C1(new_n663), .C2(new_n664), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n668), .A2(new_n664), .A3(new_n662), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT18), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n667), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2096), .B(G2100), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT85), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g261(.A(KEYINPUT85), .B1(new_n678), .B2(new_n680), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n683), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT20), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n677), .A2(new_n679), .ZN(new_n691));
  OR3_X1    g266(.A1(new_n686), .A2(new_n681), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n688), .A2(new_n689), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n686), .A2(new_n691), .ZN(new_n694));
  NAND4_X1  g269(.A1(new_n690), .A2(new_n692), .A3(new_n693), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(G1991), .B(G1996), .Z(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT86), .B(KEYINPUT87), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n697), .B(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(G229));
  NAND2_X1  g279(.A1(new_n473), .A2(G128), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n475), .A2(G140), .ZN(new_n706));
  NOR2_X1   g281(.A1(G104), .A2(G2105), .ZN(new_n707));
  OAI21_X1  g282(.A(G2104), .B1(new_n457), .B2(G116), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n705), .B(new_n706), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT93), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n712), .A2(G26), .ZN(new_n714));
  OAI21_X1  g289(.A(KEYINPUT28), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(KEYINPUT28), .B2(new_n714), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(G2067), .ZN(new_n717));
  AOI22_X1  g292(.A1(G129), .A2(new_n473), .B1(new_n475), .B2(G141), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n631), .A2(G105), .ZN(new_n719));
  NAND3_X1  g294(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT26), .Z(new_n721));
  NAND3_X1  g296(.A1(new_n718), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n722), .A2(KEYINPUT96), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(KEYINPUT96), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G29), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G29), .B2(G32), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT27), .B(G1996), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT24), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n712), .B1(new_n729), .B2(G34), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT95), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n729), .B2(G34), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G160), .B2(G29), .ZN(new_n736));
  OAI22_X1  g311(.A1(new_n727), .A2(new_n728), .B1(G2084), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(G171), .A2(G16), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G5), .B2(G16), .ZN(new_n739));
  INV_X1    g314(.A(G1961), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR3_X1   g316(.A1(new_n717), .A2(new_n737), .A3(new_n741), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT30), .B(G28), .Z(new_n743));
  MUX2_X1   g318(.A(new_n743), .B(new_n646), .S(G29), .Z(new_n744));
  INV_X1    g319(.A(G16), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n554), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n745), .B2(G19), .ZN(new_n747));
  INV_X1    g322(.A(G1341), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n712), .A2(G35), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G162), .B2(new_n712), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT29), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G2090), .ZN(new_n752));
  OAI221_X1 g327(.A(new_n744), .B1(new_n747), .B2(new_n748), .C1(new_n752), .C2(KEYINPUT98), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n727), .A2(new_n728), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n747), .A2(new_n748), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n739), .A2(new_n740), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  AOI211_X1 g332(.A(new_n753), .B(new_n757), .C1(G2084), .C2(new_n736), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n751), .A2(G2090), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT31), .B(G11), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n742), .A2(new_n758), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(KEYINPUT97), .B1(G16), .B2(G21), .ZN(new_n762));
  NOR2_X1   g337(.A1(G286), .A2(new_n745), .ZN(new_n763));
  MUX2_X1   g338(.A(new_n762), .B(KEYINPUT97), .S(new_n763), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G1966), .ZN(new_n765));
  NOR2_X1   g340(.A1(G164), .A2(new_n712), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G27), .B2(new_n712), .ZN(new_n767));
  INV_X1    g342(.A(G2078), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n631), .A2(G103), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT25), .ZN(new_n772));
  INV_X1    g347(.A(G139), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(new_n486), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT94), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n630), .A2(G127), .ZN(new_n776));
  NAND2_X1  g351(.A1(G115), .A2(G2104), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n457), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  MUX2_X1   g355(.A(G33), .B(new_n780), .S(G29), .Z(new_n781));
  AOI22_X1  g356(.A1(new_n781), .A2(G2072), .B1(KEYINPUT98), .B2(new_n752), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n765), .A2(new_n769), .A3(new_n770), .A4(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n781), .A2(G2072), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n745), .A2(G20), .ZN(new_n785));
  OAI211_X1 g360(.A(KEYINPUT23), .B(new_n785), .C1(new_n580), .C2(new_n745), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(KEYINPUT23), .B2(new_n785), .ZN(new_n787));
  INV_X1    g362(.A(G1956), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NOR4_X1   g364(.A1(new_n761), .A2(new_n783), .A3(new_n784), .A4(new_n789), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n745), .A2(G24), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G290), .B2(G16), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT88), .B(G1986), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT89), .ZN(new_n794));
  AOI21_X1  g369(.A(KEYINPUT91), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n794), .B2(new_n792), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n745), .A2(G23), .ZN(new_n797));
  INV_X1    g372(.A(G288), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(new_n745), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT33), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1976), .ZN(new_n801));
  NOR2_X1   g376(.A1(G16), .A2(G22), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G166), .B2(G16), .ZN(new_n803));
  INV_X1    g378(.A(G1971), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n745), .A2(G6), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n591), .B2(new_n745), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT32), .B(G1981), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n801), .A2(new_n805), .A3(new_n809), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT90), .B(KEYINPUT34), .Z(new_n811));
  AOI21_X1  g386(.A(new_n796), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n712), .A2(G25), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n473), .A2(G119), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n475), .A2(G131), .ZN(new_n815));
  OR2_X1    g390(.A1(G95), .A2(G2105), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n816), .B(G2104), .C1(G107), .C2(new_n457), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n814), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n813), .B1(new_n819), .B2(new_n712), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT35), .B(G1991), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n812), .B(new_n822), .C1(new_n811), .C2(new_n810), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT36), .ZN(new_n824));
  NOR2_X1   g399(.A1(G4), .A2(G16), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(new_n617), .B2(G16), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT92), .B(G1348), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  AND3_X1   g403(.A1(new_n790), .A2(new_n824), .A3(new_n828), .ZN(G311));
  NAND3_X1  g404(.A1(new_n790), .A2(new_n824), .A3(new_n828), .ZN(G150));
  NAND2_X1  g405(.A1(new_n543), .A2(G93), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT100), .B(G55), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n536), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(G80), .A2(G543), .ZN(new_n834));
  INV_X1    g409(.A(G67), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n517), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(G651), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n831), .A2(new_n833), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(G860), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT37), .Z(new_n840));
  NAND2_X1  g415(.A1(new_n617), .A2(G559), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT39), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n838), .B1(new_n552), .B2(new_n551), .ZN(new_n843));
  AND3_X1   g418(.A1(new_n831), .A2(new_n833), .A3(new_n837), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n844), .A2(new_n553), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n842), .B(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n840), .B1(new_n849), .B2(G860), .ZN(G145));
  XOR2_X1   g425(.A(G160), .B(new_n646), .Z(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT102), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n780), .A2(new_n725), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n775), .B(new_n779), .C1(new_n723), .C2(new_n724), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n710), .A2(G164), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n711), .A2(new_n500), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n858), .A2(new_n857), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n860), .A2(new_n854), .A3(new_n855), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n636), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n473), .A2(G130), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n475), .A2(G142), .ZN(new_n865));
  NOR2_X1   g440(.A1(G106), .A2(G2105), .ZN(new_n866));
  OAI21_X1  g441(.A(G2104), .B1(new_n457), .B2(G118), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n864), .B(new_n865), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  AND2_X1   g443(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n863), .A2(new_n868), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n818), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n636), .B(new_n868), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(new_n819), .ZN(new_n873));
  AOI21_X1  g448(.A(KEYINPUT101), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n853), .B1(new_n862), .B2(new_n875), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n871), .A2(new_n873), .A3(KEYINPUT101), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n859), .B(new_n861), .C1(new_n877), .C2(new_n874), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n876), .A2(new_n479), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n479), .B1(new_n876), .B2(new_n878), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n852), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(G37), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n862), .A2(new_n875), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n883), .A2(new_n878), .A3(KEYINPUT102), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(G162), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n876), .A2(new_n479), .A3(new_n878), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(new_n851), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n881), .A2(new_n882), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g464(.A(G868), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n838), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n626), .B(new_n846), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n611), .A2(new_n615), .ZN(new_n893));
  NOR3_X1   g468(.A1(new_n893), .A2(new_n609), .A3(new_n604), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(G299), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n616), .A2(new_n580), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n892), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT41), .B1(new_n895), .B2(new_n896), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n895), .A2(KEYINPUT41), .A3(new_n896), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n897), .B1(new_n901), .B2(new_n892), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n591), .A2(G290), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n591), .A2(G290), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n527), .B(new_n525), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n591), .A2(G290), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n591), .A2(G290), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(G166), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(G288), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n905), .A2(new_n908), .A3(new_n798), .ZN(new_n911));
  AOI21_X1  g486(.A(KEYINPUT42), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n905), .A2(new_n908), .A3(new_n798), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n798), .B1(new_n905), .B2(new_n908), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n910), .A2(KEYINPUT103), .A3(new_n911), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n912), .B1(new_n918), .B2(KEYINPUT42), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n902), .B(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n891), .B1(new_n920), .B2(new_n890), .ZN(G295));
  OAI21_X1  g496(.A(new_n891), .B1(new_n920), .B2(new_n890), .ZN(G331));
  XNOR2_X1  g497(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n918), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n916), .A2(new_n917), .A3(KEYINPUT106), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n844), .A2(new_n553), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n838), .A2(new_n552), .A3(new_n551), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(G301), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(G301), .B1(new_n927), .B2(new_n928), .ZN(new_n931));
  OAI21_X1  g506(.A(G286), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(G171), .B1(new_n843), .B2(new_n845), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n933), .A2(G168), .A3(new_n929), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n900), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n935), .B1(new_n936), .B2(new_n898), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n895), .A2(new_n896), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n932), .A2(new_n938), .A3(new_n934), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n932), .A2(new_n938), .A3(new_n934), .A4(KEYINPUT105), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n937), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n925), .A2(new_n926), .A3(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n918), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n882), .B1(new_n945), .B2(new_n943), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n923), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n937), .A2(new_n941), .A3(new_n942), .ZN(new_n949));
  AOI21_X1  g524(.A(G37), .B1(new_n949), .B2(new_n918), .ZN(new_n950));
  INV_X1    g525(.A(new_n923), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n937), .A2(new_n939), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n925), .A2(new_n926), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n950), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n947), .A2(new_n948), .A3(new_n954), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n925), .A2(new_n926), .A3(new_n952), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT107), .B1(new_n956), .B2(new_n946), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT107), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n950), .A2(new_n958), .A3(new_n953), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n957), .A2(new_n959), .A3(KEYINPUT43), .ZN(new_n960));
  OR3_X1    g535(.A1(new_n944), .A2(new_n946), .A3(new_n923), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n955), .B1(new_n962), .B2(KEYINPUT44), .ZN(G397));
  NAND2_X1  g538(.A1(G286), .A2(G8), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT121), .ZN(new_n965));
  INV_X1    g540(.A(G1384), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n500), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G40), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n466), .A2(new_n970), .A3(new_n470), .ZN(new_n971));
  AOI21_X1  g546(.A(G1384), .B1(new_n489), .B2(new_n499), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT45), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n969), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G1966), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n967), .A2(KEYINPUT50), .ZN(new_n977));
  INV_X1    g552(.A(G2084), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n972), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n977), .A2(new_n978), .A3(new_n971), .A4(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT122), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n965), .A2(new_n976), .A3(new_n981), .A4(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT45), .B1(new_n500), .B2(new_n966), .ZN(new_n986));
  AOI211_X1 g561(.A(new_n968), .B(G1384), .C1(new_n489), .C2(new_n499), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(G1966), .B1(new_n988), .B2(new_n971), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n972), .A2(new_n979), .ZN(new_n990));
  AOI211_X1 g565(.A(KEYINPUT50), .B(G1384), .C1(new_n489), .C2(new_n499), .ZN(new_n991));
  INV_X1    g566(.A(new_n971), .ZN(new_n992));
  NOR4_X1   g567(.A1(new_n990), .A2(new_n991), .A3(G2084), .A4(new_n992), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n983), .B(G8), .C1(new_n989), .C2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n965), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n984), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n976), .A2(new_n981), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n997), .B1(new_n998), .B2(G8), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n985), .B1(new_n996), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT62), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n986), .A2(new_n987), .A3(new_n992), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT109), .B1(new_n1003), .B2(G1971), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n1005));
  INV_X1    g580(.A(G2090), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(KEYINPUT110), .A3(new_n1006), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n977), .A2(new_n1006), .A3(new_n971), .A4(new_n980), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT110), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT109), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n974), .A2(new_n1011), .A3(new_n804), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1004), .A2(new_n1007), .A3(new_n1010), .A4(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n525), .A2(new_n527), .A3(G8), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT55), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1013), .A2(G8), .A3(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1008), .B1(new_n1003), .B2(G1971), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1016), .B1(new_n1018), .B2(G8), .ZN(new_n1019));
  INV_X1    g594(.A(G8), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1020), .B1(new_n972), .B2(new_n971), .ZN(new_n1021));
  INV_X1    g596(.A(G1981), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n591), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT113), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT49), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT114), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(G1981), .B1(new_n588), .B2(new_n590), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1023), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1025), .A2(KEYINPUT114), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n1023), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1021), .B(new_n1028), .C1(new_n1030), .C2(new_n1026), .ZN(new_n1031));
  INV_X1    g606(.A(G1976), .ZN(new_n1032));
  NOR2_X1   g607(.A1(G288), .A2(new_n1032), .ZN(new_n1033));
  AOI211_X1 g608(.A(new_n1020), .B(new_n1033), .C1(new_n972), .C2(new_n971), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT112), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n1036));
  XOR2_X1   g611(.A(KEYINPUT111), .B(G1976), .Z(new_n1037));
  NAND2_X1  g612(.A1(G288), .A2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n500), .A2(new_n971), .A3(new_n966), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1033), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(G8), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1038), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n1042), .A2(KEYINPUT52), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT112), .B1(new_n1042), .B2(KEYINPUT52), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1031), .B(new_n1039), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1019), .A2(new_n1046), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n1017), .A2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n969), .A2(new_n768), .A3(new_n971), .A4(new_n973), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1049), .A2(KEYINPUT123), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1050), .B1(new_n1049), .B2(KEYINPUT123), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n977), .A2(new_n971), .A3(new_n980), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n740), .ZN(new_n1055));
  AOI21_X1  g630(.A(G301), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1002), .A2(new_n1048), .A3(KEYINPUT125), .A4(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT125), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1056), .A2(new_n1017), .A3(new_n1047), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1020), .B1(new_n976), .B2(new_n981), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n994), .B(new_n995), .C1(new_n1060), .C2(new_n997), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT62), .B1(new_n1061), .B2(new_n985), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1058), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1061), .A2(KEYINPUT62), .A3(new_n985), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1057), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1031), .A2(new_n1032), .A3(new_n798), .ZN(new_n1066));
  XOR2_X1   g641(.A(new_n1023), .B(KEYINPUT115), .Z(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT116), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1066), .A2(new_n1070), .A3(new_n1067), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1069), .A2(new_n1021), .A3(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(new_n1017), .B2(new_n1046), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT63), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1013), .A2(G8), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1016), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1046), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1077), .A2(G168), .A3(new_n1078), .A4(new_n1060), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1017), .A2(new_n1047), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1060), .A2(G168), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1074), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1073), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1040), .A2(G2067), .ZN(new_n1084));
  INV_X1    g659(.A(G1348), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1084), .B1(new_n1054), .B2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1086), .A2(new_n616), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1054), .A2(new_n788), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n579), .A2(new_n1089), .A3(new_n575), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1089), .B1(new_n579), .B2(new_n575), .ZN(new_n1092));
  NOR3_X1   g667(.A1(new_n1091), .A2(new_n573), .A3(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT118), .B1(new_n1093), .B2(KEYINPUT57), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1092), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n1090), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1095), .B(new_n1096), .C1(new_n1098), .C2(new_n573), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n580), .A2(KEYINPUT57), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1094), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT56), .B(G2072), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n988), .A2(new_n971), .A3(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1088), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1087), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1088), .A2(new_n1103), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1101), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1105), .A2(KEYINPUT119), .A3(new_n1108), .ZN(new_n1112));
  INV_X1    g687(.A(G1996), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n969), .A2(new_n1113), .A3(new_n971), .A4(new_n973), .ZN(new_n1114));
  XOR2_X1   g689(.A(KEYINPUT58), .B(G1341), .Z(new_n1115));
  NAND2_X1  g690(.A1(new_n1040), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT120), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1040), .A2(KEYINPUT120), .A3(new_n1115), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1114), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n554), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(KEYINPUT59), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT59), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1120), .A2(new_n1123), .A3(new_n554), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  AOI211_X1 g700(.A(new_n894), .B(new_n1084), .C1(new_n1054), .C2(new_n1085), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT60), .B1(new_n1087), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT60), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1086), .A2(new_n1128), .A3(new_n894), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1125), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT61), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1088), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1101), .B1(new_n1088), .B2(new_n1103), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1131), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1108), .A2(KEYINPUT61), .A3(new_n1104), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1111), .B(new_n1112), .C1(new_n1130), .C2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1017), .A2(new_n1061), .A3(new_n1047), .A4(new_n985), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT124), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT54), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1049), .A2(KEYINPUT123), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(KEYINPUT53), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1049), .A2(KEYINPUT123), .A3(new_n1050), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1143), .A2(new_n1055), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(G171), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1143), .A2(G301), .A3(new_n1055), .A4(new_n1144), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1141), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1138), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1147), .ZN(new_n1150));
  OAI22_X1  g725(.A1(new_n1056), .A2(new_n1150), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n1141), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1137), .A2(new_n1149), .A3(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1065), .A2(new_n1083), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n986), .A2(new_n971), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1155), .A2(G1996), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n725), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n1157), .A2(KEYINPUT108), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1155), .ZN(new_n1159));
  XOR2_X1   g734(.A(new_n710), .B(G2067), .Z(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n725), .A2(new_n1113), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1159), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1157), .A2(KEYINPUT108), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1158), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  XOR2_X1   g740(.A(new_n818), .B(new_n821), .Z(new_n1166));
  AND2_X1   g741(.A1(new_n1159), .A2(new_n1166), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(G290), .B(G1986), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1168), .B1(new_n1159), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1154), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n725), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1159), .B1(new_n1161), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1156), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n1174), .A2(KEYINPUT46), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1174), .A2(KEYINPUT46), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1173), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  XOR2_X1   g752(.A(new_n1177), .B(KEYINPUT47), .Z(new_n1178));
  NAND2_X1  g753(.A1(new_n819), .A2(new_n821), .ZN(new_n1179));
  OAI22_X1  g754(.A1(new_n1165), .A2(new_n1179), .B1(G2067), .B2(new_n710), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1180), .A2(new_n1159), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1168), .B(KEYINPUT126), .ZN(new_n1182));
  NOR3_X1   g757(.A1(new_n1155), .A2(G1986), .A3(G290), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT127), .ZN(new_n1184));
  XOR2_X1   g759(.A(new_n1184), .B(KEYINPUT48), .Z(new_n1185));
  AOI211_X1 g760(.A(new_n1178), .B(new_n1181), .C1(new_n1182), .C2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1171), .A2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g762(.A(G227), .B1(new_n947), .B2(new_n954), .ZN(new_n1189));
  INV_X1    g763(.A(G319), .ZN(new_n1190));
  NOR2_X1   g764(.A1(G401), .A2(new_n1190), .ZN(new_n1191));
  NAND4_X1  g765(.A1(new_n1189), .A2(new_n703), .A3(new_n888), .A4(new_n1191), .ZN(G225));
  INV_X1    g766(.A(G225), .ZN(G308));
endmodule


