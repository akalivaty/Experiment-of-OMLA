//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 0 1 0 0 1 1 0 0 1 1 0 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n757,
    new_n758, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1028, new_n1029, new_n1030, new_n1031;
  INV_X1    g000(.A(G148gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G141gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT76), .B(G141gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(new_n204), .B2(new_n202), .ZN(new_n205));
  NOR2_X1   g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT2), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G141gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G148gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n203), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g013(.A(new_n206), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n215), .A2(new_n209), .ZN(new_n216));
  AOI22_X1  g015(.A1(new_n205), .A2(new_n210), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G197gat), .B(G204gat), .ZN(new_n218));
  AND2_X1   g017(.A1(G211gat), .A2(G218gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n218), .B1(KEYINPUT22), .B2(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(G211gat), .B(G218gat), .Z(new_n221));
  XNOR2_X1  g020(.A(new_n220), .B(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT29), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n217), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n217), .A2(new_n225), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n222), .B1(new_n227), .B2(new_n223), .ZN(new_n228));
  OR3_X1    g027(.A1(new_n226), .A2(G78gat), .A3(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT31), .B(G50gat), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(G78gat), .B1(new_n226), .B2(new_n228), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n229), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G228gat), .A2(G233gat), .ZN(new_n235));
  INV_X1    g034(.A(G22gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n237), .B(G106gat), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n231), .B1(new_n229), .B2(new_n232), .ZN(new_n240));
  OR3_X1    g039(.A1(new_n234), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n239), .B1(new_n234), .B2(new_n240), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(G15gat), .B(G43gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(G71gat), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n246), .B(G99gat), .Z(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT72), .ZN(new_n249));
  NAND2_X1  g048(.A1(G183gat), .A2(G190gat), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT27), .ZN(new_n251));
  INV_X1    g050(.A(G183gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n254));
  AOI21_X1  g053(.A(G190gat), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT28), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n250), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  OR2_X1    g058(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n260), .A2(KEYINPUT27), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n259), .B1(new_n262), .B2(new_n253), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G169gat), .A2(G176gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(G169gat), .A2(G176gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT26), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT66), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n266), .A2(new_n267), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT66), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n271), .B(new_n265), .C1(new_n266), .C2(new_n267), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n269), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  AND2_X1   g072(.A1(G169gat), .A2(G176gat), .ZN(new_n274));
  INV_X1    g073(.A(G169gat), .ZN(new_n275));
  INV_X1    g074(.A(G176gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT23), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n274), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT24), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n250), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G190gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n252), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n281), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n278), .A2(G176gat), .ZN(new_n286));
  AND2_X1   g085(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n279), .A2(new_n285), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT25), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n291), .B1(new_n266), .B2(KEYINPUT23), .ZN(new_n293));
  AOI21_X1  g092(.A(G190gat), .B1(new_n260), .B2(new_n261), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n281), .A2(new_n284), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n279), .B(new_n293), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  AOI22_X1  g095(.A1(new_n264), .A2(new_n273), .B1(new_n292), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G127gat), .B(G134gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT70), .ZN(new_n299));
  OR2_X1    g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(G113gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G120gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT69), .B(G120gat), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n302), .B1(new_n303), .B2(new_n301), .ZN(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT71), .B(KEYINPUT1), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n298), .A2(new_n299), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n300), .A2(new_n304), .A3(new_n305), .A4(new_n306), .ZN(new_n307));
  XOR2_X1   g106(.A(KEYINPUT67), .B(G127gat), .Z(new_n308));
  INV_X1    g107(.A(KEYINPUT68), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n308), .A2(new_n309), .A3(G134gat), .ZN(new_n310));
  INV_X1    g109(.A(G134gat), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n309), .B1(G127gat), .B2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(KEYINPUT67), .B(G127gat), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n312), .B1(new_n313), .B2(new_n311), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT1), .ZN(new_n315));
  INV_X1    g114(.A(new_n302), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n301), .A2(G120gat), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n310), .A2(new_n314), .A3(new_n318), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n307), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n249), .B1(new_n297), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n297), .A2(new_n320), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n292), .A2(new_n296), .ZN(new_n323));
  INV_X1    g122(.A(new_n261), .ZN(new_n324));
  NOR2_X1   g123(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n325));
  NOR3_X1   g124(.A1(new_n324), .A2(new_n325), .A3(new_n251), .ZN(new_n326));
  NOR2_X1   g125(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n258), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n254), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n282), .B1(new_n329), .B2(new_n327), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n330), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n273), .A2(new_n328), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n323), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n307), .A2(new_n319), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(KEYINPUT72), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n321), .A2(new_n322), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(G227gat), .A2(G233gat), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT33), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n248), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT32), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n342), .B1(new_n336), .B2(new_n338), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n321), .A2(new_n335), .A3(new_n337), .A4(new_n322), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT34), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT33), .B1(new_n336), .B2(new_n338), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n343), .B1(new_n349), .B2(new_n248), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n345), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n348), .ZN(new_n352));
  NOR3_X1   g151(.A1(new_n343), .A2(new_n349), .A3(new_n248), .ZN(new_n353));
  AOI221_X4 g152(.A(new_n342), .B1(KEYINPUT33), .B2(new_n247), .C1(new_n336), .C2(new_n338), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n244), .A2(new_n351), .A3(new_n355), .ZN(new_n356));
  AND2_X1   g155(.A1(new_n211), .A2(KEYINPUT76), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n211), .A2(KEYINPUT76), .ZN(new_n358));
  OAI21_X1  g157(.A(G148gat), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n359), .A2(new_n203), .B1(new_n209), .B2(new_n208), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n215), .A2(new_n209), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n361), .B1(new_n213), .B2(new_n207), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT3), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n334), .A2(new_n227), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n307), .A2(new_n217), .A3(new_n319), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(KEYINPUT4), .A3(new_n365), .ZN(new_n366));
  XOR2_X1   g165(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n367));
  OR2_X1    g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G225gat), .A2(G233gat), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n371), .A2(KEYINPUT5), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n365), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n374), .B1(new_n364), .B2(new_n367), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT4), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n365), .A2(new_n376), .ZN(new_n377));
  NOR3_X1   g176(.A1(new_n375), .A2(new_n371), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n217), .B1(new_n319), .B2(new_n307), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n371), .B1(new_n374), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT5), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n373), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(G85gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(G1gat), .B(G29gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n384), .B(KEYINPUT0), .ZN(new_n385));
  INV_X1    g184(.A(G57gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n385), .A2(new_n386), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n383), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n389), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n391), .A2(new_n387), .A3(G85gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n382), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT6), .ZN(new_n395));
  INV_X1    g194(.A(new_n393), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n373), .B(new_n396), .C1(new_n378), .C2(new_n381), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n394), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n364), .A2(new_n367), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n371), .B1(new_n399), .B2(new_n365), .ZN(new_n400));
  INV_X1    g199(.A(new_n377), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n381), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n372), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n403), .B1(new_n366), .B2(new_n368), .ZN(new_n404));
  OAI211_X1 g203(.A(KEYINPUT6), .B(new_n393), .C1(new_n402), .C2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT78), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT78), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n382), .A2(new_n407), .A3(KEYINPUT6), .A4(new_n393), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n398), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n222), .ZN(new_n410));
  INV_X1    g209(.A(G226gat), .ZN(new_n411));
  INV_X1    g210(.A(G233gat), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n413), .A2(KEYINPUT29), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT74), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n273), .A2(new_n328), .A3(new_n331), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n265), .B1(new_n266), .B2(KEYINPUT23), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n281), .A2(new_n284), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n282), .B1(new_n324), .B2(new_n325), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AOI22_X1  g220(.A1(new_n421), .A2(new_n293), .B1(new_n290), .B2(new_n291), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n416), .B1(new_n417), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n323), .A2(KEYINPUT74), .A3(new_n332), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n415), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n297), .A2(new_n413), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n410), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n423), .A2(new_n413), .A3(new_n424), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n333), .A2(new_n414), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(new_n222), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT30), .ZN(new_n433));
  XNOR2_X1  g232(.A(G8gat), .B(G36gat), .ZN(new_n434));
  INV_X1    g233(.A(G64gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n434), .B(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(G92gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n436), .B(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n432), .A2(new_n433), .A3(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n438), .B(KEYINPUT75), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n428), .A2(new_n431), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT30), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n438), .B1(new_n428), .B2(new_n431), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n440), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n409), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT35), .B1(new_n356), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT87), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT73), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n355), .A2(new_n449), .A3(new_n351), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n345), .A2(KEYINPUT73), .A3(new_n348), .A4(new_n350), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n244), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT86), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n445), .A2(KEYINPUT80), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT80), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n456), .B(new_n440), .C1(new_n443), .C2(new_n444), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n399), .A2(new_n365), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n459), .A2(new_n370), .A3(new_n401), .ZN(new_n460));
  INV_X1    g259(.A(new_n381), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n404), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n390), .A2(new_n392), .A3(KEYINPUT81), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT81), .B1(new_n390), .B2(new_n392), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n397), .B(new_n395), .C1(new_n462), .C2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n406), .A2(new_n466), .A3(new_n408), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n454), .B1(new_n458), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n453), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n457), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n429), .A2(new_n222), .A3(new_n430), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n323), .A2(KEYINPUT74), .A3(new_n332), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT74), .B1(new_n323), .B2(new_n332), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n414), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n222), .B1(new_n474), .B2(new_n426), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n439), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n476), .A2(KEYINPUT30), .A3(new_n442), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n456), .B1(new_n477), .B2(new_n440), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n467), .B(new_n454), .C1(new_n470), .C2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT35), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n448), .B1(new_n469), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n467), .B1(new_n470), .B2(new_n478), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT86), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n243), .B1(new_n450), .B2(new_n451), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n484), .A2(new_n480), .A3(new_n485), .A4(new_n479), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n486), .A2(KEYINPUT87), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n447), .B1(new_n482), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT79), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT36), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n450), .A2(new_n490), .A3(new_n451), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n355), .A2(KEYINPUT36), .A3(new_n351), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n446), .A2(new_n243), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n489), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n374), .A2(new_n379), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT39), .B1(new_n497), .B2(new_n371), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT83), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g299(.A(KEYINPUT83), .B(KEYINPUT39), .C1(new_n497), .C2(new_n371), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n500), .B(new_n501), .C1(new_n370), .C2(new_n369), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT39), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n366), .A2(new_n503), .A3(new_n371), .A4(new_n368), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n465), .A2(KEYINPUT82), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT82), .B1(new_n465), .B2(new_n504), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n502), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT40), .ZN(new_n508));
  OR2_X1    g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n462), .A2(new_n465), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n510), .B1(new_n507), .B2(new_n508), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n509), .A2(new_n511), .A3(new_n457), .A4(new_n455), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n406), .A2(new_n408), .ZN(new_n513));
  XOR2_X1   g312(.A(KEYINPUT85), .B(KEYINPUT37), .Z(new_n514));
  NAND2_X1  g313(.A1(new_n432), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT37), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n515), .B(new_n438), .C1(new_n516), .C2(new_n432), .ZN(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT84), .B(KEYINPUT38), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n444), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n518), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n474), .A2(new_n222), .A3(new_n426), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n429), .A2(new_n430), .ZN(new_n522));
  OAI211_X1 g321(.A(KEYINPUT37), .B(new_n521), .C1(new_n522), .C2(new_n222), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n515), .A2(new_n441), .A3(new_n520), .A4(new_n523), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n513), .A2(new_n519), .A3(new_n466), .A4(new_n524), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n512), .A2(new_n525), .A3(new_n244), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n493), .A2(new_n489), .A3(new_n494), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n496), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n488), .A2(KEYINPUT88), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT88), .ZN(new_n531));
  INV_X1    g330(.A(new_n447), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n486), .A2(KEYINPUT87), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n481), .A2(new_n448), .A3(new_n485), .A4(new_n484), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n493), .A2(new_n489), .A3(new_n494), .ZN(new_n536));
  NOR3_X1   g335(.A1(new_n536), .A2(new_n495), .A3(new_n526), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n531), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  OR2_X1    g337(.A1(KEYINPUT89), .A2(G36gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(KEYINPUT89), .A2(G36gat), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n539), .A2(G29gat), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT14), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n542), .B1(G29gat), .B2(G36gat), .ZN(new_n543));
  INV_X1    g342(.A(G29gat), .ZN(new_n544));
  INV_X1    g343(.A(G36gat), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(new_n545), .A3(KEYINPUT14), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n541), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT15), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n541), .A2(KEYINPUT15), .A3(new_n543), .A4(new_n546), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G43gat), .B(G50gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT90), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT16), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n555), .A2(G1gat), .ZN(new_n556));
  INV_X1    g355(.A(G15gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(G22gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n236), .A2(G15gat), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n556), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(G1gat), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n561), .B1(new_n558), .B2(new_n559), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n554), .B(G8gat), .C1(new_n560), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n558), .A2(new_n559), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(G1gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n554), .A2(G8gat), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n556), .A2(new_n558), .A3(new_n559), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n554), .A2(G8gat), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n565), .A2(new_n566), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n563), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n552), .ZN(new_n572));
  AND2_X1   g371(.A1(new_n550), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n553), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT92), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n573), .B1(new_n551), .B2(new_n552), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT92), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n577), .A2(new_n578), .A3(new_n571), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT93), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n580), .B1(new_n577), .B2(new_n571), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n572), .B1(new_n549), .B2(new_n550), .ZN(new_n582));
  OAI211_X1 g381(.A(KEYINPUT93), .B(new_n570), .C1(new_n582), .C2(new_n573), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n576), .A2(new_n579), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G229gat), .A2(G233gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT13), .ZN(new_n586));
  NOR3_X1   g385(.A1(new_n584), .A2(KEYINPUT94), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT94), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n553), .A2(new_n574), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT93), .B1(new_n589), .B2(new_n570), .ZN(new_n590));
  INV_X1    g389(.A(new_n583), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n578), .B1(new_n577), .B2(new_n571), .ZN(new_n592));
  NOR4_X1   g391(.A1(new_n582), .A2(new_n570), .A3(new_n573), .A4(KEYINPUT92), .ZN(new_n593));
  OAI22_X1  g392(.A1(new_n590), .A2(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n586), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n588), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n587), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT17), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n553), .A2(new_n598), .A3(new_n574), .ZN(new_n599));
  OAI21_X1  g398(.A(KEYINPUT17), .B1(new_n582), .B2(new_n573), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(new_n600), .A3(new_n570), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n601), .A2(new_n585), .A3(new_n575), .ZN(new_n602));
  NOR2_X1   g401(.A1(KEYINPUT91), .A2(KEYINPUT18), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n601), .A2(new_n585), .A3(new_n575), .A4(new_n603), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n597), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G113gat), .B(G141gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(G197gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT11), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(new_n275), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT12), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n611), .B(G169gat), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT12), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n608), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(KEYINPUT94), .B1(new_n584), .B2(new_n586), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n594), .A2(new_n588), .A3(new_n595), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n607), .A2(new_n620), .A3(new_n617), .A4(new_n621), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n622), .A2(KEYINPUT95), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(KEYINPUT95), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n619), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT104), .ZN(new_n626));
  NAND2_X1  g425(.A1(G85gat), .A2(G92gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G99gat), .A2(G106gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(KEYINPUT8), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n383), .A2(new_n437), .ZN(new_n632));
  NAND4_X1  g431(.A1(KEYINPUT102), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n629), .A2(new_n631), .A3(new_n632), .A4(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT103), .ZN(new_n635));
  XOR2_X1   g434(.A(G99gat), .B(G106gat), .Z(new_n636));
  AOI22_X1  g435(.A1(KEYINPUT8), .A2(new_n630), .B1(new_n383), .B2(new_n437), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT103), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n637), .A2(new_n638), .A3(new_n629), .A4(new_n633), .ZN(new_n639));
  AND3_X1   g438(.A1(new_n635), .A2(new_n636), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n636), .B1(new_n635), .B2(new_n639), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n626), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n635), .A2(new_n639), .ZN(new_n643));
  INV_X1    g442(.A(new_n636), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n635), .A2(new_n636), .A3(new_n639), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n645), .A2(KEYINPUT104), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n648), .A2(new_n600), .A3(new_n599), .ZN(new_n649));
  NAND3_X1  g448(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n642), .A2(new_n647), .A3(new_n577), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(G134gat), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n649), .A2(new_n311), .A3(new_n650), .A4(new_n651), .ZN(new_n654));
  XNOR2_X1  g453(.A(G190gat), .B(G218gat), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n653), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(G162gat), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n656), .B1(new_n653), .B2(new_n654), .ZN(new_n662));
  OR3_X1    g461(.A1(new_n658), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n661), .B1(new_n658), .B2(new_n662), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g464(.A(G71gat), .B(G78gat), .Z(new_n666));
  NAND2_X1  g465(.A1(new_n435), .A2(G57gat), .ZN(new_n667));
  AND2_X1   g466(.A1(KEYINPUT97), .A2(G57gat), .ZN(new_n668));
  NOR2_X1   g467(.A1(KEYINPUT97), .A2(G57gat), .ZN(new_n669));
  OAI21_X1  g468(.A(G64gat), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n666), .B1(new_n667), .B2(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT96), .ZN(new_n673));
  AND2_X1   g472(.A1(G71gat), .A2(G78gat), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT96), .B1(new_n674), .B2(KEYINPUT9), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT96), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n386), .A2(G64gat), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n667), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n675), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  AOI22_X1  g479(.A1(new_n671), .A2(new_n673), .B1(new_n666), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(KEYINPUT21), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n570), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(KEYINPUT100), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT100), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n682), .A2(new_n685), .A3(new_n570), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT101), .B(KEYINPUT20), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n684), .A2(new_n686), .A3(new_n688), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(KEYINPUT99), .B(KEYINPUT19), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n691), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(G127gat), .B(G155gat), .ZN(new_n696));
  NAND2_X1  g495(.A1(G231gat), .A2(G233gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(G183gat), .B(G211gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n670), .A2(new_n667), .ZN(new_n701));
  INV_X1    g500(.A(new_n666), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n673), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n680), .A2(new_n666), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(KEYINPUT98), .B(KEYINPUT21), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n700), .B(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n694), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n709), .B1(new_n690), .B2(new_n692), .ZN(new_n710));
  OR3_X1    g509(.A1(new_n695), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n708), .B1(new_n695), .B2(new_n710), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n665), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n530), .A2(new_n538), .A3(new_n625), .A4(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n634), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n645), .A2(new_n681), .A3(new_n717), .A4(new_n646), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n704), .A3(new_n717), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n640), .B2(new_n641), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(G230gat), .A2(G233gat), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(G120gat), .B(G148gat), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(new_n276), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(G204gat), .ZN(new_n727));
  INV_X1    g526(.A(new_n722), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT10), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n718), .A2(new_n720), .A3(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n705), .A2(new_n729), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n642), .A2(new_n647), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n728), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI211_X1 g534(.A(KEYINPUT106), .B(new_n728), .C1(new_n730), .C2(new_n732), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n724), .B(new_n727), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n727), .B(KEYINPUT107), .Z(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n723), .B2(new_n733), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n715), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n409), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g543(.A(KEYINPUT16), .B(G8gat), .ZN(new_n745));
  NOR4_X1   g544(.A1(new_n715), .A2(new_n740), .A3(new_n458), .A4(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n747));
  OR3_X1    g546(.A1(new_n746), .A2(new_n747), .A3(KEYINPUT42), .ZN(new_n748));
  INV_X1    g547(.A(new_n458), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n741), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(G8gat), .ZN(new_n751));
  OAI21_X1  g550(.A(KEYINPUT42), .B1(new_n746), .B2(new_n747), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n748), .A2(new_n751), .A3(new_n752), .ZN(G1325gat));
  AOI21_X1  g552(.A(G15gat), .B1(new_n741), .B2(new_n452), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n493), .A2(new_n557), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n754), .B1(new_n741), .B2(new_n755), .ZN(G1326gat));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n243), .ZN(new_n757));
  XNOR2_X1  g556(.A(KEYINPUT43), .B(G22gat), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(G1327gat));
  INV_X1    g558(.A(new_n740), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n665), .A2(new_n760), .A3(new_n713), .ZN(new_n761));
  XOR2_X1   g560(.A(new_n761), .B(KEYINPUT109), .Z(new_n762));
  AND4_X1   g561(.A1(new_n530), .A2(new_n538), .A3(new_n625), .A4(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n763), .A2(new_n544), .A3(new_n742), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT45), .ZN(new_n765));
  INV_X1    g564(.A(new_n665), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT44), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n530), .A2(new_n538), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n493), .A2(new_n494), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n526), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n665), .B1(new_n535), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n767), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n713), .B(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT95), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n597), .A2(new_n776), .A3(new_n617), .A4(new_n607), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n622), .A2(KEYINPUT95), .ZN(new_n778));
  AOI22_X1  g577(.A1(new_n777), .A2(new_n778), .B1(new_n608), .B2(new_n618), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n775), .A2(new_n740), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT111), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n769), .A2(new_n773), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(G29gat), .B1(new_n782), .B2(new_n409), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n765), .A2(new_n783), .ZN(G1328gat));
  NAND2_X1  g583(.A1(new_n539), .A2(new_n540), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n763), .A2(new_n749), .A3(new_n785), .ZN(new_n786));
  OR2_X1    g585(.A1(new_n786), .A2(KEYINPUT46), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(KEYINPUT46), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n782), .A2(new_n458), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n787), .B(new_n788), .C1(new_n785), .C2(new_n789), .ZN(G1329gat));
  INV_X1    g589(.A(new_n493), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n769), .A2(new_n791), .A3(new_n773), .A4(new_n781), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(G43gat), .ZN(new_n793));
  INV_X1    g592(.A(new_n452), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n794), .A2(G43gat), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n763), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT112), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT47), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AOI22_X1  g598(.A1(new_n792), .A2(G43gat), .B1(new_n763), .B2(new_n795), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT47), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n800), .A2(KEYINPUT112), .A3(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n799), .A2(new_n802), .ZN(G1330gat));
  NAND4_X1  g602(.A1(new_n769), .A2(new_n243), .A3(new_n773), .A4(new_n781), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(G50gat), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n530), .A2(new_n538), .A3(new_n625), .A4(new_n762), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n244), .A2(G50gat), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n806), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n763), .A2(KEYINPUT113), .A3(new_n808), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n805), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT48), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n763), .B2(new_n808), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n805), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n813), .B1(new_n805), .B2(new_n815), .ZN(new_n817));
  OAI22_X1  g616(.A1(KEYINPUT48), .A2(new_n812), .B1(new_n816), .B2(new_n817), .ZN(G1331gat));
  NOR3_X1   g617(.A1(new_n665), .A2(new_n625), .A3(new_n713), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n740), .B(new_n819), .C1(new_n535), .C2(new_n771), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n742), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n668), .A2(new_n669), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n826), .B(new_n827), .ZN(G1332gat));
  NAND2_X1  g627(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n822), .A2(new_n749), .A3(new_n823), .A4(new_n829), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n830), .A2(KEYINPUT116), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n830), .A2(KEYINPUT116), .ZN(new_n832));
  OAI22_X1  g631(.A1(new_n831), .A2(new_n832), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n830), .A2(KEYINPUT116), .ZN(new_n834));
  NOR2_X1   g633(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n830), .A2(KEYINPUT116), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n833), .A2(new_n837), .ZN(G1333gat));
  INV_X1    g637(.A(G71gat), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n839), .B1(new_n824), .B2(new_n794), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n822), .A2(G71gat), .A3(new_n791), .A4(new_n823), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(KEYINPUT50), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT50), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n840), .A2(new_n844), .A3(new_n841), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(G1334gat));
  NAND2_X1  g645(.A1(new_n825), .A2(new_n243), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g647(.A1(new_n779), .A2(new_n713), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n769), .A2(new_n773), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n409), .A2(new_n760), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(G85gat), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n665), .B(new_n850), .C1(new_n535), .C2(new_n771), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT51), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n855), .B(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(new_n383), .A3(new_n852), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n854), .A2(new_n858), .ZN(G1336gat));
  NAND4_X1  g658(.A1(new_n769), .A2(new_n740), .A3(new_n773), .A4(new_n850), .ZN(new_n860));
  OAI21_X1  g659(.A(G92gat), .B1(new_n860), .B2(new_n458), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n458), .A2(G92gat), .A3(new_n760), .ZN(new_n862));
  AOI22_X1  g661(.A1(new_n857), .A2(new_n862), .B1(KEYINPUT117), .B2(KEYINPUT52), .ZN(new_n863));
  OR2_X1    g662(.A1(KEYINPUT117), .A2(KEYINPUT52), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n861), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n864), .B1(new_n861), .B2(new_n863), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(G1337gat));
  OAI21_X1  g666(.A(G99gat), .B1(new_n860), .B2(new_n493), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n760), .A2(G99gat), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n857), .A2(new_n452), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(G1338gat));
  OAI21_X1  g670(.A(G106gat), .B1(new_n860), .B2(new_n244), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n244), .A2(new_n760), .A3(G106gat), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT118), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n857), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT53), .ZN(new_n877));
  INV_X1    g676(.A(new_n873), .ZN(new_n878));
  OR2_X1    g677(.A1(new_n855), .A2(new_n856), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n855), .A2(new_n856), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT53), .B1(new_n881), .B2(KEYINPUT119), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n857), .A2(new_n873), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n882), .A2(new_n885), .A3(new_n872), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n877), .A2(new_n886), .ZN(G1339gat));
  NAND2_X1  g686(.A1(new_n584), .A2(new_n586), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n601), .A2(new_n575), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(G229gat), .A3(G233gat), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n614), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n891), .B1(new_n777), .B2(new_n778), .ZN(new_n892));
  INV_X1    g691(.A(new_n737), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n730), .A2(new_n732), .A3(new_n728), .ZN(new_n894));
  OAI211_X1 g693(.A(KEYINPUT54), .B(new_n894), .C1(new_n735), .C2(new_n736), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n727), .B1(new_n733), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT55), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT55), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n895), .A2(new_n900), .A3(new_n897), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n893), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n665), .A2(new_n892), .A3(new_n902), .ZN(new_n903));
  AOI22_X1  g702(.A1(new_n625), .A2(new_n902), .B1(new_n892), .B2(new_n740), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n903), .B1(new_n904), .B2(new_n665), .ZN(new_n905));
  INV_X1    g704(.A(new_n775), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR4_X1   g706(.A1(new_n665), .A2(new_n625), .A3(new_n740), .A4(new_n713), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n749), .A2(new_n409), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n912), .A2(new_n453), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(G113gat), .B1(new_n914), .B2(new_n779), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n912), .A2(new_n356), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n301), .A3(new_n625), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(G1340gat));
  OAI21_X1  g717(.A(G120gat), .B1(new_n914), .B2(new_n760), .ZN(new_n919));
  INV_X1    g718(.A(new_n303), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n916), .A2(new_n920), .A3(new_n740), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(G1341gat));
  INV_X1    g721(.A(new_n713), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n313), .B1(new_n916), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n906), .A2(new_n308), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n924), .B1(new_n913), .B2(new_n925), .ZN(G1342gat));
  NAND3_X1  g725(.A1(new_n916), .A2(new_n311), .A3(new_n665), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT56), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n912), .A2(new_n766), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n311), .B1(new_n929), .B2(new_n485), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n928), .A2(new_n930), .ZN(G1343gat));
  INV_X1    g730(.A(KEYINPUT121), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n244), .B1(new_n907), .B2(new_n909), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n911), .A2(new_n493), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n933), .A2(new_n211), .A3(new_n625), .A4(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT58), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n908), .B1(new_n905), .B2(new_n713), .ZN(new_n938));
  OAI21_X1  g737(.A(KEYINPUT57), .B1(new_n938), .B2(new_n244), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT57), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n895), .A2(new_n900), .A3(new_n897), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n900), .B1(new_n895), .B2(new_n897), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n737), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n779), .A2(new_n943), .ZN(new_n944));
  AOI221_X4 g743(.A(new_n891), .B1(new_n737), .B2(new_n739), .C1(new_n777), .C2(new_n778), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n766), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n775), .B1(new_n946), .B2(new_n903), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n940), .B(new_n243), .C1(new_n947), .C2(new_n908), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n939), .A2(new_n625), .A3(new_n948), .A4(new_n934), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT120), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n937), .B1(new_n950), .B2(new_n204), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n204), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n936), .B1(new_n952), .B2(new_n935), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n932), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT120), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n949), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n949), .A2(new_n955), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n956), .A2(new_n204), .A3(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(new_n937), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(new_n953), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n960), .A2(new_n961), .A3(KEYINPUT121), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n954), .A2(new_n962), .ZN(G1344gat));
  AND2_X1   g762(.A1(new_n933), .A2(KEYINPUT57), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n938), .A2(new_n244), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n965), .A2(KEYINPUT57), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n934), .A2(new_n740), .ZN(new_n968));
  OAI211_X1 g767(.A(KEYINPUT59), .B(G148gat), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n933), .A2(new_n202), .A3(new_n740), .A4(new_n934), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n939), .A2(new_n934), .A3(new_n948), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n971), .A2(new_n760), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n972), .A2(new_n202), .ZN(new_n973));
  OAI211_X1 g772(.A(new_n969), .B(new_n970), .C1(KEYINPUT59), .C2(new_n973), .ZN(G1345gat));
  INV_X1    g773(.A(G155gat), .ZN(new_n975));
  NOR3_X1   g774(.A1(new_n971), .A2(new_n975), .A3(new_n906), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n933), .A2(new_n923), .A3(new_n934), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n976), .B1(new_n975), .B2(new_n977), .ZN(G1346gat));
  NOR2_X1   g777(.A1(new_n244), .A2(G162gat), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n929), .A2(new_n493), .A3(new_n979), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n980), .B(KEYINPUT122), .ZN(new_n981));
  OAI21_X1  g780(.A(G162gat), .B1(new_n971), .B2(new_n766), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(G1347gat));
  NOR2_X1   g782(.A1(new_n742), .A2(new_n458), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n910), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n985), .A2(new_n356), .ZN(new_n986));
  OAI211_X1 g785(.A(new_n986), .B(new_n625), .C1(new_n288), .C2(new_n287), .ZN(new_n987));
  XOR2_X1   g786(.A(new_n987), .B(KEYINPUT123), .Z(new_n988));
  NAND3_X1  g787(.A1(new_n910), .A2(new_n485), .A3(new_n984), .ZN(new_n989));
  OAI21_X1  g788(.A(G169gat), .B1(new_n989), .B2(new_n779), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n988), .A2(new_n990), .ZN(G1348gat));
  NOR3_X1   g790(.A1(new_n989), .A2(new_n276), .A3(new_n760), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n986), .A2(new_n740), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n992), .B1(new_n993), .B2(new_n276), .ZN(G1349gat));
  OAI211_X1 g793(.A(new_n986), .B(new_n923), .C1(new_n327), .C2(new_n329), .ZN(new_n995));
  OAI211_X1 g794(.A(new_n260), .B(new_n261), .C1(new_n989), .C2(new_n906), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  XNOR2_X1  g796(.A(new_n997), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g797(.A(G190gat), .B1(new_n989), .B2(new_n766), .ZN(new_n999));
  AOI21_X1  g798(.A(new_n999), .B1(KEYINPUT124), .B2(KEYINPUT61), .ZN(new_n1000));
  NOR2_X1   g799(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n1001));
  XNOR2_X1  g800(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n986), .A2(new_n282), .A3(new_n665), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1002), .A2(new_n1003), .ZN(G1351gat));
  INV_X1    g803(.A(KEYINPUT126), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n967), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n493), .A2(new_n984), .ZN(new_n1007));
  INV_X1    g806(.A(new_n1007), .ZN(new_n1008));
  OAI21_X1  g807(.A(KEYINPUT126), .B1(new_n964), .B2(new_n966), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n1006), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  OAI21_X1  g809(.A(G197gat), .B1(new_n1010), .B2(new_n779), .ZN(new_n1011));
  AND2_X1   g810(.A1(new_n933), .A2(new_n1008), .ZN(new_n1012));
  XNOR2_X1  g811(.A(new_n1012), .B(KEYINPUT125), .ZN(new_n1013));
  INV_X1    g812(.A(G197gat), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n1013), .A2(new_n1014), .A3(new_n625), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1011), .A2(new_n1015), .ZN(G1352gat));
  OAI21_X1  g815(.A(G204gat), .B1(new_n1010), .B2(new_n760), .ZN(new_n1017));
  INV_X1    g816(.A(G204gat), .ZN(new_n1018));
  NAND3_X1  g817(.A1(new_n1012), .A2(new_n1018), .A3(new_n740), .ZN(new_n1019));
  XOR2_X1   g818(.A(new_n1019), .B(KEYINPUT62), .Z(new_n1020));
  NAND2_X1  g819(.A1(new_n1017), .A2(new_n1020), .ZN(G1353gat));
  INV_X1    g820(.A(G211gat), .ZN(new_n1022));
  NAND3_X1  g821(.A1(new_n1013), .A2(new_n1022), .A3(new_n923), .ZN(new_n1023));
  OAI211_X1 g822(.A(new_n923), .B(new_n1008), .C1(new_n964), .C2(new_n966), .ZN(new_n1024));
  AND3_X1   g823(.A1(new_n1024), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1025));
  AOI21_X1  g824(.A(KEYINPUT63), .B1(new_n1024), .B2(G211gat), .ZN(new_n1026));
  OAI21_X1  g825(.A(new_n1023), .B1(new_n1025), .B2(new_n1026), .ZN(G1354gat));
  AOI21_X1  g826(.A(G218gat), .B1(new_n1013), .B2(new_n665), .ZN(new_n1028));
  INV_X1    g827(.A(new_n1010), .ZN(new_n1029));
  NAND2_X1  g828(.A1(new_n665), .A2(G218gat), .ZN(new_n1030));
  XNOR2_X1  g829(.A(new_n1030), .B(KEYINPUT127), .ZN(new_n1031));
  AOI21_X1  g830(.A(new_n1028), .B1(new_n1029), .B2(new_n1031), .ZN(G1355gat));
endmodule


