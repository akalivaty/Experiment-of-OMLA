//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 0 0 0 0 0 1 1 1 0 1 1 0 0 1 1 1 1 0 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n840, new_n841, new_n842,
    new_n843, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(G29gat), .A2(G36gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT14), .ZN(new_n204));
  NAND2_X1  g003(.A1(G29gat), .A2(G36gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  OAI211_X1 g005(.A(KEYINPUT15), .B(new_n202), .C1(new_n204), .C2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT89), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  XOR2_X1   g010(.A(new_n205), .B(KEYINPUT90), .Z(new_n212));
  NOR2_X1   g011(.A1(new_n212), .A2(new_n204), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  AND2_X1   g013(.A1(new_n214), .A2(KEYINPUT91), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(KEYINPUT91), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n207), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT17), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G15gat), .B(G22gat), .ZN(new_n220));
  INV_X1    g019(.A(G1gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT16), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(G1gat), .B2(new_n220), .ZN(new_n224));
  INV_X1    g023(.A(G8gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n224), .B(new_n225), .ZN(new_n226));
  OAI211_X1 g025(.A(KEYINPUT17), .B(new_n207), .C1(new_n215), .C2(new_n216), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n219), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G229gat), .A2(G233gat), .ZN(new_n229));
  INV_X1    g028(.A(new_n226), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n217), .A2(new_n230), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n228), .A2(KEYINPUT18), .A3(new_n229), .A4(new_n231), .ZN(new_n232));
  XOR2_X1   g031(.A(new_n229), .B(KEYINPUT13), .Z(new_n233));
  INV_X1    g032(.A(new_n231), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n217), .A2(new_n230), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G113gat), .B(G141gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(G169gat), .B(G197gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n241), .B(KEYINPUT12), .Z(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n232), .A2(new_n236), .A3(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n228), .A2(new_n229), .A3(new_n231), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT18), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT92), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT92), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n245), .A2(new_n249), .A3(new_n246), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n244), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n247), .A2(new_n232), .A3(new_n236), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(new_n242), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G230gat), .ZN(new_n256));
  INV_X1    g055(.A(G233gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(G85gat), .ZN(new_n259));
  INV_X1    g058(.A(G92gat), .ZN(new_n260));
  OAI21_X1  g059(.A(KEYINPUT98), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT98), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n262), .A2(G85gat), .A3(G92gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n261), .A2(KEYINPUT7), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G99gat), .A2(G106gat), .ZN(new_n265));
  AOI22_X1  g064(.A1(KEYINPUT8), .A2(new_n265), .B1(new_n259), .B2(new_n260), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT7), .ZN(new_n267));
  OAI211_X1 g066(.A(KEYINPUT98), .B(new_n267), .C1(new_n259), .C2(new_n260), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n264), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  XOR2_X1   g068(.A(G99gat), .B(G106gat), .Z(new_n270));
  XOR2_X1   g069(.A(new_n269), .B(new_n270), .Z(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT93), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G71gat), .B(G78gat), .ZN(new_n276));
  INV_X1    g075(.A(G64gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(G57gat), .ZN(new_n278));
  OR2_X1    g077(.A1(new_n277), .A2(G57gat), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n276), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT94), .B(G57gat), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n278), .B1(new_n281), .B2(new_n277), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT95), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n275), .B(new_n280), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n275), .A2(new_n282), .A3(new_n284), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(new_n276), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT100), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n269), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n272), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT10), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n271), .A2(new_n288), .A3(new_n290), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n271), .A2(KEYINPUT10), .A3(new_n288), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n258), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n292), .A2(new_n294), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(new_n258), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G120gat), .B(G148gat), .ZN(new_n302));
  INV_X1    g101(.A(G176gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G204gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n304), .B(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n306), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n298), .A2(new_n300), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G127gat), .B(G134gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT71), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT1), .ZN(new_n314));
  INV_X1    g113(.A(G113gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n315), .A2(G120gat), .ZN(new_n316));
  INV_X1    g115(.A(G120gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n317), .A2(G113gat), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n314), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT72), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n316), .B1(new_n321), .B2(new_n318), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT72), .B1(new_n317), .B2(G113gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n324), .A2(new_n314), .A3(new_n311), .ZN(new_n325));
  AND2_X1   g124(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G155gat), .ZN(new_n327));
  INV_X1    g126(.A(G162gat), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT2), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT77), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  XOR2_X1   g130(.A(G141gat), .B(G148gat), .Z(new_n332));
  XNOR2_X1  g131(.A(G155gat), .B(G162gat), .ZN(new_n333));
  OAI211_X1 g132(.A(KEYINPUT77), .B(KEYINPUT2), .C1(new_n327), .C2(new_n328), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n331), .A2(new_n332), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n333), .ZN(new_n336));
  XNOR2_X1  g135(.A(G141gat), .B(G148gat), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n336), .B1(KEYINPUT2), .B2(new_n337), .ZN(new_n338));
  AND2_X1   g137(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n326), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n340), .A2(KEYINPUT4), .ZN(new_n341));
  NAND2_X1  g140(.A1(G225gat), .A2(G233gat), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n320), .A2(new_n325), .ZN(new_n344));
  INV_X1    g143(.A(new_n339), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n340), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n341), .B1(new_n343), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n345), .A2(KEYINPUT3), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT3), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n339), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(new_n344), .A3(new_n351), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n352), .A2(KEYINPUT4), .A3(new_n340), .A4(new_n342), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n348), .A2(KEYINPUT5), .A3(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(KEYINPUT0), .B(G57gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(G85gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(G1gat), .B(G29gat), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n356), .B(new_n357), .Z(new_n358));
  AOI21_X1  g157(.A(KEYINPUT78), .B1(new_n340), .B2(KEYINPUT4), .ZN(new_n359));
  OR3_X1    g158(.A1(new_n344), .A2(new_n345), .A3(KEYINPUT4), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n341), .A2(KEYINPUT78), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n343), .A2(KEYINPUT5), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n361), .A2(new_n362), .A3(new_n352), .A4(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n354), .A2(new_n358), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT6), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n358), .B1(new_n354), .B2(new_n364), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI211_X1 g168(.A(new_n366), .B(new_n358), .C1(new_n354), .C2(new_n364), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G8gat), .B(G36gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n372), .B(new_n277), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n373), .B(new_n260), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(G211gat), .ZN(new_n376));
  INV_X1    g175(.A(G218gat), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT22), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n378), .B1(new_n376), .B2(new_n377), .ZN(new_n379));
  XNOR2_X1  g178(.A(G197gat), .B(G204gat), .ZN(new_n380));
  AND2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n380), .A2(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n376), .A2(new_n377), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n381), .B1(new_n384), .B2(KEYINPUT75), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n381), .A2(KEYINPUT75), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT76), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT64), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT23), .ZN(new_n391));
  INV_X1    g190(.A(G169gat), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n392), .A3(new_n303), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AND2_X1   g194(.A1(G169gat), .A2(G176gat), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n390), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  AOI211_X1 g197(.A(KEYINPUT64), .B(new_n396), .C1(new_n393), .C2(new_n394), .ZN(new_n399));
  NAND2_X1  g198(.A1(G183gat), .A2(G190gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT24), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT24), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(G183gat), .A3(G190gat), .ZN(new_n403));
  INV_X1    g202(.A(G183gat), .ZN(new_n404));
  INV_X1    g203(.A(G190gat), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n401), .A2(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NOR3_X1   g205(.A1(new_n398), .A2(new_n399), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n396), .B1(new_n393), .B2(new_n394), .ZN(new_n408));
  XNOR2_X1  g207(.A(KEYINPUT66), .B(G183gat), .ZN(new_n409));
  AND2_X1   g208(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n410));
  NOR2_X1   g209(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT65), .ZN(new_n413));
  NOR3_X1   g212(.A1(new_n400), .A2(new_n413), .A3(KEYINPUT24), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n402), .A2(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n415));
  OAI22_X1  g214(.A1(new_n409), .A2(new_n412), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n408), .B1(new_n416), .B2(KEYINPUT68), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n404), .A2(KEYINPUT66), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT66), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(G183gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT67), .B(G190gat), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n400), .B1(new_n413), .B2(KEYINPUT24), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n402), .A2(KEYINPUT65), .A3(G183gat), .A4(G190gat), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n421), .A2(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT68), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT25), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  OAI22_X1  g226(.A1(new_n407), .A2(KEYINPUT25), .B1(new_n417), .B2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(KEYINPUT27), .B(G183gat), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n422), .A2(new_n429), .A3(KEYINPUT28), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n418), .A2(new_n420), .A3(KEYINPUT27), .ZN(new_n431));
  OR2_X1    g230(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n412), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n430), .B1(new_n433), .B2(KEYINPUT28), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n392), .A2(new_n303), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT26), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n400), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n396), .A2(KEYINPUT26), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n437), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n428), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G226gat), .A2(G233gat), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n389), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT69), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n428), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n394), .ZN(new_n447));
  NOR3_X1   g246(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n397), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT64), .ZN(new_n450));
  INV_X1    g249(.A(new_n406), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n408), .A2(new_n390), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT25), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n454), .B1(new_n416), .B2(KEYINPUT68), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n449), .B1(new_n425), .B2(new_n426), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n455), .A2(new_n458), .A3(KEYINPUT69), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n446), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n440), .A2(KEYINPUT70), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT70), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n434), .A2(new_n462), .A3(new_n439), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT29), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n444), .B1(new_n465), .B2(new_n443), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n455), .A2(new_n458), .A3(KEYINPUT69), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT69), .B1(new_n455), .B2(new_n458), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n464), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT29), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n471), .A2(new_n389), .A3(new_n442), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n388), .B1(new_n466), .B2(new_n472), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n464), .B(new_n443), .C1(new_n467), .C2(new_n468), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n441), .A2(new_n470), .A3(new_n442), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(new_n388), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n375), .B1(new_n473), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT38), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT37), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n474), .A2(new_n387), .A3(new_n475), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT85), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT85), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n474), .A2(new_n483), .A3(new_n387), .A4(new_n475), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n441), .A2(new_n443), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT76), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n488), .B1(new_n471), .B2(new_n442), .ZN(new_n489));
  AOI211_X1 g288(.A(KEYINPUT76), .B(new_n443), .C1(new_n469), .C2(new_n470), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n388), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n480), .B1(new_n486), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT86), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n479), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n387), .B1(new_n466), .B2(new_n472), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n493), .B(KEYINPUT37), .C1(new_n495), .C2(new_n485), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n480), .B1(new_n473), .B2(new_n477), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(new_n374), .A3(new_n497), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n371), .B(new_n478), .C1(new_n494), .C2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT87), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n387), .B1(new_n489), .B2(new_n490), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(new_n476), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n375), .B1(new_n503), .B2(new_n480), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n504), .B1(new_n480), .B2(new_n503), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT38), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT37), .B1(new_n495), .B2(new_n485), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT38), .B1(new_n507), .B2(KEYINPUT86), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n508), .A2(new_n504), .A3(new_n496), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n509), .A2(KEYINPUT87), .A3(new_n371), .A4(new_n478), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n501), .A2(new_n506), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n502), .A2(new_n476), .A3(new_n374), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n478), .A2(KEYINPUT30), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT30), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n503), .A2(new_n514), .A3(new_n375), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT83), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n513), .A2(KEYINPUT83), .A3(new_n515), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n362), .A2(new_n352), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n342), .B1(new_n521), .B2(new_n361), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT39), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(new_n358), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n347), .A2(new_n343), .ZN(new_n526));
  NOR3_X1   g325(.A1(new_n522), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT84), .B1(new_n528), .B2(KEYINPUT40), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n368), .B1(new_n528), .B2(KEYINPUT40), .ZN(new_n530));
  OR3_X1    g329(.A1(new_n528), .A2(KEYINPUT84), .A3(KEYINPUT40), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n520), .A2(new_n529), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(G22gat), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n470), .B1(new_n385), .B2(new_n386), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n339), .B1(new_n534), .B2(new_n350), .ZN(new_n535));
  AOI211_X1 g334(.A(new_n386), .B(new_n385), .C1(new_n351), .C2(new_n470), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n537), .A2(G228gat), .A3(G233gat), .ZN(new_n538));
  INV_X1    g337(.A(G228gat), .ZN(new_n539));
  OAI22_X1  g338(.A1(new_n535), .A2(new_n536), .B1(new_n539), .B2(new_n257), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n533), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n538), .A2(new_n533), .A3(new_n540), .ZN(new_n543));
  XNOR2_X1  g342(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(G50gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(G78gat), .ZN(new_n546));
  XOR2_X1   g345(.A(new_n546), .B(G106gat), .Z(new_n547));
  NAND3_X1  g346(.A1(new_n542), .A2(new_n543), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT81), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n543), .B1(new_n541), .B2(new_n550), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n538), .A2(KEYINPUT81), .A3(new_n533), .A4(new_n540), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n547), .B(KEYINPUT80), .Z(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT82), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n553), .A2(KEYINPUT82), .A3(new_n554), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n549), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n511), .A2(new_n532), .A3(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(G15gat), .B(G43gat), .Z(new_n562));
  XNOR2_X1  g361(.A(G71gat), .B(G99gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  AND2_X1   g363(.A1(G227gat), .A2(G233gat), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n469), .A2(new_n344), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n460), .A2(new_n326), .A3(new_n464), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n564), .B1(new_n569), .B2(KEYINPUT33), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT32), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n570), .A2(new_n572), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n567), .A2(new_n568), .A3(new_n566), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT74), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT34), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n577), .A2(KEYINPUT34), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n576), .A2(new_n580), .A3(new_n578), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT73), .ZN(new_n584));
  AOI22_X1  g383(.A1(new_n573), .A2(new_n575), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n573), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n579), .A2(new_n581), .A3(new_n584), .ZN(new_n587));
  NOR3_X1   g386(.A1(new_n586), .A2(new_n587), .A3(new_n574), .ZN(new_n588));
  OAI21_X1  g387(.A(KEYINPUT36), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n582), .B1(new_n586), .B2(new_n574), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n575), .A2(new_n583), .A3(new_n573), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT36), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n371), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(new_n516), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n559), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n561), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  NOR3_X1   g397(.A1(new_n520), .A2(new_n559), .A3(new_n371), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT35), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n590), .A2(new_n591), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n585), .A2(new_n588), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n560), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(KEYINPUT35), .B1(new_n604), .B2(new_n596), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  AOI211_X1 g405(.A(new_n255), .B(new_n310), .C1(new_n598), .C2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G134gat), .B(G162gat), .ZN(new_n608));
  AOI21_X1  g407(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n608), .B(new_n609), .Z(new_n610));
  NAND3_X1  g409(.A1(new_n219), .A2(new_n272), .A3(new_n227), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT99), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AND3_X1   g412(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n614), .B1(new_n217), .B2(new_n271), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n219), .A2(new_n227), .A3(KEYINPUT99), .A4(new_n272), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n613), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(G190gat), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n613), .A2(new_n405), .A3(new_n615), .A4(new_n616), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n618), .A2(G218gat), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(G218gat), .B1(new_n618), .B2(new_n619), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n610), .B1(new_n622), .B2(KEYINPUT97), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n618), .A2(new_n619), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(new_n377), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n618), .A2(G218gat), .A3(new_n619), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n625), .A2(KEYINPUT97), .A3(new_n626), .A4(new_n610), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n230), .B1(KEYINPUT21), .B2(new_n288), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(new_n404), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G127gat), .B(G155gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(new_n376), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n634), .B(new_n636), .Z(new_n637));
  NOR2_X1   g436(.A1(new_n288), .A2(KEYINPUT21), .ZN(new_n638));
  NAND2_X1  g437(.A1(G231gat), .A2(G233gat), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n639), .B(KEYINPUT96), .Z(new_n640));
  XNOR2_X1  g439(.A(new_n638), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n637), .B(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n630), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n607), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n645), .A2(new_n595), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT101), .B(G1gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(G1324gat));
  INV_X1    g447(.A(new_n645), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n520), .ZN(new_n650));
  NOR2_X1   g449(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT42), .ZN(new_n653));
  NAND2_X1  g452(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n654));
  AND3_X1   g453(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n653), .B1(new_n652), .B2(new_n654), .ZN(new_n656));
  AND3_X1   g455(.A1(new_n650), .A2(KEYINPUT102), .A3(G8gat), .ZN(new_n657));
  AOI21_X1  g456(.A(KEYINPUT102), .B1(new_n650), .B2(G8gat), .ZN(new_n658));
  OAI22_X1  g457(.A1(new_n655), .A2(new_n656), .B1(new_n657), .B2(new_n658), .ZN(G1325gat));
  AOI21_X1  g458(.A(G15gat), .B1(new_n649), .B2(new_n601), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT103), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n589), .A2(new_n593), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n661), .B1(new_n589), .B2(new_n593), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n645), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n660), .B1(G15gat), .B2(new_n665), .ZN(G1326gat));
  NOR2_X1   g465(.A1(new_n645), .A2(new_n560), .ZN(new_n667));
  XOR2_X1   g466(.A(KEYINPUT43), .B(G22gat), .Z(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1327gat));
  NAND3_X1  g468(.A1(new_n607), .A2(new_n643), .A3(new_n630), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n371), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n673));
  OR3_X1    g472(.A1(new_n672), .A2(G29gat), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n561), .A2(new_n597), .A3(new_n664), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n606), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n676), .A2(new_n630), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n629), .B1(new_n598), .B2(new_n606), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n310), .B(KEYINPUT105), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n643), .A2(new_n254), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n683), .B(KEYINPUT106), .Z(new_n684));
  NAND2_X1  g483(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(G29gat), .B1(new_n685), .B2(new_n595), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n673), .B1(new_n672), .B2(G29gat), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n674), .A2(new_n686), .A3(new_n687), .ZN(G1328gat));
  INV_X1    g487(.A(new_n520), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n689), .A2(G36gat), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n671), .A2(new_n690), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n691), .A2(KEYINPUT46), .ZN(new_n692));
  OAI21_X1  g491(.A(G36gat), .B1(new_n685), .B2(new_n689), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(KEYINPUT46), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(G1329gat));
  INV_X1    g494(.A(KEYINPUT108), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT47), .ZN(new_n697));
  OAI21_X1  g496(.A(G43gat), .B1(new_n685), .B2(new_n664), .ZN(new_n698));
  INV_X1    g497(.A(G43gat), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n671), .A2(new_n699), .A3(new_n601), .ZN(new_n700));
  AOI211_X1 g499(.A(new_n696), .B(new_n697), .C1(new_n698), .C2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n696), .A2(new_n697), .ZN(new_n703));
  AND4_X1   g502(.A1(new_n702), .A2(new_n698), .A3(new_n703), .A4(new_n700), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n701), .A2(new_n704), .ZN(G1330gat));
  NOR2_X1   g504(.A1(new_n670), .A2(new_n560), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n681), .A2(G50gat), .A3(new_n684), .ZN(new_n707));
  OAI22_X1  g506(.A1(new_n706), .A2(G50gat), .B1(new_n560), .B2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g508(.A1(new_n625), .A2(KEYINPUT97), .A3(new_n626), .ZN(new_n710));
  INV_X1    g509(.A(new_n610), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n712), .A2(new_n642), .A3(new_n627), .A4(new_n255), .ZN(new_n713));
  AOI211_X1 g512(.A(new_n682), .B(new_n713), .C1(new_n675), .C2(new_n606), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n371), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(new_n281), .ZN(G1332gat));
  INV_X1    g515(.A(KEYINPUT49), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n520), .B1(new_n717), .B2(new_n277), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT109), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT110), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1333gat));
  INV_X1    g525(.A(new_n664), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n714), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(G71gat), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n601), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n729), .B1(G71gat), .B2(new_n730), .ZN(new_n731));
  XOR2_X1   g530(.A(new_n731), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g531(.A1(new_n714), .A2(new_n559), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g533(.A(new_n629), .B1(new_n675), .B2(new_n606), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n642), .A2(new_n254), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT51), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(KEYINPUT51), .B1(new_n735), .B2(new_n736), .ZN(new_n740));
  OR2_X1    g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n371), .A2(new_n259), .A3(new_n310), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT113), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT112), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n736), .A2(new_n310), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT111), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n745), .B1(new_n681), .B2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n680), .A2(new_n679), .ZN(new_n750));
  INV_X1    g549(.A(new_n677), .ZN(new_n751));
  AOI211_X1 g550(.A(new_n629), .B(new_n751), .C1(new_n675), .C2(new_n606), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n745), .B(new_n747), .C1(new_n750), .C2(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n595), .B1(new_n749), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n744), .B1(new_n754), .B2(new_n259), .ZN(G1336gat));
  INV_X1    g554(.A(KEYINPUT114), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n737), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n738), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n737), .A2(new_n756), .A3(KEYINPUT51), .ZN(new_n759));
  OR3_X1    g558(.A1(new_n689), .A2(G92gat), .A3(new_n682), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  AND3_X1   g560(.A1(new_n758), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n753), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n520), .B1(new_n763), .B2(new_n748), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n762), .B1(new_n764), .B2(G92gat), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n520), .B(new_n747), .C1(new_n750), .C2(new_n752), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT52), .B1(new_n767), .B2(G92gat), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n761), .B1(new_n739), .B2(new_n740), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT115), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AND3_X1   g569(.A1(new_n768), .A2(KEYINPUT115), .A3(new_n769), .ZN(new_n771));
  OAI22_X1  g570(.A1(new_n765), .A2(new_n766), .B1(new_n770), .B2(new_n771), .ZN(G1337gat));
  INV_X1    g571(.A(G99gat), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n601), .A2(new_n773), .A3(new_n310), .ZN(new_n774));
  XOR2_X1   g573(.A(new_n774), .B(KEYINPUT116), .Z(new_n775));
  NAND2_X1  g574(.A1(new_n741), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n664), .B1(new_n749), .B2(new_n753), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n776), .B1(new_n777), .B2(new_n773), .ZN(G1338gat));
  NOR3_X1   g577(.A1(new_n560), .A2(G106gat), .A3(new_n682), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n758), .A2(new_n759), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n559), .B1(new_n763), .B2(new_n748), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n780), .B1(new_n781), .B2(G106gat), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n559), .B(new_n747), .C1(new_n750), .C2(new_n752), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT53), .B1(new_n784), .B2(G106gat), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n779), .B1(new_n739), .B2(new_n740), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT117), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n785), .A2(KEYINPUT117), .A3(new_n786), .ZN(new_n788));
  OAI22_X1  g587(.A1(new_n782), .A2(new_n783), .B1(new_n787), .B2(new_n788), .ZN(G1339gat));
  INV_X1    g588(.A(KEYINPUT120), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n713), .A2(new_n310), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT119), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n229), .B1(new_n228), .B2(new_n231), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n234), .A2(new_n235), .A3(new_n233), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n241), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT118), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI211_X1 g596(.A(KEYINPUT118), .B(new_n241), .C1(new_n793), .C2(new_n794), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n799), .A2(new_n251), .A3(new_n310), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n295), .A2(new_n258), .A3(new_n296), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n298), .A2(KEYINPUT54), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n308), .B1(new_n297), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n802), .A2(KEYINPUT55), .A3(new_n804), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(new_n309), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n809), .B1(new_n251), .B2(new_n253), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n792), .B1(new_n800), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n809), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n254), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n799), .A2(new_n251), .A3(new_n310), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n813), .A2(KEYINPUT119), .A3(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n811), .A2(new_n627), .A3(new_n712), .A4(new_n815), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n799), .A2(new_n251), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n817), .B(new_n812), .C1(new_n623), .C2(new_n628), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n791), .B1(new_n819), .B2(new_n643), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n790), .B1(new_n820), .B2(new_n559), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n642), .B1(new_n816), .B2(new_n818), .ZN(new_n822));
  OAI211_X1 g621(.A(KEYINPUT120), .B(new_n560), .C1(new_n822), .C2(new_n791), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n824), .A2(new_n601), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n520), .A2(new_n595), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(G113gat), .B1(new_n827), .B2(new_n255), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n819), .A2(new_n643), .ZN(new_n829));
  INV_X1    g628(.A(new_n791), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n604), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n831), .A2(new_n832), .A3(new_n826), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT121), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(new_n315), .A3(new_n254), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n828), .A2(new_n835), .ZN(G1340gat));
  OAI21_X1  g635(.A(G120gat), .B1(new_n827), .B2(new_n682), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n834), .A2(new_n317), .A3(new_n310), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(G1341gat));
  NAND4_X1  g638(.A1(new_n824), .A2(new_n642), .A3(new_n601), .A4(new_n826), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(G127gat), .ZN(new_n841));
  OR3_X1    g640(.A1(new_n833), .A2(G127gat), .A3(new_n643), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(KEYINPUT122), .ZN(G1342gat));
  OAI21_X1  g643(.A(G134gat), .B1(new_n827), .B2(new_n629), .ZN(new_n845));
  OR3_X1    g644(.A1(new_n833), .A2(G134gat), .A3(new_n629), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT56), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(KEYINPUT123), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n847), .A2(KEYINPUT123), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n846), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n845), .B(new_n850), .C1(new_n848), .C2(new_n846), .ZN(G1343gat));
  OAI211_X1 g650(.A(new_n712), .B(new_n627), .C1(new_n800), .C2(new_n810), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n642), .B1(new_n818), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n559), .B1(new_n853), .B2(new_n791), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT57), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n727), .A2(new_n595), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n857), .A2(new_n520), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n831), .A2(new_n559), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n855), .B(new_n858), .C1(new_n859), .C2(KEYINPUT57), .ZN(new_n860));
  OAI21_X1  g659(.A(G141gat), .B1(new_n860), .B2(new_n255), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT58), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n859), .A2(KEYINPUT124), .A3(new_n857), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT124), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n820), .A2(new_n560), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n864), .B1(new_n865), .B2(new_n856), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n689), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n255), .A2(G141gat), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n861), .B(new_n862), .C1(new_n867), .C2(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n865), .A2(new_n858), .A3(new_n868), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n861), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n870), .B1(new_n872), .B2(new_n862), .ZN(G1344gat));
  INV_X1    g672(.A(KEYINPUT59), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT57), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n854), .A2(KEYINPUT57), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(new_n310), .A3(new_n858), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n874), .B1(new_n878), .B2(G148gat), .ZN(new_n879));
  INV_X1    g678(.A(new_n310), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n874), .B1(new_n860), .B2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(G148gat), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n310), .A2(new_n882), .ZN(new_n884));
  OAI22_X1  g683(.A1(new_n879), .A2(new_n883), .B1(new_n867), .B2(new_n884), .ZN(G1345gat));
  NOR3_X1   g684(.A1(new_n860), .A2(new_n327), .A3(new_n643), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n867), .A2(new_n643), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(new_n327), .ZN(G1346gat));
  NOR3_X1   g687(.A1(new_n860), .A2(new_n328), .A3(new_n629), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n867), .A2(new_n629), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n889), .B1(new_n890), .B2(new_n328), .ZN(G1347gat));
  NOR2_X1   g690(.A1(new_n689), .A2(new_n371), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n825), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(G169gat), .B1(new_n893), .B2(new_n255), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n832), .B(new_n892), .C1(new_n822), .C2(new_n791), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n896), .A2(new_n392), .A3(new_n254), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n894), .A2(new_n897), .ZN(G1348gat));
  AOI21_X1  g697(.A(G176gat), .B1(new_n896), .B2(new_n310), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n893), .A2(new_n682), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(G176gat), .ZN(G1349gat));
  OR2_X1    g700(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n824), .A2(new_n642), .A3(new_n601), .A4(new_n892), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n409), .ZN(new_n904));
  NAND2_X1  g703(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT125), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n831), .A2(new_n429), .A3(new_n832), .A4(new_n892), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n906), .B1(new_n907), .B2(new_n643), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n896), .A2(KEYINPUT125), .A3(new_n642), .A4(new_n429), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AND4_X1   g709(.A1(new_n902), .A2(new_n904), .A3(new_n905), .A4(new_n910), .ZN(new_n911));
  AOI22_X1  g710(.A1(new_n903), .A2(new_n409), .B1(new_n908), .B2(new_n909), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n902), .B1(new_n912), .B2(new_n905), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n911), .A2(new_n913), .ZN(G1350gat));
  NAND3_X1  g713(.A1(new_n896), .A2(new_n630), .A3(new_n422), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n824), .A2(new_n630), .A3(new_n601), .A4(new_n892), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT61), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n916), .A2(new_n917), .A3(G190gat), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(new_n916), .B2(G190gat), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n915), .B1(new_n918), .B2(new_n919), .ZN(G1351gat));
  AND2_X1   g719(.A1(new_n664), .A2(new_n892), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n877), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(G197gat), .B1(new_n922), .B2(new_n255), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n865), .A2(new_n921), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n924), .A2(G197gat), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n923), .B1(new_n255), .B2(new_n925), .ZN(G1352gat));
  OAI21_X1  g725(.A(G204gat), .B1(new_n922), .B2(new_n682), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n924), .A2(G204gat), .A3(new_n880), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT62), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n929), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n927), .A2(new_n930), .A3(new_n931), .ZN(G1353gat));
  NAND4_X1  g731(.A1(new_n875), .A2(new_n876), .A3(new_n642), .A4(new_n921), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(G211gat), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT127), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n934), .A2(new_n935), .A3(KEYINPUT63), .ZN(new_n936));
  INV_X1    g735(.A(new_n924), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n937), .A2(new_n376), .A3(new_n642), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n935), .A2(KEYINPUT63), .ZN(new_n939));
  OR2_X1    g738(.A1(new_n935), .A2(KEYINPUT63), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n933), .A2(G211gat), .A3(new_n939), .A4(new_n940), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n936), .A2(new_n938), .A3(new_n941), .ZN(G1354gat));
  OAI21_X1  g741(.A(G218gat), .B1(new_n922), .B2(new_n629), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n937), .A2(new_n377), .A3(new_n630), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1355gat));
endmodule


