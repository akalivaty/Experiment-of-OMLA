//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1 0 0 0 1 1 1 0 1 1 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT32), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT69), .ZN(new_n191));
  NOR2_X1   g005(.A1(G237), .A2(G953), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G210), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n193), .B(KEYINPUT27), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT26), .B(G101), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n194), .B(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT11), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(G137), .ZN(new_n198));
  AND2_X1   g012(.A1(KEYINPUT65), .A2(G134), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT65), .A2(G134), .ZN(new_n200));
  NOR3_X1   g014(.A1(new_n198), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G137), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT11), .A3(G134), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n197), .A2(G137), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g019(.A(G131), .B1(new_n201), .B2(new_n205), .ZN(new_n206));
  OR2_X1    g020(.A1(KEYINPUT65), .A2(G134), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n202), .A2(KEYINPUT11), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT65), .A2(G134), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G131), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n210), .A2(new_n211), .A3(new_n203), .A4(new_n204), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n206), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT64), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G143), .ZN(new_n216));
  INV_X1    g030(.A(G143), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G146), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(KEYINPUT0), .A2(G128), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n214), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(G143), .B(G146), .ZN(new_n222));
  AND2_X1   g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(KEYINPUT64), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(KEYINPUT0), .A2(G128), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  AOI22_X1  g040(.A1(new_n221), .A2(new_n224), .B1(new_n219), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n213), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n229));
  INV_X1    g043(.A(G116), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n229), .B1(new_n230), .B2(G119), .ZN(new_n231));
  INV_X1    g045(.A(G119), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(KEYINPUT67), .A3(G116), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n231), .B(new_n233), .C1(G116), .C2(new_n232), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT2), .B(G113), .ZN(new_n235));
  XOR2_X1   g049(.A(new_n234), .B(new_n235), .Z(new_n236));
  XNOR2_X1  g050(.A(KEYINPUT66), .B(G128), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT1), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n238), .B1(G143), .B2(new_n215), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n219), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n216), .A2(new_n218), .A3(new_n238), .A4(G128), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n211), .B1(G134), .B2(G137), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n207), .A2(new_n209), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n243), .B1(new_n244), .B2(G137), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n212), .A3(new_n245), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n228), .A2(new_n236), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n236), .B1(new_n228), .B2(new_n246), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT28), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n228), .A2(new_n236), .A3(new_n246), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT28), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n196), .B1(new_n249), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n228), .A2(new_n246), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT30), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n236), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n212), .A2(new_n245), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n242), .A2(new_n258), .B1(new_n213), .B2(new_n227), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n257), .B1(new_n259), .B2(KEYINPUT30), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n228), .A2(new_n257), .A3(KEYINPUT30), .A4(new_n246), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n256), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n250), .A2(new_n196), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n253), .B1(new_n266), .B2(KEYINPUT31), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n228), .A2(KEYINPUT30), .A3(new_n246), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT68), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n261), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n264), .B1(new_n270), .B2(new_n256), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT31), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n191), .B1(new_n267), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n196), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n234), .B(new_n235), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n219), .A2(new_n226), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT64), .B1(new_n222), .B2(new_n223), .ZN(new_n278));
  AND4_X1   g092(.A1(KEYINPUT64), .A2(new_n216), .A3(new_n218), .A4(new_n223), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n280), .B1(new_n206), .B2(new_n212), .ZN(new_n281));
  INV_X1    g095(.A(new_n246), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n276), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n251), .B1(new_n283), .B2(new_n250), .ZN(new_n284));
  INV_X1    g098(.A(new_n252), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n275), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n286), .B1(new_n271), .B2(new_n272), .ZN(new_n287));
  AOI211_X1 g101(.A(KEYINPUT31), .B(new_n264), .C1(new_n270), .C2(new_n256), .ZN(new_n288));
  NOR3_X1   g102(.A1(new_n287), .A2(KEYINPUT69), .A3(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n190), .B1(new_n274), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT29), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n249), .A2(new_n196), .A3(new_n252), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n247), .B1(new_n270), .B2(new_n256), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n291), .B(new_n292), .C1(new_n293), .C2(new_n196), .ZN(new_n294));
  INV_X1    g108(.A(G902), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n294), .B(new_n295), .C1(new_n291), .C2(new_n292), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G472), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT69), .B1(new_n287), .B2(new_n288), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n266), .A2(KEYINPUT31), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n299), .A2(new_n191), .A3(new_n273), .A4(new_n286), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n188), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n290), .B(new_n297), .C1(KEYINPUT32), .C2(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT9), .B(G234), .ZN(new_n303));
  OAI21_X1  g117(.A(G221), .B1(new_n303), .B2(G902), .ZN(new_n304));
  INV_X1    g118(.A(G469), .ZN(new_n305));
  XNOR2_X1  g119(.A(G110), .B(G140), .ZN(new_n306));
  INV_X1    g120(.A(G953), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n307), .A2(G227), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n306), .B(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G101), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT3), .ZN(new_n312));
  INV_X1    g126(.A(G107), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n312), .B1(G104), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n312), .A2(G104), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n315), .B1(new_n316), .B2(KEYINPUT77), .ZN(new_n317));
  NAND2_X1  g131(.A1(KEYINPUT78), .A2(G107), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(KEYINPUT78), .A2(G107), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n314), .B1(new_n317), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G104), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G107), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n311), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT77), .B1(new_n323), .B2(KEYINPUT3), .ZN(new_n326));
  OR2_X1    g140(.A1(KEYINPUT78), .A2(G107), .ZN(new_n327));
  OR2_X1    g141(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n326), .A2(new_n327), .A3(new_n328), .A4(new_n318), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n311), .A2(KEYINPUT79), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT79), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G101), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n330), .A2(new_n332), .A3(new_n324), .ZN(new_n333));
  INV_X1    g147(.A(new_n314), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n329), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT4), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n325), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n329), .A2(new_n334), .A3(new_n324), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT4), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n339), .A3(G101), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n227), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(G104), .B1(new_n327), .B2(new_n318), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n313), .A2(G104), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(G101), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G128), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n347), .B1(new_n216), .B2(KEYINPUT1), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n241), .B1(new_n348), .B2(new_n222), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n335), .A2(new_n346), .A3(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT10), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n242), .A2(new_n335), .A3(KEYINPUT10), .A4(new_n346), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(KEYINPUT81), .B1(new_n342), .B2(new_n354), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n227), .B(new_n340), .C1(new_n325), .C2(new_n336), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT81), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n356), .A2(new_n357), .A3(new_n352), .A4(new_n353), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n355), .A2(new_n213), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n213), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n356), .A2(new_n360), .A3(new_n352), .A4(new_n353), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n310), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n310), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n242), .B1(new_n335), .B2(new_n346), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT80), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n360), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n335), .A2(new_n346), .ZN(new_n367));
  OAI211_X1 g181(.A(KEYINPUT80), .B(new_n350), .C1(new_n367), .C2(new_n242), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n366), .A2(KEYINPUT12), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(KEYINPUT12), .B1(new_n366), .B2(new_n368), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n363), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n305), .B(new_n295), .C1(new_n362), .C2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n361), .B1(new_n369), .B2(new_n371), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n309), .ZN(new_n377));
  INV_X1    g191(.A(new_n363), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n359), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(G469), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(G469), .A2(G902), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n304), .B1(new_n375), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(G214), .B1(G237), .B2(G902), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n276), .B(new_n340), .C1(new_n325), .C2(new_n336), .ZN(new_n385));
  OR2_X1    g199(.A1(new_n234), .A2(new_n235), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT5), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(new_n232), .A3(G116), .ZN(new_n388));
  OAI211_X1 g202(.A(G113), .B(new_n388), .C1(new_n234), .C2(new_n387), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n367), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n385), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT82), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT6), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n385), .A2(new_n390), .A3(KEYINPUT82), .ZN(new_n395));
  XNOR2_X1  g209(.A(G110), .B(G122), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n393), .A2(new_n394), .A3(new_n395), .A4(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G125), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n242), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n400), .B1(new_n399), .B2(new_n280), .ZN(new_n401));
  XNOR2_X1  g215(.A(KEYINPUT83), .B(G224), .ZN(new_n402));
  OR2_X1    g216(.A1(new_n402), .A2(G953), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n401), .B(new_n403), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n385), .A2(KEYINPUT82), .A3(new_n390), .ZN(new_n405));
  AOI21_X1  g219(.A(KEYINPUT82), .B1(new_n385), .B2(new_n390), .ZN(new_n406));
  NOR3_X1   g220(.A1(new_n405), .A2(new_n406), .A3(new_n396), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n385), .A2(new_n390), .A3(new_n396), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT6), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n398), .B(new_n404), .C1(new_n407), .C2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n403), .A2(KEYINPUT7), .ZN(new_n411));
  INV_X1    g225(.A(new_n401), .ZN(new_n412));
  AND2_X1   g226(.A1(KEYINPUT85), .A2(KEYINPUT7), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT85), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n401), .A2(new_n415), .A3(KEYINPUT7), .A4(new_n403), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n414), .A2(new_n416), .A3(new_n408), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n396), .B(KEYINPUT8), .ZN(new_n418));
  AND4_X1   g232(.A1(new_n386), .A2(new_n389), .A3(new_n335), .A4(new_n346), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n389), .A2(new_n386), .B1(new_n335), .B2(new_n346), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT84), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT84), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n423), .B(new_n418), .C1(new_n419), .C2(new_n420), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(G902), .B1(new_n417), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(G210), .B1(G237), .B2(G902), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n410), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n427), .B1(new_n410), .B2(new_n426), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n384), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n383), .A2(new_n430), .ZN(new_n431));
  XOR2_X1   g245(.A(KEYINPUT70), .B(G217), .Z(new_n432));
  AOI21_X1  g246(.A(new_n432), .B1(G234), .B2(new_n295), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n347), .A2(KEYINPUT66), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT66), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(G128), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n435), .A2(new_n437), .A3(KEYINPUT23), .A4(G119), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n232), .A2(G128), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT23), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n440), .B1(new_n232), .B2(G128), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n438), .A2(KEYINPUT71), .A3(new_n439), .A4(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT71), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n237), .A2(new_n443), .A3(KEYINPUT23), .A4(G119), .ZN(new_n444));
  AOI21_X1  g258(.A(G110), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  XOR2_X1   g259(.A(KEYINPUT24), .B(G110), .Z(new_n446));
  NAND2_X1  g260(.A1(new_n237), .A2(G119), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n446), .B1(new_n447), .B2(new_n439), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G140), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G125), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n399), .A2(G140), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n452), .A3(KEYINPUT72), .ZN(new_n453));
  OR3_X1    g267(.A1(new_n450), .A2(KEYINPUT72), .A3(G125), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(new_n454), .A3(KEYINPUT16), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT16), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n451), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G146), .ZN(new_n459));
  XNOR2_X1  g273(.A(G125), .B(G140), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n460), .A2(KEYINPUT74), .A3(new_n215), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT74), .B1(new_n460), .B2(new_n215), .ZN(new_n462));
  OR2_X1    g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  OR2_X1    g278(.A1(new_n449), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n442), .A2(G110), .A3(new_n444), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n447), .A2(new_n439), .A3(new_n446), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n455), .A2(new_n215), .A3(new_n457), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n459), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT73), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n455), .A2(new_n215), .A3(new_n457), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n215), .B1(new_n455), .B2(new_n457), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n466), .A2(new_n467), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT73), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n465), .B1(new_n471), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT75), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n449), .A2(new_n464), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n476), .B1(new_n474), .B2(new_n475), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n468), .A2(new_n470), .A3(KEYINPUT73), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT75), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n307), .A2(G221), .A3(G234), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(KEYINPUT76), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT22), .B(G137), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n487), .B(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n480), .A2(new_n485), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(G902), .B1(new_n484), .B2(new_n489), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n434), .B1(new_n493), .B2(KEYINPUT25), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT25), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n491), .A2(new_n495), .A3(new_n492), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n433), .A2(G902), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n484), .A2(new_n489), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n491), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  AOI22_X1  g314(.A1(new_n494), .A2(new_n496), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT87), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n192), .A2(G143), .A3(G214), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(G143), .B1(new_n192), .B2(G214), .ZN(new_n505));
  OAI21_X1  g319(.A(G131), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n192), .A2(G214), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n217), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(new_n211), .A3(new_n503), .ZN(new_n509));
  AOI22_X1  g323(.A1(new_n458), .A2(G146), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT19), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n511), .B1(new_n453), .B2(new_n454), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n460), .A2(KEYINPUT19), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n215), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(KEYINPUT18), .A2(G131), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n508), .A2(new_n503), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n516), .B1(new_n508), .B2(new_n503), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n453), .A2(new_n454), .A3(G146), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n520), .B1(new_n461), .B2(new_n462), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n515), .A2(new_n522), .ZN(new_n523));
  XOR2_X1   g337(.A(KEYINPUT86), .B(G104), .Z(new_n524));
  XNOR2_X1  g338(.A(G113), .B(G122), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n524), .B(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n502), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT17), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n506), .A2(new_n509), .A3(new_n528), .ZN(new_n529));
  OAI211_X1 g343(.A(KEYINPUT17), .B(G131), .C1(new_n504), .C2(new_n505), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n459), .A2(new_n529), .A3(new_n469), .A4(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n526), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n532), .A3(new_n522), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT20), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n523), .A2(new_n502), .A3(new_n526), .ZN(new_n536));
  NOR2_X1   g350(.A1(G475), .A2(G902), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n534), .A2(new_n535), .A3(new_n536), .A4(new_n537), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n510), .A2(new_n514), .B1(new_n521), .B2(new_n519), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT87), .B1(new_n539), .B2(new_n532), .ZN(new_n540));
  INV_X1    g354(.A(new_n533), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n536), .B(new_n537), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT20), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n538), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n531), .A2(new_n522), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n526), .ZN(new_n546));
  AOI21_X1  g360(.A(G902), .B1(new_n546), .B2(new_n533), .ZN(new_n547));
  XOR2_X1   g361(.A(KEYINPUT88), .B(G475), .Z(new_n548));
  NOR2_X1   g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n544), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(G116), .B(G122), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n321), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n321), .A2(new_n552), .ZN(new_n555));
  OR2_X1    g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n435), .A2(new_n437), .A3(G143), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n199), .A2(new_n200), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n217), .A2(G128), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT89), .B(KEYINPUT13), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n557), .B1(new_n561), .B2(new_n559), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT13), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT89), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT89), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT13), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n559), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT90), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n561), .A2(KEYINPUT90), .A3(new_n559), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n562), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(G134), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n556), .B(new_n560), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT91), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n230), .A2(KEYINPUT14), .A3(G122), .ZN(new_n575));
  INV_X1    g389(.A(new_n552), .ZN(new_n576));
  OAI211_X1 g390(.A(G107), .B(new_n575), .C1(new_n576), .C2(KEYINPUT14), .ZN(new_n577));
  INV_X1    g391(.A(new_n560), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n558), .B1(new_n557), .B2(new_n559), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n577), .B(new_n553), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  NOR3_X1   g394(.A1(new_n432), .A2(G953), .A3(new_n303), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n573), .A2(new_n574), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n562), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n569), .A2(new_n570), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n572), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n560), .B1(new_n554), .B2(new_n555), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n580), .B(new_n581), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT91), .ZN(new_n588));
  INV_X1    g402(.A(new_n581), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n585), .A2(new_n586), .ZN(new_n590));
  INV_X1    g404(.A(new_n580), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n582), .A2(new_n588), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n295), .ZN(new_n594));
  INV_X1    g408(.A(G478), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(KEYINPUT15), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(G234), .A2(G237), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(G952), .A3(new_n307), .ZN(new_n599));
  OR2_X1    g413(.A1(new_n599), .A2(KEYINPUT92), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(KEYINPUT92), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT21), .B(G898), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n598), .A2(G902), .A3(G953), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n593), .B(new_n295), .C1(KEYINPUT15), .C2(new_n595), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n597), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(KEYINPUT93), .B1(new_n551), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n597), .A2(new_n607), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n549), .B1(new_n538), .B2(new_n543), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT93), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n611), .A2(new_n612), .A3(new_n613), .A4(new_n606), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n302), .A2(new_n431), .A3(new_n501), .A4(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n330), .A2(new_n332), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G3));
  INV_X1    g432(.A(new_n304), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n376), .A2(new_n309), .B1(new_n359), .B2(new_n378), .ZN(new_n620));
  OAI21_X1  g434(.A(G469), .B1(new_n620), .B2(G902), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n619), .B1(new_n621), .B2(new_n374), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n493), .A2(KEYINPUT25), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n623), .A2(new_n433), .A3(new_n496), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n500), .A2(new_n497), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n622), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n298), .A2(new_n300), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n295), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n301), .B1(new_n628), .B2(G472), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n606), .B(new_n384), .C1(new_n428), .C2(new_n429), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT33), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n593), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(KEYINPUT94), .B1(new_n590), .B2(new_n591), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n581), .ZN(new_n635));
  OAI211_X1 g449(.A(KEYINPUT94), .B(new_n589), .C1(new_n590), .C2(new_n591), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n635), .A2(KEYINPUT33), .A3(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n633), .A2(new_n637), .A3(G478), .A4(new_n295), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n594), .A2(new_n595), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n551), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n631), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n630), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT34), .B(G104), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G6));
  NAND3_X1  g459(.A1(new_n538), .A2(new_n543), .A3(KEYINPUT95), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT95), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n542), .A2(new_n647), .A3(KEYINPUT20), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n646), .A2(new_n550), .A3(new_n610), .A4(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n631), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n630), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT35), .B(G107), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  NOR2_X1   g467(.A1(new_n490), .A2(KEYINPUT36), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n478), .A2(new_n479), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n484), .A2(KEYINPUT75), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n654), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n480), .A2(new_n485), .A3(new_n658), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n657), .A2(new_n497), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(new_n494), .B2(new_n496), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n629), .A2(new_n431), .A3(new_n615), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT96), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT37), .B(G110), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G12));
  NAND2_X1  g480(.A1(new_n627), .A2(new_n187), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n189), .ZN(new_n668));
  AOI22_X1  g482(.A1(new_n627), .A2(new_n190), .B1(G472), .B2(new_n296), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n661), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT97), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n646), .A2(new_n610), .A3(new_n648), .ZN(new_n672));
  INV_X1    g486(.A(G900), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n602), .B1(new_n673), .B2(new_n604), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n550), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n671), .B1(new_n678), .B2(new_n430), .ZN(new_n679));
  INV_X1    g493(.A(new_n430), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n680), .A2(KEYINPUT97), .A3(new_n677), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n670), .A2(new_n679), .A3(new_n622), .A4(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT98), .B(G128), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G30));
  NOR2_X1   g498(.A1(new_n293), .A2(new_n275), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n247), .A2(new_n248), .ZN(new_n686));
  AOI21_X1  g500(.A(G902), .B1(new_n686), .B2(new_n275), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g502(.A(G472), .B1(new_n685), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n668), .A2(new_n290), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n410), .A2(new_n426), .ZN(new_n691));
  INV_X1    g505(.A(new_n427), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n410), .A2(new_n426), .A3(new_n427), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n384), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n611), .A2(new_n612), .A3(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n690), .A2(new_n697), .A3(new_n661), .A4(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT100), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT101), .B(KEYINPUT39), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n674), .B(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n622), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n706), .B(KEYINPUT40), .Z(new_n707));
  NAND3_X1  g521(.A1(new_n702), .A2(new_n703), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(KEYINPUT102), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT102), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n702), .A2(new_n710), .A3(new_n703), .A4(new_n707), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(new_n217), .ZN(G45));
  NAND3_X1  g527(.A1(new_n551), .A2(new_n640), .A3(new_n675), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n670), .A2(new_n680), .A3(new_n622), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G146), .ZN(G48));
  OAI21_X1  g531(.A(new_n295), .B1(new_n362), .B2(new_n373), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(G469), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n304), .A3(new_n374), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n302), .A2(new_n642), .A3(new_n501), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT41), .B(G113), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G15));
  NAND4_X1  g538(.A1(new_n302), .A2(new_n650), .A3(new_n501), .A4(new_n721), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G116), .ZN(G18));
  NOR2_X1   g540(.A1(new_n720), .A2(new_n430), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n302), .A2(new_n615), .A3(new_n727), .A4(new_n662), .ZN(new_n728));
  XNOR2_X1  g542(.A(KEYINPUT103), .B(G119), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(G21));
  AOI21_X1  g544(.A(new_n272), .B1(new_n263), .B2(new_n265), .ZN(new_n731));
  OAI21_X1  g545(.A(KEYINPUT104), .B1(new_n731), .B2(new_n253), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT104), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n286), .B(new_n733), .C1(new_n271), .C2(new_n272), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n732), .A2(new_n273), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n187), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT105), .ZN(new_n737));
  AOI22_X1  g551(.A1(new_n628), .A2(G472), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n719), .A2(new_n606), .A3(new_n304), .A4(new_n374), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n698), .B1(new_n597), .B2(new_n607), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n551), .B(new_n740), .C1(new_n428), .C2(new_n429), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n735), .A2(KEYINPUT105), .A3(new_n187), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n738), .A2(new_n742), .A3(new_n501), .A4(new_n743), .ZN(new_n744));
  XOR2_X1   g558(.A(KEYINPUT106), .B(G122), .Z(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G24));
  NOR3_X1   g560(.A1(new_n720), .A2(new_n430), .A3(new_n714), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n747), .A2(new_n738), .A3(new_n662), .A4(new_n743), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G125), .ZN(G27));
  INV_X1    g563(.A(KEYINPUT42), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n290), .A2(new_n297), .ZN(new_n751));
  AOI21_X1  g565(.A(KEYINPUT32), .B1(new_n627), .B2(new_n187), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n501), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n693), .A2(new_n384), .A3(new_n694), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(new_n715), .A3(new_n622), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n750), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n624), .A2(new_n625), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n758), .B1(new_n668), .B2(new_n669), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n383), .A2(new_n754), .A3(new_n714), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(KEYINPUT42), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n757), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G131), .ZN(G33));
  NOR2_X1   g577(.A1(new_n383), .A2(new_n754), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n302), .A2(new_n764), .A3(new_n501), .A4(new_n677), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G134), .ZN(G36));
  OR2_X1    g580(.A1(new_n620), .A2(KEYINPUT45), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n620), .A2(KEYINPUT45), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(G469), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT46), .B1(new_n769), .B2(new_n381), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n770), .A2(new_n375), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n769), .A2(KEYINPUT46), .A3(new_n381), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n619), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n705), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT107), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n612), .A2(new_n640), .ZN(new_n776));
  XOR2_X1   g590(.A(new_n776), .B(KEYINPUT43), .Z(new_n777));
  INV_X1    g591(.A(G472), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n778), .B1(new_n627), .B2(new_n295), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n777), .B(new_n662), .C1(new_n301), .C2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n754), .B1(new_n781), .B2(KEYINPUT44), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n782), .B1(KEYINPUT44), .B2(new_n781), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n775), .A2(new_n783), .ZN(new_n784));
  XOR2_X1   g598(.A(KEYINPUT108), .B(G137), .Z(new_n785));
  XNOR2_X1  g599(.A(new_n784), .B(new_n785), .ZN(G39));
  XNOR2_X1  g600(.A(new_n773), .B(KEYINPUT47), .ZN(new_n787));
  NOR4_X1   g601(.A1(new_n302), .A2(new_n501), .A3(new_n714), .A4(new_n754), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT109), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n787), .A2(KEYINPUT109), .A3(new_n788), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G140), .ZN(G42));
  AND2_X1   g608(.A1(new_n738), .A2(new_n743), .ZN(new_n795));
  AND4_X1   g609(.A1(new_n501), .A2(new_n795), .A3(new_n602), .A4(new_n777), .ZN(new_n796));
  INV_X1    g610(.A(new_n697), .ZN(new_n797));
  OAI21_X1  g611(.A(KEYINPUT116), .B1(new_n720), .B2(new_n384), .ZN(new_n798));
  OR3_X1    g612(.A1(new_n720), .A2(KEYINPUT116), .A3(new_n384), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT117), .B1(new_n796), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT50), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n795), .A2(new_n662), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  AND4_X1   g619(.A1(new_n602), .A2(new_n777), .A3(new_n721), .A4(new_n755), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n501), .A2(new_n602), .ZN(new_n807));
  NOR4_X1   g621(.A1(new_n690), .A2(new_n720), .A3(new_n807), .A4(new_n754), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n551), .A2(new_n640), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n805), .A2(new_n806), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n803), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n802), .A2(KEYINPUT50), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n719), .A2(new_n374), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(new_n304), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n755), .B(new_n796), .C1(new_n787), .C2(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT51), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n806), .A2(new_n759), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(KEYINPUT48), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n796), .A2(new_n727), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n307), .A2(G952), .ZN(new_n821));
  AOI22_X1  g635(.A1(new_n544), .A2(new_n550), .B1(new_n638), .B2(new_n639), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n821), .B1(new_n808), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n819), .A2(new_n820), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n817), .A2(new_n824), .ZN(new_n825));
  OR3_X1    g639(.A1(new_n811), .A2(KEYINPUT118), .A3(new_n812), .ZN(new_n826));
  OAI21_X1  g640(.A(KEYINPUT118), .B1(new_n811), .B2(new_n812), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n826), .A2(KEYINPUT51), .A3(new_n827), .A4(new_n816), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT112), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n615), .A2(new_n680), .A3(new_n622), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n779), .A2(new_n661), .A3(new_n301), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n830), .B1(new_n759), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n612), .A2(new_n610), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n833), .A2(new_n822), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n834), .A2(new_n631), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n835), .A2(new_n626), .A3(new_n629), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT111), .B1(new_n832), .B2(new_n836), .ZN(new_n837));
  AND4_X1   g651(.A1(KEYINPUT111), .A2(new_n616), .A3(new_n663), .A4(new_n836), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n760), .A2(new_n738), .A3(new_n662), .A4(new_n743), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n646), .A2(new_n648), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n841), .A2(new_n610), .A3(new_n676), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n302), .A2(new_n764), .A3(new_n662), .A4(new_n842), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n840), .A2(new_n765), .A3(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n722), .A2(new_n725), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n744), .A2(new_n728), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n844), .A2(new_n762), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n829), .B1(new_n839), .B2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT111), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n616), .A2(new_n663), .ZN(new_n850));
  INV_X1    g664(.A(new_n836), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n832), .A2(KEYINPUT111), .A3(new_n836), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n846), .A2(new_n845), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n840), .A2(new_n765), .A3(new_n843), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n856), .B1(new_n757), .B2(new_n761), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n854), .A2(new_n855), .A3(new_n857), .A4(KEYINPUT112), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT53), .B1(new_n848), .B2(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n716), .A2(new_n748), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n674), .B(KEYINPUT113), .Z(new_n861));
  NOR3_X1   g675(.A1(new_n383), .A2(new_n741), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n690), .A2(new_n862), .A3(new_n661), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n860), .A2(KEYINPUT52), .A3(new_n682), .A4(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n682), .A2(new_n716), .A3(new_n863), .A4(new_n748), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT115), .ZN(new_n866));
  XNOR2_X1  g680(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n866), .B1(new_n865), .B2(new_n867), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n859), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT52), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n865), .A2(new_n875), .ZN(new_n876));
  AOI22_X1  g690(.A1(new_n848), .A2(new_n858), .B1(new_n864), .B2(new_n876), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n873), .B(KEYINPUT54), .C1(new_n874), .C2(new_n877), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n839), .A2(new_n847), .A3(new_n874), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n864), .A2(new_n868), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n879), .B1(new_n870), .B2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT54), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n881), .B(new_n882), .C1(new_n877), .C2(KEYINPUT53), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n825), .A2(new_n828), .A3(new_n878), .A4(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n884), .B1(G952), .B2(G953), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n776), .A2(new_n698), .A3(new_n619), .ZN(new_n886));
  INV_X1    g700(.A(new_n814), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT49), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n886), .B(new_n501), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(KEYINPUT110), .Z(new_n890));
  AOI21_X1  g704(.A(new_n690), .B1(new_n888), .B2(new_n887), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n890), .A2(new_n797), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n885), .A2(new_n892), .ZN(G75));
  OAI21_X1  g707(.A(new_n881), .B1(new_n877), .B2(KEYINPUT53), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n894), .A2(G210), .A3(G902), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n407), .A2(new_n409), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n896), .B1(new_n394), .B2(new_n407), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(new_n404), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT55), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n895), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n900), .B1(new_n895), .B2(new_n901), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n307), .A2(G952), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(G51));
  NAND2_X1  g719(.A1(new_n894), .A2(KEYINPUT54), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n883), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n381), .B(KEYINPUT57), .ZN(new_n909));
  OAI22_X1  g723(.A1(new_n908), .A2(new_n909), .B1(new_n362), .B2(new_n373), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n854), .A2(new_n855), .A3(new_n857), .A4(KEYINPUT53), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n911), .B1(new_n869), .B2(new_n871), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n848), .A2(new_n858), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n864), .A2(new_n876), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n912), .B1(new_n915), .B2(new_n874), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n916), .A2(new_n295), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n769), .B(KEYINPUT120), .Z(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n904), .B1(new_n910), .B2(new_n919), .ZN(G54));
  INV_X1    g734(.A(new_n536), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n527), .B2(new_n533), .ZN(new_n922));
  NAND2_X1  g736(.A1(KEYINPUT58), .A2(G475), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT121), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n917), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n922), .B1(new_n917), .B2(new_n924), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n925), .A2(new_n926), .A3(new_n904), .ZN(G60));
  INV_X1    g741(.A(new_n904), .ZN(new_n928));
  NAND2_X1  g742(.A1(G478), .A2(G902), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT59), .Z(new_n930));
  AOI21_X1  g744(.A(new_n930), .B1(new_n878), .B2(new_n883), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n633), .A2(new_n637), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n928), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n932), .A2(new_n930), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(KEYINPUT122), .B1(new_n908), .B2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT122), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n907), .A2(new_n938), .A3(new_n935), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n934), .B1(new_n937), .B2(new_n939), .ZN(G63));
  NAND2_X1  g754(.A1(new_n928), .A2(KEYINPUT61), .ZN(new_n941));
  NAND2_X1  g755(.A1(G217), .A2(G902), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT60), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n499), .B1(new_n916), .B2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT124), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n941), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n657), .A2(new_n659), .ZN(new_n947));
  INV_X1    g761(.A(new_n943), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT53), .B1(new_n913), .B2(new_n914), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n947), .B(new_n948), .C1(new_n949), .C2(new_n912), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT123), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n894), .A2(KEYINPUT123), .A3(new_n947), .A4(new_n948), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n500), .B1(new_n894), .B2(new_n948), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(KEYINPUT124), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n946), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  AOI211_X1 g771(.A(new_n904), .B(new_n955), .C1(new_n952), .C2(new_n953), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n957), .B1(new_n958), .B2(KEYINPUT61), .ZN(G66));
  OAI21_X1  g773(.A(G953), .B1(new_n603), .B2(new_n402), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n854), .A2(new_n855), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n960), .B1(new_n961), .B2(G953), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT125), .Z(new_n963));
  INV_X1    g777(.A(G898), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n897), .B1(new_n964), .B2(G953), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n963), .B(new_n965), .ZN(G69));
  OAI21_X1  g780(.A(new_n270), .B1(KEYINPUT30), .B2(new_n259), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n512), .A2(new_n513), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n969), .B1(new_n673), .B2(new_n307), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n759), .A2(new_n695), .A3(new_n699), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n783), .A2(new_n971), .ZN(new_n972));
  OR2_X1    g786(.A1(new_n972), .A2(new_n775), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n860), .A2(new_n682), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n974), .A2(new_n762), .A3(new_n765), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n973), .A2(new_n793), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n970), .B1(new_n976), .B2(new_n307), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n709), .A2(new_n711), .A3(new_n974), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n978), .A2(KEYINPUT62), .ZN(new_n979));
  OR4_X1    g793(.A1(new_n753), .A2(new_n706), .A3(new_n754), .A4(new_n834), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n775), .B2(new_n783), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n981), .B1(new_n791), .B2(new_n792), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n978), .A2(KEYINPUT62), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n979), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n969), .B1(new_n984), .B2(new_n307), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n307), .B1(G227), .B2(G900), .ZN(new_n986));
  OR3_X1    g800(.A1(new_n977), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n986), .B1(new_n977), .B2(new_n985), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(G72));
  AND4_X1   g803(.A1(new_n961), .A2(new_n979), .A3(new_n982), .A4(new_n983), .ZN(new_n990));
  XNOR2_X1  g804(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n778), .A2(new_n295), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n991), .B(new_n992), .Z(new_n993));
  OAI21_X1  g807(.A(new_n685), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n973), .A2(new_n793), .A3(new_n961), .A4(new_n975), .ZN(new_n995));
  INV_X1    g809(.A(new_n993), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n293), .A2(new_n275), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n904), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n994), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n915), .A2(KEYINPUT53), .ZN(new_n1001));
  NOR3_X1   g815(.A1(new_n998), .A2(new_n685), .A3(new_n993), .ZN(new_n1002));
  AND3_X1   g816(.A1(new_n1001), .A2(new_n873), .A3(new_n1002), .ZN(new_n1003));
  OR2_X1    g817(.A1(new_n1003), .A2(KEYINPUT127), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(KEYINPUT127), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1000), .B1(new_n1004), .B2(new_n1005), .ZN(G57));
endmodule


