//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 0 1 0 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 1 1 0 1 1 1 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n625,
    new_n626, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT67), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n450), .B(new_n451), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND3_X1  g032(.A1(new_n454), .A2(KEYINPUT69), .A3(G567), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT69), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n453), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n457), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(KEYINPUT70), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n466), .B1(new_n467), .B2(G125), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n464), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(G125), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(new_n465), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n469), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  OAI211_X1 g053(.A(G137), .B(new_n469), .C1(new_n471), .C2(new_n472), .ZN(new_n479));
  AND3_X1   g054(.A1(new_n476), .A2(new_n478), .A3(new_n479), .ZN(G160));
  NAND2_X1  g055(.A1(new_n467), .A2(new_n469), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n472), .ZN(new_n483));
  NAND2_X1  g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n469), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI22_X1  g060(.A1(new_n482), .A2(G136), .B1(G124), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(G100), .ZN(new_n487));
  AND3_X1   g062(.A1(new_n487), .A2(new_n469), .A3(KEYINPUT71), .ZN(new_n488));
  AOI21_X1  g063(.A(KEYINPUT71), .B1(new_n487), .B2(new_n469), .ZN(new_n489));
  OAI221_X1 g064(.A(G2104), .B1(G112), .B2(new_n469), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  XOR2_X1   g066(.A(new_n491), .B(KEYINPUT72), .Z(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  OAI211_X1 g068(.A(G126), .B(G2105), .C1(new_n471), .C2(new_n472), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n500), .B1(new_n471), .B2(new_n472), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n467), .A2(new_n503), .A3(new_n500), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n498), .B1(new_n502), .B2(new_n504), .ZN(G164));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G50), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n510), .A2(KEYINPUT73), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n512), .B1(new_n509), .B2(G50), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(new_n506), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n507), .A2(new_n508), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G88), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n516), .A2(new_n517), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n519), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n514), .A2(new_n523), .ZN(G166));
  INV_X1    g099(.A(KEYINPUT75), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT74), .B(G51), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n509), .A2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n521), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n525), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n509), .A2(new_n526), .B1(new_n521), .B2(new_n528), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(KEYINPUT75), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n518), .A2(G89), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n530), .A2(new_n532), .A3(new_n534), .A4(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  AOI22_X1  g112(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n520), .ZN(new_n539));
  XNOR2_X1  g114(.A(KEYINPUT6), .B(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n521), .A2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G52), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n541), .A2(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g120(.A(KEYINPUT76), .B1(new_n539), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n518), .A2(G90), .B1(new_n509), .B2(G52), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT76), .ZN(new_n548));
  OAI211_X1 g123(.A(new_n547), .B(new_n548), .C1(new_n520), .C2(new_n538), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n546), .A2(new_n549), .ZN(G171));
  NAND2_X1  g125(.A1(new_n521), .A2(G56), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G651), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(KEYINPUT77), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT77), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n553), .A2(new_n556), .A3(G651), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n518), .A2(G81), .B1(new_n509), .B2(G43), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n555), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n509), .A2(G53), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n566), .B1(new_n567), .B2(KEYINPUT78), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n567), .A2(KEYINPUT79), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT79), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n566), .A2(KEYINPUT78), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n509), .A2(new_n571), .A3(G53), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n518), .A2(G91), .ZN(new_n574));
  INV_X1    g149(.A(G65), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(new_n516), .B2(new_n517), .ZN(new_n576));
  AND2_X1   g151(.A1(G78), .A2(G543), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n573), .A2(new_n574), .A3(new_n578), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n570), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G299));
  INV_X1    g156(.A(G171), .ZN(G301));
  OAI221_X1 g157(.A(new_n519), .B1(new_n520), .B2(new_n522), .C1(new_n511), .C2(new_n513), .ZN(G303));
  NAND2_X1  g158(.A1(new_n518), .A2(G87), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n509), .A2(G49), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(G288));
  AOI22_X1  g162(.A1(new_n518), .A2(G86), .B1(new_n509), .B2(G48), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(new_n516), .B2(new_n517), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(KEYINPUT80), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n593), .A2(G73), .A3(G543), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(G651), .B1(new_n590), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n588), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n597), .B(new_n598), .ZN(G305));
  AOI22_X1  g174(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(new_n520), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  INV_X1    g177(.A(G47), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n541), .A2(new_n602), .B1(new_n543), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(G290));
  INV_X1    g181(.A(G92), .ZN(new_n607));
  OAI21_X1  g182(.A(KEYINPUT82), .B1(new_n541), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT82), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n518), .A2(new_n609), .A3(G92), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n608), .A2(KEYINPUT10), .A3(new_n610), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n521), .A2(G66), .ZN(new_n615));
  INV_X1    g190(.A(G79), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(new_n506), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n617), .A2(G651), .B1(G54), .B2(new_n509), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n613), .A2(new_n614), .A3(new_n618), .ZN(new_n619));
  MUX2_X1   g194(.A(new_n619), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g195(.A(new_n619), .B(G301), .S(G868), .Z(G321));
  NAND2_X1  g196(.A1(G286), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n580), .ZN(G297));
  OAI21_X1  g198(.A(new_n622), .B1(G868), .B2(new_n580), .ZN(G280));
  AND3_X1   g199(.A1(new_n613), .A2(new_n614), .A3(new_n618), .ZN(new_n625));
  XOR2_X1   g200(.A(KEYINPUT83), .B(G559), .Z(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(G860), .B2(new_n626), .ZN(G148));
  NAND4_X1  g202(.A1(new_n613), .A2(new_n614), .A3(new_n618), .A4(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G868), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G868), .B2(new_n560), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n467), .A2(new_n477), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  INV_X1    g209(.A(G2100), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n485), .A2(G123), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n469), .A2(G111), .ZN(new_n639));
  OAI21_X1  g214(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n640));
  INV_X1    g215(.A(G135), .ZN(new_n641));
  OAI221_X1 g216(.A(new_n638), .B1(new_n639), .B2(new_n640), .C1(new_n641), .C2(new_n481), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2096), .Z(new_n643));
  NAND3_X1  g218(.A1(new_n636), .A2(new_n637), .A3(new_n643), .ZN(G156));
  INV_X1    g219(.A(KEYINPUT14), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2427), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2430), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n649), .B1(new_n648), .B2(new_n647), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT85), .ZN(new_n652));
  XOR2_X1   g227(.A(G2443), .B(G2446), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n650), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2451), .B(G2454), .Z(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(G14), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n655), .A2(new_n658), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(G401));
  XOR2_X1   g238(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(KEYINPUT17), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n664), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2072), .B(G2078), .Z(new_n671));
  INV_X1    g246(.A(new_n664), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n671), .B1(new_n667), .B2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n670), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2096), .B(G2100), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XNOR2_X1  g251(.A(G1961), .B(G1966), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT87), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1956), .B(G2474), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT20), .Z(new_n685));
  OR2_X1    g260(.A1(new_n678), .A2(new_n680), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n686), .A2(new_n683), .A3(new_n681), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n685), .B(new_n687), .C1(new_n683), .C2(new_n686), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT88), .B(KEYINPUT89), .Z(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G1981), .B(G1986), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n690), .B(new_n695), .ZN(G229));
  NOR2_X1   g271(.A1(G16), .A2(G19), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n560), .B2(G16), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(G1341), .Z(new_n699));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G26), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT28), .Z(new_n702));
  NAND2_X1  g277(.A1(new_n485), .A2(G128), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT94), .ZN(new_n704));
  OAI21_X1  g279(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n705));
  INV_X1    g280(.A(G116), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(G2105), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(new_n482), .B2(G140), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n702), .B1(new_n709), .B2(G29), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(G2067), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT98), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n700), .A2(G27), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G164), .B2(new_n700), .ZN(new_n714));
  INV_X1    g289(.A(G2078), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n699), .B(new_n711), .C1(new_n712), .C2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n700), .A2(G33), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT25), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G139), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(new_n481), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n467), .A2(G127), .ZN(new_n724));
  NAND2_X1  g299(.A1(G115), .A2(G2104), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n469), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT95), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n718), .B1(new_n728), .B2(new_n700), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n729), .A2(G2072), .B1(new_n712), .B2(new_n716), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G2072), .B2(new_n729), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n717), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(G171), .A2(G16), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G5), .B2(G16), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n734), .A2(KEYINPUT97), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n734), .A2(KEYINPUT97), .ZN(new_n736));
  OR3_X1    g311(.A1(new_n735), .A2(new_n736), .A3(G1961), .ZN(new_n737));
  NOR2_X1   g312(.A1(G160), .A2(new_n700), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n700), .B1(KEYINPUT24), .B2(G34), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(KEYINPUT24), .B2(G34), .ZN(new_n740));
  OAI21_X1  g315(.A(G2084), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT96), .ZN(new_n742));
  OAI21_X1  g317(.A(G1961), .B1(new_n735), .B2(new_n736), .ZN(new_n743));
  AND3_X1   g318(.A1(new_n737), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NOR3_X1   g319(.A1(new_n738), .A2(G2084), .A3(new_n740), .ZN(new_n745));
  INV_X1    g320(.A(G16), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G21), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G168), .B2(new_n746), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n745), .B1(G1966), .B2(new_n748), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n700), .A2(G32), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n482), .A2(G141), .B1(G105), .B2(new_n477), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n485), .A2(G129), .ZN(new_n752));
  NAND3_X1  g327(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT26), .Z(new_n754));
  NAND3_X1  g329(.A1(new_n751), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n750), .B1(new_n755), .B2(G29), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT27), .B(G1996), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT30), .B(G28), .ZN(new_n760));
  OR2_X1    g335(.A1(KEYINPUT31), .A2(G11), .ZN(new_n761));
  NAND2_X1  g336(.A1(KEYINPUT31), .A2(G11), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n760), .A2(new_n700), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n642), .B2(new_n700), .ZN(new_n764));
  NOR3_X1   g339(.A1(new_n758), .A2(new_n759), .A3(new_n764), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n749), .B(new_n765), .C1(G1966), .C2(new_n748), .ZN(new_n766));
  NOR2_X1   g341(.A1(G4), .A2(G16), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n625), .B2(G16), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G1348), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  AND3_X1   g345(.A1(new_n732), .A2(new_n744), .A3(new_n770), .ZN(new_n771));
  OR2_X1    g346(.A1(G29), .A2(G35), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n492), .B2(new_n700), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n773), .A2(KEYINPUT29), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(KEYINPUT29), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G2090), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT99), .ZN(new_n779));
  OAI21_X1  g354(.A(KEYINPUT100), .B1(new_n776), .B2(new_n777), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT102), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT101), .B(KEYINPUT23), .Z(new_n782));
  NAND2_X1  g357(.A1(new_n746), .A2(G20), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n580), .B2(new_n746), .ZN(new_n785));
  INV_X1    g360(.A(G1956), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT100), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n774), .A2(new_n788), .A3(G2090), .A4(new_n775), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n780), .A2(new_n781), .A3(new_n787), .A4(new_n789), .ZN(new_n790));
  AND3_X1   g365(.A1(new_n771), .A2(new_n779), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n746), .A2(G23), .ZN(new_n792));
  AND3_X1   g367(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n792), .B1(new_n793), .B2(new_n746), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT33), .B(G1976), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT92), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n746), .A2(G22), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT93), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G166), .B2(new_n746), .ZN(new_n802));
  INV_X1    g377(.A(G1971), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  AND3_X1   g379(.A1(new_n798), .A2(new_n799), .A3(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(G6), .A2(G16), .ZN(new_n806));
  INV_X1    g381(.A(G305), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(G16), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT32), .B(G1981), .Z(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n805), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(KEYINPUT34), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT34), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n805), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n700), .A2(G25), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n482), .A2(G131), .ZN(new_n816));
  OAI21_X1  g391(.A(KEYINPUT90), .B1(G95), .B2(G2105), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  NOR3_X1   g393(.A1(KEYINPUT90), .A2(G95), .A3(G2105), .ZN(new_n819));
  OAI221_X1 g394(.A(G2104), .B1(G107), .B2(new_n469), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n485), .A2(G119), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n816), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n815), .B1(new_n823), .B2(new_n700), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT91), .Z(new_n825));
  XOR2_X1   g400(.A(KEYINPUT35), .B(G1991), .Z(new_n826));
  AND2_X1   g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n825), .A2(new_n826), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n746), .A2(G24), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n605), .B2(new_n746), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(G1986), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n827), .A2(new_n828), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n812), .A2(new_n814), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(KEYINPUT36), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT36), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n812), .A2(new_n835), .A3(new_n814), .A4(new_n832), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n780), .A2(new_n787), .A3(new_n789), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT102), .ZN(new_n839));
  AND3_X1   g414(.A1(new_n791), .A2(new_n837), .A3(new_n839), .ZN(G311));
  NAND3_X1  g415(.A1(new_n791), .A2(new_n837), .A3(new_n839), .ZN(G150));
  AOI22_X1  g416(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n842), .A2(new_n520), .ZN(new_n843));
  INV_X1    g418(.A(G93), .ZN(new_n844));
  INV_X1    g419(.A(G55), .ZN(new_n845));
  OAI22_X1  g420(.A1(new_n541), .A2(new_n844), .B1(new_n543), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g421(.A(KEYINPUT103), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n518), .A2(G93), .B1(new_n509), .B2(G55), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT103), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n848), .B(new_n849), .C1(new_n520), .C2(new_n842), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(new_n559), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n843), .A2(new_n846), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n853), .A2(new_n555), .A3(new_n557), .A4(new_n558), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT38), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n625), .A2(G559), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT39), .ZN(new_n859));
  AOI21_X1  g434(.A(G860), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(new_n859), .B2(new_n858), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n851), .A2(G860), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(KEYINPUT37), .Z(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(G145));
  XOR2_X1   g439(.A(KEYINPUT105), .B(G37), .Z(new_n865));
  OAI21_X1  g440(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n866));
  INV_X1    g441(.A(G118), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n866), .B1(new_n867), .B2(G2105), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n485), .A2(G130), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT104), .ZN(new_n870));
  AOI211_X1 g445(.A(new_n868), .B(new_n870), .C1(G142), .C2(new_n482), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n822), .B(new_n633), .Z(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n502), .A2(new_n504), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n494), .A2(new_n497), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n709), .B(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n755), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n879), .A2(new_n727), .ZN(new_n880));
  INV_X1    g455(.A(new_n728), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n877), .A2(new_n878), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n877), .A2(new_n878), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n873), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(G160), .B(new_n642), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(G162), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n879), .A2(new_n728), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n882), .B(new_n883), .C1(new_n726), .C2(new_n723), .ZN(new_n889));
  INV_X1    g464(.A(new_n873), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n885), .A2(new_n887), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n887), .B1(new_n885), .B2(new_n891), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n865), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g470(.A(KEYINPUT110), .ZN(new_n896));
  INV_X1    g471(.A(G868), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n851), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT109), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n899), .A2(KEYINPUT109), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n605), .A2(G288), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n793), .B1(new_n601), .B2(new_n604), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n902), .A2(G166), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(G166), .B1(new_n903), .B2(new_n902), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n905), .A2(new_n906), .A3(KEYINPUT108), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT108), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n902), .A2(new_n903), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(G303), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n908), .B1(new_n910), .B2(new_n904), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n907), .A2(new_n911), .A3(new_n807), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT108), .B1(new_n905), .B2(new_n906), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n910), .A2(new_n908), .A3(new_n904), .ZN(new_n914));
  AOI21_X1  g489(.A(G305), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n900), .B(new_n901), .C1(new_n912), .C2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n807), .B1(new_n907), .B2(new_n911), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n913), .A2(G305), .A3(new_n914), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n917), .A2(KEYINPUT109), .A3(new_n899), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n852), .A2(new_n628), .A3(new_n854), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n628), .B1(new_n852), .B2(new_n854), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT106), .B1(new_n619), .B2(new_n580), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n625), .A2(G299), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n619), .A2(KEYINPUT106), .A3(new_n580), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n921), .B1(new_n924), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n928), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT41), .B1(new_n931), .B2(new_n925), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT41), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n926), .A2(new_n933), .A3(new_n927), .A4(new_n928), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n930), .B1(new_n935), .B2(new_n924), .ZN(new_n936));
  INV_X1    g511(.A(new_n924), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n937), .A2(new_n921), .A3(new_n932), .A4(new_n934), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n920), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n938), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n940), .A2(new_n919), .A3(new_n916), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n896), .B(new_n898), .C1(new_n942), .C2(new_n897), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n897), .B1(new_n939), .B2(new_n941), .ZN(new_n944));
  INV_X1    g519(.A(new_n898), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT110), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n943), .A2(new_n946), .ZN(G295));
  OAI21_X1  g522(.A(new_n898), .B1(new_n942), .B2(new_n897), .ZN(G331));
  NAND2_X1  g523(.A1(G168), .A2(G171), .ZN(new_n949));
  NAND3_X1  g524(.A1(G286), .A2(new_n549), .A3(new_n546), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n855), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n949), .A2(new_n852), .A3(new_n854), .A4(new_n950), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n932), .A2(new_n954), .A3(new_n934), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n929), .A2(new_n953), .A3(new_n952), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n917), .A2(new_n918), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT111), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n912), .A2(new_n915), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT111), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n960), .A2(new_n961), .A3(new_n956), .A4(new_n955), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n865), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n964), .B1(new_n957), .B2(new_n958), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n963), .A2(KEYINPUT43), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(G37), .B1(new_n957), .B2(new_n958), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT43), .B1(new_n963), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT44), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT43), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n963), .A2(new_n971), .A3(new_n965), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n971), .B1(new_n963), .B2(new_n967), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n970), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n969), .A2(new_n974), .ZN(G397));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT120), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n479), .A2(new_n478), .A3(G40), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT114), .B1(new_n476), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT114), .ZN(new_n981));
  AOI211_X1 g556(.A(new_n981), .B(new_n978), .C1(new_n470), .C2(new_n475), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G2084), .ZN(new_n984));
  INV_X1    g559(.A(G1384), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT50), .B1(new_n876), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n987));
  AOI211_X1 g562(.A(new_n987), .B(G1384), .C1(new_n874), .C2(new_n875), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n984), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n977), .B1(new_n983), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G1966), .ZN(new_n991));
  XNOR2_X1  g566(.A(KEYINPUT113), .B(KEYINPUT45), .ZN(new_n992));
  NOR3_X1   g567(.A1(G164), .A2(G1384), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n994), .B1(new_n876), .B2(new_n985), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n991), .B1(new_n983), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT70), .B1(new_n474), .B2(G2105), .ZN(new_n998));
  AOI211_X1 g573(.A(new_n464), .B(new_n469), .C1(new_n473), .C2(new_n465), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n979), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n981), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n476), .A2(KEYINPUT114), .A3(new_n979), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n987), .B1(G164), .B2(G1384), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n876), .A2(KEYINPUT50), .A3(new_n985), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1003), .A2(KEYINPUT120), .A3(new_n984), .A4(new_n1006), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n990), .A2(new_n997), .A3(G168), .A4(new_n1007), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n1008), .A2(G8), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n990), .A2(new_n997), .A3(new_n1007), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(G286), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n976), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1008), .A2(G8), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1013), .A2(KEYINPUT51), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT62), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1011), .ZN(new_n1016));
  OAI21_X1  g591(.A(KEYINPUT51), .B1(new_n1016), .B2(new_n1013), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT62), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1009), .A2(new_n976), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1981), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n521), .A2(new_n540), .A3(G86), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n509), .A2(G48), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n596), .A2(new_n1021), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT118), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n588), .A2(KEYINPUT118), .A3(new_n1021), .A4(new_n596), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n597), .A2(G1981), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT49), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n876), .A2(new_n985), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n980), .B2(new_n982), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1028), .A2(KEYINPUT49), .A3(new_n1029), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1032), .A2(G8), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n793), .A2(G1976), .ZN(new_n1038));
  INV_X1    g613(.A(G1976), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT52), .B1(G288), .B2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1035), .A2(G8), .A3(new_n1038), .A4(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1037), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1035), .A2(G8), .A3(new_n1038), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT52), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1043), .A2(KEYINPUT117), .A3(KEYINPUT52), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1042), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n992), .ZN(new_n1049));
  XOR2_X1   g624(.A(KEYINPUT112), .B(G1384), .Z(new_n1050));
  AOI21_X1  g625(.A(new_n1050), .B1(new_n874), .B2(new_n875), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1033), .A2(new_n1049), .B1(new_n1051), .B2(KEYINPUT45), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1003), .A2(new_n1052), .ZN(new_n1053));
  AOI22_X1  g628(.A1(new_n1001), .A2(new_n1002), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n1053), .A2(new_n803), .B1(new_n1054), .B2(new_n777), .ZN(new_n1055));
  INV_X1    g630(.A(G8), .ZN(new_n1056));
  AND2_X1   g631(.A1(KEYINPUT119), .A2(G8), .ZN(new_n1057));
  OAI21_X1  g632(.A(G8), .B1(new_n514), .B2(new_n523), .ZN(new_n1058));
  XNOR2_X1  g633(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1059), .B1(G303), .B2(G8), .ZN(new_n1062));
  OR2_X1    g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  OAI22_X1  g638(.A1(new_n1055), .A2(new_n1056), .B1(new_n1057), .B2(new_n1063), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n1061), .A2(new_n1062), .A3(new_n1057), .ZN(new_n1065));
  OAI22_X1  g640(.A1(new_n980), .A2(new_n982), .B1(new_n986), .B2(new_n988), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1066), .A2(G2090), .ZN(new_n1067));
  AOI21_X1  g642(.A(G1971), .B1(new_n1003), .B2(new_n1052), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1065), .B(G8), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1064), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1048), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(new_n1053), .B2(G2078), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1072), .A2(G2078), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1003), .B(new_n1075), .C1(new_n993), .C2(new_n995), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1076), .B1(G1961), .B2(new_n1054), .ZN(new_n1077));
  OAI21_X1  g652(.A(G171), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1071), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1015), .A2(new_n1020), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1063), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1037), .A2(new_n1041), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT117), .B1(new_n1043), .B2(KEYINPUT52), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1043), .A2(KEYINPUT117), .A3(KEYINPUT52), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1082), .B(new_n1083), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(KEYINPUT122), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1063), .B(G8), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT63), .ZN(new_n1089));
  NOR2_X1   g664(.A1(G286), .A2(new_n1056), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1010), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT121), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1010), .A2(KEYINPUT121), .A3(new_n1090), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1089), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT122), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1048), .A2(new_n1096), .A3(new_n1082), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1087), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT63), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1010), .A2(KEYINPUT121), .A3(new_n1090), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT121), .B1(new_n1010), .B2(new_n1090), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1099), .B1(new_n1071), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1098), .A2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(KEYINPUT56), .B(G2072), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1003), .A2(new_n1052), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(G1956), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n574), .A2(new_n578), .A3(KEYINPUT123), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n579), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1111), .B(new_n1112), .C1(new_n569), .C2(new_n568), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1110), .B(new_n1109), .C1(new_n570), .C2(new_n579), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT124), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1115), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1108), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1066), .A2(new_n786), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1003), .A2(new_n1052), .A3(new_n1105), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(G2067), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1003), .A2(new_n1124), .A3(new_n1034), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(G1348), .B2(new_n1054), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1126), .A2(new_n625), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1119), .B1(new_n1123), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT61), .ZN(new_n1129));
  AND2_X1   g704(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1106), .A2(new_n1107), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1122), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1129), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT60), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1126), .A2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1125), .B(KEYINPUT60), .C1(G1348), .C2(new_n1054), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1135), .A2(new_n625), .A3(new_n1136), .ZN(new_n1137));
  OAI211_X1 g712(.A(KEYINPUT61), .B(new_n1123), .C1(new_n1108), .C2(new_n1118), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1133), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT59), .ZN(new_n1140));
  XOR2_X1   g715(.A(KEYINPUT58), .B(G1341), .Z(new_n1141));
  NAND2_X1  g716(.A1(new_n1035), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(G1996), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1003), .A2(new_n1143), .A3(new_n1052), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1140), .B1(new_n1145), .B2(new_n560), .ZN(new_n1146));
  AOI211_X1 g721(.A(KEYINPUT59), .B(new_n559), .C1(new_n1142), .C2(new_n1144), .ZN(new_n1147));
  OAI22_X1  g722(.A1(new_n1146), .A2(new_n1147), .B1(new_n625), .B2(new_n1136), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1128), .B1(new_n1139), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT54), .ZN(new_n1151));
  XNOR2_X1  g726(.A(G171), .B(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1051), .A2(new_n992), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT126), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n979), .B1(new_n469), .B2(new_n468), .ZN(new_n1155));
  OR3_X1    g730(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1154), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  AOI211_X1 g733(.A(new_n1072), .B(G2078), .C1(new_n1051), .C2(KEYINPUT45), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1152), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1054), .A2(G1961), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n1161), .A2(KEYINPUT125), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1161), .A2(KEYINPUT125), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1160), .B(new_n1073), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1152), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1165));
  AND4_X1   g740(.A1(new_n1048), .A2(new_n1070), .A3(new_n1164), .A4(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1149), .A2(new_n1150), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1035), .A2(G8), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1037), .A2(new_n1039), .A3(new_n793), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1168), .B1(new_n1169), .B2(new_n1028), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1088), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1170), .B1(new_n1171), .B2(new_n1048), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1080), .A2(new_n1104), .A3(new_n1167), .A4(new_n1172), .ZN(new_n1173));
  AND2_X1   g748(.A1(new_n1003), .A2(new_n1153), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n709), .A2(G2067), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n704), .A2(new_n1124), .A3(new_n708), .ZN(new_n1176));
  AND2_X1   g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n755), .B(G1996), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1180), .ZN(new_n1181));
  XOR2_X1   g756(.A(new_n822), .B(new_n826), .Z(new_n1182));
  OAI21_X1  g757(.A(new_n1174), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(G290), .A2(G1986), .ZN(new_n1184));
  AND2_X1   g759(.A1(G290), .A2(G1986), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1174), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1183), .A2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n1187), .B(KEYINPUT115), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1173), .A2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1174), .B1(new_n1178), .B2(new_n755), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1174), .A2(new_n1143), .ZN(new_n1191));
  AND2_X1   g766(.A1(new_n1191), .A2(KEYINPUT46), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1191), .A2(KEYINPUT46), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1190), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n1194), .B(KEYINPUT47), .ZN(new_n1195));
  AND2_X1   g770(.A1(new_n1174), .A2(new_n1184), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1196), .A2(KEYINPUT48), .ZN(new_n1197));
  OR2_X1    g772(.A1(new_n1196), .A2(KEYINPUT48), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1183), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n823), .A2(new_n826), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1176), .B1(new_n1181), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n1174), .ZN(new_n1202));
  AND3_X1   g777(.A1(new_n1195), .A2(new_n1199), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1189), .A2(new_n1203), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g779(.A1(G227), .A2(new_n462), .ZN(new_n1206));
  AND2_X1   g780(.A1(new_n662), .A2(new_n1206), .ZN(new_n1207));
  OR2_X1    g781(.A1(new_n1207), .A2(KEYINPUT127), .ZN(new_n1208));
  NAND2_X1  g782(.A1(new_n1207), .A2(KEYINPUT127), .ZN(new_n1209));
  AOI21_X1  g783(.A(G229), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  OAI211_X1 g784(.A(new_n894), .B(new_n1210), .C1(new_n972), .C2(new_n973), .ZN(G225));
  INV_X1    g785(.A(G225), .ZN(G308));
endmodule


