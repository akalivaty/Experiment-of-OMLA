//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n787, new_n788, new_n789, new_n790, new_n791, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n818, new_n819, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1017, new_n1018, new_n1019, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1087;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT3), .B1(new_n190), .B2(G107), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G104), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n190), .A2(G107), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n191), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G101), .ZN(new_n197));
  INV_X1    g011(.A(G101), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n191), .A2(new_n194), .A3(new_n198), .A4(new_n195), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n197), .A2(KEYINPUT4), .A3(new_n199), .ZN(new_n200));
  OR2_X1    g014(.A1(KEYINPUT2), .A2(G113), .ZN(new_n201));
  NAND2_X1  g015(.A1(KEYINPUT2), .A2(G113), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(G116), .A2(G119), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(G116), .A2(G119), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n206), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n201), .B(new_n202), .C1(new_n208), .C2(new_n204), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT4), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n196), .A2(new_n211), .A3(G101), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n200), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT80), .ZN(new_n214));
  XNOR2_X1  g028(.A(G110), .B(G122), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT80), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n200), .A2(new_n216), .A3(new_n210), .A4(new_n212), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT5), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n218), .B1(new_n205), .B2(new_n206), .ZN(new_n219));
  INV_X1    g033(.A(G119), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n218), .A2(new_n220), .A3(G116), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G113), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n209), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n190), .A2(G107), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n193), .A2(G104), .ZN(new_n225));
  OAI21_X1  g039(.A(G101), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n199), .A2(new_n226), .ZN(new_n227));
  OR2_X1    g041(.A1(new_n223), .A2(new_n227), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n214), .A2(new_n215), .A3(new_n217), .A4(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G143), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G146), .ZN(new_n231));
  INV_X1    g045(.A(G128), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n231), .B1(KEYINPUT1), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(G143), .B(G146), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n233), .B1(new_n234), .B2(KEYINPUT1), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n230), .A2(G146), .ZN(new_n236));
  INV_X1    g050(.A(G146), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(G143), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n232), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT76), .B(G125), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n235), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n237), .A2(G143), .ZN(new_n242));
  AND2_X1   g056(.A1(KEYINPUT0), .A2(G128), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n242), .A2(new_n231), .A3(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT0), .B(G128), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n244), .B1(new_n234), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G125), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT76), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT76), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G125), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n241), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G224), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n254), .A2(G953), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT7), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n215), .B(KEYINPUT8), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n199), .A2(new_n226), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n258), .B1(new_n259), .B2(new_n223), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT82), .ZN(new_n261));
  INV_X1    g075(.A(G116), .ZN(new_n262));
  NOR3_X1   g076(.A1(new_n262), .A2(KEYINPUT5), .A3(G119), .ZN(new_n263));
  INV_X1    g077(.A(G113), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT5), .B1(new_n208), .B2(new_n204), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n221), .A2(KEYINPUT82), .A3(G113), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n227), .B1(new_n268), .B2(new_n209), .ZN(new_n269));
  OAI22_X1  g083(.A1(new_n253), .A2(new_n257), .B1(new_n260), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT81), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n252), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n246), .A2(KEYINPUT81), .A3(new_n251), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n272), .A2(new_n241), .A3(new_n273), .A4(new_n257), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT83), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n273), .A2(new_n241), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n277), .A2(KEYINPUT83), .A3(new_n272), .A4(new_n257), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n270), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT84), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n229), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n276), .A2(new_n278), .ZN(new_n282));
  INV_X1    g096(.A(new_n270), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n282), .A2(new_n283), .A3(new_n280), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n189), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n214), .A2(new_n217), .A3(new_n228), .ZN(new_n286));
  INV_X1    g100(.A(new_n215), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(KEYINPUT6), .A3(new_n229), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n277), .A2(new_n272), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n290), .B(new_n255), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT6), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n286), .A2(new_n292), .A3(new_n287), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n289), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n188), .B1(new_n285), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n282), .A2(new_n283), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT84), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n279), .A2(new_n280), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n229), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n289), .A2(new_n291), .A3(new_n293), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n299), .A2(new_n189), .A3(new_n300), .A4(new_n187), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n295), .A2(KEYINPUT85), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n285), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT85), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n303), .A2(new_n304), .A3(new_n300), .A4(new_n187), .ZN(new_n305));
  OAI21_X1  g119(.A(G214), .B1(G237), .B2(G902), .ZN(new_n306));
  INV_X1    g120(.A(G952), .ZN(new_n307));
  AOI211_X1 g121(.A(G953), .B(new_n307), .C1(G234), .C2(G237), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT67), .B(G953), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n189), .B1(G234), .B2(G237), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(KEYINPUT96), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT21), .B(G898), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n308), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n302), .A2(new_n305), .A3(new_n306), .A4(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(G113), .B(G122), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n318), .B(new_n190), .ZN(new_n319));
  INV_X1    g133(.A(G953), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT67), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT67), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G953), .ZN(new_n323));
  INV_X1    g137(.A(G237), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n321), .A2(new_n323), .A3(G214), .A4(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n230), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n309), .A2(G143), .A3(G214), .A4(new_n324), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G131), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT64), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT64), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G131), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT88), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT88), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n328), .A2(new_n336), .A3(new_n333), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n330), .A2(new_n332), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n326), .A2(new_n327), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n335), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G140), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n341), .B1(new_n248), .B2(new_n250), .ZN(new_n342));
  NOR2_X1   g156(.A1(G125), .A2(G140), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT16), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OR2_X1    g158(.A1(KEYINPUT16), .A2(G140), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n345), .B1(new_n248), .B2(new_n250), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(G146), .A3(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(G125), .B(G140), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT19), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT89), .ZN(new_n351));
  OR2_X1    g165(.A1(new_n350), .A2(KEYINPUT89), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n349), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n343), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n354), .B1(new_n240), .B2(new_n341), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n353), .B1(new_n355), .B2(new_n350), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n340), .B(new_n348), .C1(G146), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(KEYINPUT18), .A2(G131), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n326), .A2(new_n327), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n328), .A2(KEYINPUT18), .A3(G131), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n349), .A2(new_n237), .ZN(new_n361));
  OAI211_X1 g175(.A(G146), .B(new_n354), .C1(new_n240), .C2(new_n341), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n361), .B1(new_n362), .B2(KEYINPUT86), .ZN(new_n363));
  INV_X1    g177(.A(new_n342), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT86), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n364), .A2(new_n365), .A3(G146), .A4(new_n354), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n363), .A2(KEYINPUT87), .A3(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(KEYINPUT87), .B1(new_n363), .B2(new_n366), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n359), .B(new_n360), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n319), .B1(new_n357), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n360), .A2(new_n359), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n363), .A2(new_n366), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT87), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n373), .B1(new_n376), .B2(new_n367), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n344), .A2(new_n347), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n237), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n348), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n335), .A2(new_n337), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n380), .B1(new_n381), .B2(KEYINPUT17), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT17), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n335), .A2(new_n383), .A3(new_n337), .A4(new_n339), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n377), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(KEYINPUT90), .B1(new_n385), .B2(new_n319), .ZN(new_n386));
  INV_X1    g200(.A(new_n380), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n336), .B1(new_n328), .B2(new_n333), .ZN(new_n388));
  AOI211_X1 g202(.A(KEYINPUT88), .B(new_n338), .C1(new_n326), .C2(new_n327), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT17), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n384), .A2(new_n387), .A3(new_n390), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n391), .A2(new_n370), .A3(KEYINPUT90), .A4(new_n319), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n372), .B1(new_n386), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT20), .ZN(new_n395));
  NOR2_X1   g209(.A1(G475), .A2(G902), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n391), .A2(new_n319), .A3(new_n370), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT90), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n371), .B1(new_n400), .B2(new_n392), .ZN(new_n401));
  INV_X1    g215(.A(new_n396), .ZN(new_n402));
  OAI21_X1  g216(.A(KEYINPUT20), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n397), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n319), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n391), .A2(new_n370), .ZN(new_n406));
  AOI22_X1  g220(.A1(new_n400), .A2(new_n392), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(G475), .B1(new_n407), .B2(G902), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT93), .ZN(new_n409));
  INV_X1    g223(.A(G122), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G116), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n262), .A2(G122), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n411), .B1(new_n412), .B2(KEYINPUT14), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT92), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n410), .A2(G116), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT14), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI211_X1 g231(.A(KEYINPUT92), .B(KEYINPUT14), .C1(new_n410), .C2(G116), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n413), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n409), .B1(new_n419), .B2(new_n193), .ZN(new_n420));
  INV_X1    g234(.A(new_n418), .ZN(new_n421));
  AOI21_X1  g235(.A(KEYINPUT92), .B1(new_n412), .B2(KEYINPUT14), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g237(.A(KEYINPUT93), .B(G107), .C1(new_n423), .C2(new_n413), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n230), .A2(G128), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n232), .A2(G143), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G134), .ZN(new_n429));
  XNOR2_X1  g243(.A(G128), .B(G143), .ZN(new_n430));
  INV_X1    g244(.A(G134), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n411), .A2(new_n412), .A3(new_n193), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT91), .ZN(new_n435));
  OR2_X1    g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n434), .A2(new_n435), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n433), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n425), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n430), .A2(KEYINPUT13), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n441), .B(G134), .C1(KEYINPUT13), .C2(new_n426), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n411), .A2(new_n412), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(G107), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n434), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n442), .A2(new_n445), .A3(new_n432), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n440), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(KEYINPUT9), .B(G234), .ZN(new_n448));
  INV_X1    g262(.A(G217), .ZN(new_n449));
  NOR3_X1   g263(.A1(new_n448), .A2(new_n449), .A3(G953), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(KEYINPUT95), .B1(new_n447), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n438), .B1(new_n420), .B2(new_n424), .ZN(new_n453));
  INV_X1    g267(.A(new_n446), .ZN(new_n454));
  OAI211_X1 g268(.A(KEYINPUT95), .B(new_n451), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n453), .A2(new_n454), .ZN(new_n457));
  AOI21_X1  g271(.A(KEYINPUT94), .B1(new_n457), .B2(new_n450), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT94), .ZN(new_n459));
  NOR4_X1   g273(.A1(new_n453), .A2(new_n454), .A3(new_n459), .A4(new_n451), .ZN(new_n460));
  OAI22_X1  g274(.A1(new_n452), .A2(new_n456), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G478), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n461), .B(new_n189), .C1(KEYINPUT15), .C2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(KEYINPUT15), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT95), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n465), .B1(new_n457), .B2(new_n450), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n440), .A2(new_n450), .A3(new_n446), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n459), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n457), .A2(KEYINPUT94), .A3(new_n450), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n466), .A2(new_n455), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n464), .B1(new_n470), .B2(G902), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n463), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n404), .A2(new_n408), .A3(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n317), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n220), .A2(KEYINPUT74), .A3(G128), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n232), .A2(G119), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(KEYINPUT24), .B(G110), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT75), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT74), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n482), .B1(new_n232), .B2(G119), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n478), .A2(new_n480), .A3(new_n481), .A4(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(new_n477), .A3(new_n476), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT75), .B1(new_n485), .B2(new_n479), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT23), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n477), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n220), .A2(G128), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n232), .A2(KEYINPUT23), .A3(G119), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI22_X1  g305(.A1(new_n484), .A2(new_n486), .B1(G110), .B2(new_n491), .ZN(new_n492));
  AOI211_X1 g306(.A(new_n237), .B(new_n346), .C1(new_n355), .C2(KEYINPUT16), .ZN(new_n493));
  AOI21_X1  g307(.A(G146), .B1(new_n344), .B2(new_n347), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n485), .A2(new_n479), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT77), .B(G110), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n497), .A2(new_n488), .A3(new_n489), .A4(new_n490), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n361), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n348), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G137), .ZN(new_n502));
  AND2_X1   g316(.A1(G221), .A2(G234), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n321), .A2(new_n323), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT78), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT78), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n309), .A2(new_n506), .A3(new_n503), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT22), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n505), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n508), .B1(new_n505), .B2(new_n507), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n502), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n505), .A2(new_n507), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT22), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n505), .A2(new_n507), .A3(new_n508), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n514), .A3(G137), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n501), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n495), .A2(new_n500), .A3(new_n515), .A4(new_n511), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(new_n189), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT25), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT25), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n517), .A2(new_n521), .A3(new_n189), .A4(new_n518), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n449), .B1(G234), .B2(new_n189), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n520), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n523), .A2(G902), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n517), .A2(new_n518), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT30), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT11), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n529), .B1(new_n431), .B2(G137), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n431), .A2(G137), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n502), .A2(KEYINPUT11), .A3(G134), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(G131), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT66), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT66), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n533), .A2(new_n536), .A3(G131), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n532), .A2(new_n531), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT65), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n539), .A2(new_n338), .A3(new_n540), .A4(new_n530), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT65), .B1(new_n533), .B2(new_n333), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n246), .B1(new_n538), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n502), .A2(G134), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n329), .B1(new_n545), .B2(new_n531), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(new_n235), .B2(new_n239), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n528), .B1(new_n544), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n543), .A2(new_n547), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n535), .A2(new_n537), .B1(new_n541), .B2(new_n542), .ZN(new_n551));
  OAI211_X1 g365(.A(KEYINPUT30), .B(new_n550), .C1(new_n551), .C2(new_n246), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n549), .A2(new_n210), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n210), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n554), .B(new_n550), .C1(new_n551), .C2(new_n246), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT26), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n321), .A2(new_n323), .A3(G210), .A4(new_n324), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT27), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT27), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n309), .A2(new_n559), .A3(G210), .A4(new_n324), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n556), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n558), .A2(new_n560), .A3(new_n556), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(G101), .A3(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n563), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n198), .B1(new_n565), .B2(new_n561), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(KEYINPUT68), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n553), .A2(new_n555), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(KEYINPUT31), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT31), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n572), .A2(new_n555), .A3(new_n553), .A4(new_n568), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT28), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n555), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n210), .B1(new_n544), .B2(new_n548), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n580), .A2(new_n555), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n579), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n567), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n576), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(G472), .A2(G902), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(KEYINPUT32), .A3(new_n587), .ZN(new_n588));
  XOR2_X1   g402(.A(KEYINPUT70), .B(KEYINPUT32), .Z(new_n589));
  AOI22_X1  g403(.A1(new_n574), .A2(new_n575), .B1(new_n584), .B2(new_n567), .ZN(new_n590));
  INV_X1    g404(.A(new_n587), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n567), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n583), .B1(new_n580), .B2(new_n555), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n594), .B1(new_n595), .B2(new_n578), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n553), .A2(new_n555), .A3(new_n567), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT29), .ZN(new_n599));
  AOI21_X1  g413(.A(G902), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n578), .B(KEYINPUT73), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n567), .A2(new_n599), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n555), .A2(KEYINPUT71), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n540), .B1(new_n604), .B2(new_n338), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n533), .A2(KEYINPUT65), .A3(new_n333), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n533), .A2(new_n536), .A3(G131), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n536), .B1(new_n533), .B2(G131), .ZN(new_n608));
  OAI22_X1  g422(.A1(new_n605), .A2(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n246), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT71), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n611), .A2(new_n612), .A3(new_n554), .A4(new_n550), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n603), .A2(new_n580), .A3(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT72), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n614), .A2(new_n615), .A3(KEYINPUT28), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n615), .B1(new_n614), .B2(KEYINPUT28), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n601), .B(new_n602), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n600), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(G472), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n527), .B1(new_n593), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(G221), .B1(new_n448), .B2(G902), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(G469), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n624), .A2(new_n189), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n309), .A2(G227), .ZN(new_n626));
  XOR2_X1   g440(.A(G110), .B(G140), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(G128), .B1(new_n242), .B2(new_n231), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT1), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n630), .B1(new_n236), .B2(new_n238), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n629), .B1(new_n631), .B2(new_n233), .ZN(new_n632));
  OAI21_X1  g446(.A(KEYINPUT10), .B1(new_n632), .B2(new_n227), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT10), .ZN(new_n634));
  AOI21_X1  g448(.A(KEYINPUT1), .B1(new_n242), .B2(new_n231), .ZN(new_n635));
  AOI22_X1  g449(.A1(new_n630), .A2(G128), .B1(new_n230), .B2(G146), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n239), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n259), .A2(new_n634), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n200), .A2(new_n610), .A3(new_n212), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n639), .A2(new_n551), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n551), .B1(new_n639), .B2(new_n640), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n628), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n639), .A2(new_n551), .A3(new_n640), .ZN(new_n644));
  INV_X1    g458(.A(new_n628), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n259), .A2(new_n637), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n632), .A2(new_n227), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n648), .A2(new_n609), .A3(KEYINPUT12), .ZN(new_n649));
  AOI21_X1  g463(.A(KEYINPUT12), .B1(new_n648), .B2(new_n609), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n644), .B(new_n645), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(G902), .B1(new_n643), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n625), .B1(new_n652), .B2(new_n624), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n644), .B1(new_n649), .B2(new_n650), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n628), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n644), .A2(KEYINPUT79), .A3(new_n645), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n639), .A2(new_n640), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n656), .B1(new_n551), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(KEYINPUT79), .B1(new_n644), .B2(new_n645), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n655), .B(G469), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n623), .B1(new_n653), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n475), .A2(new_n621), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT97), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G101), .ZN(G3));
  OAI21_X1  g478(.A(G472), .B1(new_n590), .B2(G902), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n665), .B1(new_n591), .B2(new_n590), .ZN(new_n666));
  INV_X1    g480(.A(new_n661), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n666), .A2(new_n527), .A3(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n306), .ZN(new_n669));
  AOI211_X1 g483(.A(new_n669), .B(new_n315), .C1(new_n295), .C2(new_n301), .ZN(new_n670));
  INV_X1    g484(.A(new_n467), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n457), .A2(new_n450), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT33), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n462), .A2(G902), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT98), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n470), .A2(new_n677), .A3(KEYINPUT33), .ZN(new_n678));
  AOI21_X1  g492(.A(KEYINPUT98), .B1(new_n461), .B2(new_n673), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n675), .B(new_n676), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  AOI21_X1  g494(.A(G478), .B1(new_n461), .B2(new_n189), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  AOI22_X1  g496(.A1(new_n404), .A2(new_n408), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n668), .A2(new_n670), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT34), .B(G104), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT99), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n684), .B(new_n686), .ZN(G6));
  AND2_X1   g501(.A1(new_n408), .A2(new_n472), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n670), .A2(new_n404), .A3(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n668), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n691), .B(KEYINPUT100), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT101), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT35), .B(G107), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G9));
  INV_X1    g509(.A(new_n666), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n511), .A2(new_n515), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT36), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n697), .A2(new_n698), .A3(new_n495), .A4(new_n500), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n501), .B1(KEYINPUT36), .B2(new_n516), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n699), .A2(new_n700), .A3(new_n525), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n524), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT102), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT102), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n524), .A2(new_n702), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n475), .A2(new_n661), .A3(new_n696), .A4(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(KEYINPUT37), .B(G110), .Z(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G12));
  AOI21_X1  g524(.A(new_n395), .B1(new_n394), .B2(new_n396), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n401), .A2(KEYINPUT20), .A3(new_n402), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n408), .B(new_n472), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(G900), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n308), .B1(new_n313), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g529(.A(KEYINPUT103), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n620), .A2(new_n592), .A3(new_n588), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT103), .ZN(new_n718));
  INV_X1    g532(.A(new_n715), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n688), .A2(new_n404), .A3(new_n718), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n295), .A2(new_n301), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n306), .ZN(new_n722));
  INV_X1    g536(.A(new_n523), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n723), .B1(new_n519), .B2(KEYINPUT25), .ZN(new_n724));
  AOI211_X1 g538(.A(KEYINPUT102), .B(new_n701), .C1(new_n724), .C2(new_n522), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n705), .B1(new_n524), .B2(new_n702), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n661), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n722), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n716), .A2(new_n717), .A3(new_n720), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G128), .ZN(G30));
  OAI22_X1  g544(.A1(new_n386), .A2(new_n393), .B1(new_n319), .B2(new_n385), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n189), .ZN(new_n732));
  AOI22_X1  g546(.A1(new_n397), .A2(new_n403), .B1(new_n732), .B2(G475), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n472), .A2(new_n306), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n553), .A2(new_n555), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n594), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n737), .B(new_n189), .C1(new_n614), .C2(new_n594), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(G472), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n588), .A2(new_n592), .A3(new_n739), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n735), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n715), .B(KEYINPUT39), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n667), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(KEYINPUT40), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n725), .A2(new_n726), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n302), .A2(new_n305), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT38), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n741), .A2(new_n744), .A3(new_n745), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G143), .ZN(G45));
  NAND4_X1  g564(.A1(new_n728), .A2(new_n683), .A3(new_n717), .A4(new_n719), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G146), .ZN(G48));
  NOR2_X1   g566(.A1(new_n652), .A2(new_n624), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n643), .A2(new_n651), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(new_n624), .A3(new_n189), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n754), .A2(new_n622), .A3(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n757), .A2(new_n527), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n588), .A2(new_n592), .ZN(new_n759));
  INV_X1    g573(.A(G472), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n760), .B1(new_n600), .B2(new_n618), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n758), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n408), .B1(new_n711), .B2(new_n712), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n680), .A2(new_n682), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n670), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(KEYINPUT41), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G113), .ZN(G15));
  OR2_X1    g582(.A1(new_n762), .A2(new_n689), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G116), .ZN(G18));
  NOR2_X1   g584(.A1(new_n759), .A2(new_n761), .ZN(new_n771));
  AOI211_X1 g585(.A(G469), .B(G902), .C1(new_n643), .C2(new_n651), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n753), .A2(new_n772), .A3(new_n623), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n707), .A2(new_n721), .A3(new_n306), .A4(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n404), .A2(new_n408), .A3(new_n473), .A4(new_n316), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n771), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(new_n220), .ZN(G21));
  INV_X1    g591(.A(new_n734), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n757), .A2(new_n315), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n763), .A2(new_n778), .A3(new_n779), .A4(new_n721), .ZN(new_n780));
  INV_X1    g594(.A(new_n527), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n601), .B1(new_n616), .B2(new_n617), .ZN(new_n782));
  AOI22_X1  g596(.A1(new_n782), .A2(new_n567), .B1(new_n575), .B2(new_n574), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n781), .B(new_n665), .C1(new_n783), .C2(new_n591), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n780), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(new_n410), .ZN(G24));
  NAND3_X1  g600(.A1(new_n721), .A2(new_n306), .A3(new_n773), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(new_n745), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n665), .B1(new_n783), .B2(new_n591), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n788), .A2(new_n790), .A3(new_n683), .A4(new_n719), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G125), .ZN(G27));
  INV_X1    g606(.A(KEYINPUT42), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n669), .B1(new_n302), .B2(new_n305), .ZN(new_n794));
  AOI211_X1 g608(.A(KEYINPUT104), .B(new_n623), .C1(new_n653), .C2(new_n660), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT104), .ZN(new_n796));
  INV_X1    g610(.A(new_n625), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n660), .A2(new_n756), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n796), .B1(new_n798), .B2(new_n622), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n717), .A2(new_n794), .A3(new_n800), .A4(new_n781), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n763), .A2(new_n764), .A3(new_n719), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n793), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT105), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT32), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n805), .B1(new_n590), .B2(new_n591), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n588), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n804), .B(new_n781), .C1(new_n807), .C2(new_n761), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n620), .A2(new_n588), .A3(new_n806), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n804), .B1(new_n810), .B2(new_n781), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n794), .A2(new_n800), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n763), .A2(new_n764), .A3(new_n719), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(new_n814), .A3(KEYINPUT42), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n803), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G131), .ZN(G33));
  AND2_X1   g631(.A1(new_n716), .A2(new_n720), .ZN(new_n818));
  INV_X1    g632(.A(new_n801), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G134), .ZN(G36));
  INV_X1    g635(.A(KEYINPUT43), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n822), .B1(new_n763), .B2(KEYINPUT106), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n677), .B1(new_n470), .B2(KEYINPUT33), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n461), .A2(KEYINPUT98), .A3(new_n673), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n674), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n681), .B1(new_n826), .B2(new_n676), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n763), .A2(new_n827), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n823), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n823), .A2(new_n828), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n696), .A2(new_n745), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT44), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n794), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n655), .B1(new_n658), .B2(new_n659), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT45), .ZN(new_n838));
  OR2_X1    g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n624), .B1(new_n837), .B2(new_n838), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n625), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n841), .A2(KEYINPUT46), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n756), .B1(new_n841), .B2(KEYINPUT46), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n622), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n844), .A2(new_n742), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n833), .A2(new_n834), .ZN(new_n846));
  OR3_X1    g660(.A1(new_n836), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(G137), .ZN(G39));
  OR2_X1    g662(.A1(new_n844), .A2(KEYINPUT47), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n844), .A2(KEYINPUT47), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n814), .A2(new_n771), .A3(new_n527), .A4(new_n794), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(new_n341), .ZN(G42));
  NOR3_X1   g668(.A1(new_n527), .A2(new_n669), .A3(new_n623), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT107), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n753), .A2(new_n772), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT49), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR4_X1   g673(.A1(new_n856), .A2(new_n763), .A3(new_n827), .A4(new_n859), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(KEYINPUT108), .ZN(new_n861));
  AOI211_X1 g675(.A(new_n740), .B(new_n748), .C1(new_n858), .C2(new_n857), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n667), .A2(new_n703), .A3(new_n715), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n735), .A2(new_n721), .A3(new_n740), .A4(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n729), .A2(new_n751), .A3(new_n791), .A4(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT52), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n728), .A2(new_n717), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n774), .A2(new_n789), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n814), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n871), .A2(KEYINPUT52), .A3(new_n729), .A4(new_n865), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n781), .B1(new_n807), .B2(new_n761), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT105), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n808), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n794), .A2(new_n800), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n877), .A2(new_n802), .A3(new_n793), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n813), .A2(new_n621), .A3(new_n814), .ZN(new_n879));
  AOI22_X1  g693(.A1(new_n876), .A2(new_n878), .B1(new_n879), .B2(new_n793), .ZN(new_n880));
  INV_X1    g694(.A(new_n474), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n881), .A2(new_n788), .A3(new_n717), .A4(new_n316), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n763), .A2(new_n778), .A3(new_n721), .ZN(new_n883));
  INV_X1    g697(.A(new_n784), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n883), .A2(new_n884), .A3(new_n779), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n766), .A2(new_n769), .A3(new_n882), .A4(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n880), .A2(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n873), .A2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n317), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n889), .A2(KEYINPUT109), .A3(new_n404), .A4(new_n688), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT109), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n891), .B1(new_n317), .B2(new_n713), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n890), .A2(new_n668), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n668), .A2(new_n889), .A3(new_n683), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n893), .A2(new_n662), .A3(new_n708), .A4(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT111), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n463), .A2(new_n471), .A3(new_n719), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n727), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n717), .A2(new_n898), .A3(new_n733), .A4(new_n794), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(KEYINPUT110), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n763), .A2(new_n727), .A3(new_n897), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT110), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n901), .A2(new_n902), .A3(new_n717), .A4(new_n794), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n716), .A2(new_n720), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n683), .A2(new_n719), .A3(new_n794), .A4(new_n800), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n789), .A2(new_n745), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  OAI22_X1  g723(.A1(new_n906), .A2(new_n801), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n896), .B1(new_n905), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n877), .A2(new_n802), .ZN(new_n912));
  AOI22_X1  g726(.A1(new_n818), .A2(new_n819), .B1(new_n912), .B2(new_n908), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n913), .A2(KEYINPUT111), .A3(new_n904), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n895), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n888), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT112), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT53), .B1(new_n873), .B2(new_n917), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n916), .B(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(KEYINPUT54), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT53), .B1(new_n888), .B2(new_n915), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT114), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n922), .B1(new_n880), .B2(new_n886), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n762), .B1(new_n689), .B2(new_n765), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n924), .A2(new_n776), .A3(new_n785), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n816), .A2(KEYINPUT114), .A3(new_n925), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n923), .A2(new_n873), .A3(KEYINPUT53), .A4(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n895), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n912), .A2(new_n908), .ZN(new_n929));
  AND4_X1   g743(.A1(KEYINPUT111), .A2(new_n904), .A3(new_n820), .A4(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(KEYINPUT111), .B1(new_n913), .B2(new_n904), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n927), .B1(KEYINPUT113), .B2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT113), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n934), .B(new_n928), .C1(new_n930), .C2(new_n931), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n921), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  XOR2_X1   g750(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n920), .A2(new_n938), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n794), .A2(new_n773), .ZN(new_n940));
  INV_X1    g754(.A(new_n308), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n740), .A2(new_n527), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n683), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n945), .A2(new_n307), .A3(G953), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n941), .B1(new_n829), .B2(new_n830), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n884), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n947), .A2(new_n876), .A3(new_n940), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n949), .A2(KEYINPUT48), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n831), .A2(new_n308), .A3(new_n940), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n951), .A2(KEYINPUT48), .A3(new_n812), .ZN(new_n952));
  OAI221_X1 g766(.A(new_n946), .B1(new_n787), .B2(new_n948), .C1(new_n950), .C2(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n947), .A2(new_n884), .A3(new_n794), .ZN(new_n954));
  AOI22_X1  g768(.A1(new_n849), .A2(new_n850), .B1(new_n623), .B2(new_n857), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n733), .A2(new_n827), .ZN(new_n957));
  OAI22_X1  g771(.A1(new_n951), .A2(new_n909), .B1(new_n943), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g773(.A(KEYINPUT117), .B(KEYINPUT50), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n773), .A2(new_n669), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n748), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n947), .A2(new_n884), .A3(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT116), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n947), .A2(KEYINPUT116), .A3(new_n884), .A4(new_n962), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n960), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT50), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n963), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n959), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT51), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n953), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n959), .B(KEYINPUT51), .C1(new_n967), .C2(new_n969), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT118), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n973), .A2(new_n974), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n972), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(KEYINPUT119), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT119), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n979), .B(new_n972), .C1(new_n975), .C2(new_n976), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n939), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  NOR2_X1   g795(.A1(G952), .A2(G953), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n863), .B1(new_n981), .B2(new_n982), .ZN(G75));
  NOR2_X1   g797(.A1(new_n309), .A2(G952), .ZN(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n936), .A2(new_n189), .ZN(new_n986));
  AOI21_X1  g800(.A(KEYINPUT56), .B1(new_n986), .B2(G210), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n289), .A2(new_n293), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(new_n291), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(KEYINPUT120), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT55), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n985), .B1(new_n987), .B2(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n992), .B1(new_n987), .B2(new_n991), .ZN(G51));
  NAND2_X1  g807(.A1(new_n932), .A2(KEYINPUT113), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT53), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n995), .B1(new_n868), .B2(new_n872), .ZN(new_n996));
  AND3_X1   g810(.A1(new_n996), .A2(new_n926), .A3(new_n923), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n994), .A2(new_n997), .A3(new_n935), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n873), .A2(new_n887), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n995), .B1(new_n932), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n937), .ZN(new_n1002));
  OAI21_X1  g816(.A(KEYINPUT121), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT121), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n936), .A2(new_n1004), .A3(new_n937), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1003), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n625), .B(KEYINPUT57), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n755), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n839), .A2(new_n840), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  AND3_X1   g826(.A1(new_n986), .A2(KEYINPUT122), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(KEYINPUT122), .B1(new_n986), .B2(new_n1012), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n984), .B1(new_n1010), .B2(new_n1015), .ZN(G54));
  NAND3_X1  g830(.A1(new_n986), .A2(KEYINPUT58), .A3(G475), .ZN(new_n1017));
  AND2_X1   g831(.A1(new_n1017), .A2(new_n401), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1017), .A2(new_n401), .ZN(new_n1019));
  NOR3_X1   g833(.A1(new_n1018), .A2(new_n1019), .A3(new_n984), .ZN(G60));
  NAND2_X1  g834(.A1(G478), .A2(G902), .ZN(new_n1021));
  XOR2_X1   g835(.A(new_n1021), .B(KEYINPUT59), .Z(new_n1022));
  AOI21_X1  g836(.A(new_n1022), .B1(new_n920), .B2(new_n938), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n985), .B1(new_n1023), .B2(new_n826), .ZN(new_n1024));
  AOI211_X1 g838(.A(new_n674), .B(new_n1022), .C1(new_n824), .C2(new_n825), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1024), .B1(new_n1007), .B2(new_n1025), .ZN(G63));
  NAND2_X1  g840(.A1(new_n699), .A2(new_n700), .ZN(new_n1027));
  XNOR2_X1  g841(.A(new_n1027), .B(KEYINPUT124), .ZN(new_n1028));
  INV_X1    g842(.A(KEYINPUT123), .ZN(new_n1029));
  NAND2_X1  g843(.A1(G217), .A2(G902), .ZN(new_n1030));
  XNOR2_X1  g844(.A(new_n1030), .B(KEYINPUT60), .ZN(new_n1031));
  INV_X1    g845(.A(new_n1031), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1029), .B1(new_n1001), .B2(new_n1032), .ZN(new_n1033));
  AOI211_X1 g847(.A(KEYINPUT123), .B(new_n1031), .C1(new_n998), .C2(new_n1000), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1028), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g849(.A(KEYINPUT123), .B1(new_n936), .B2(new_n1031), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n517), .A2(new_n518), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1001), .A2(new_n1029), .A3(new_n1032), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n1035), .A2(new_n1039), .A3(new_n985), .ZN(new_n1040));
  INV_X1    g854(.A(KEYINPUT61), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g856(.A1(new_n1035), .A2(new_n1039), .A3(KEYINPUT61), .A4(new_n985), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1042), .A2(new_n1043), .ZN(G66));
  OAI21_X1  g858(.A(G953), .B1(new_n314), .B2(new_n254), .ZN(new_n1045));
  NOR2_X1   g859(.A1(new_n895), .A2(new_n886), .ZN(new_n1046));
  OAI21_X1  g860(.A(new_n1045), .B1(new_n1046), .B2(new_n310), .ZN(new_n1047));
  INV_X1    g861(.A(G898), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n988), .B1(new_n1048), .B2(new_n310), .ZN(new_n1049));
  XOR2_X1   g863(.A(new_n1047), .B(new_n1049), .Z(G69));
  AND2_X1   g864(.A1(new_n871), .A2(new_n729), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1051), .A2(new_n749), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n1052), .A2(KEYINPUT62), .ZN(new_n1053));
  OR2_X1    g867(.A1(new_n1052), .A2(KEYINPUT62), .ZN(new_n1054));
  NAND3_X1  g868(.A1(new_n621), .A2(new_n743), .A3(new_n794), .ZN(new_n1055));
  AOI21_X1  g869(.A(new_n1055), .B1(new_n944), .B2(new_n713), .ZN(new_n1056));
  NOR2_X1   g870(.A1(new_n853), .A2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g871(.A1(new_n847), .A2(new_n1053), .A3(new_n1054), .A4(new_n1057), .ZN(new_n1058));
  NAND2_X1  g872(.A1(new_n1058), .A2(new_n309), .ZN(new_n1059));
  NAND2_X1  g873(.A1(new_n549), .A2(new_n552), .ZN(new_n1060));
  XOR2_X1   g874(.A(new_n1060), .B(new_n356), .Z(new_n1061));
  INV_X1    g875(.A(KEYINPUT125), .ZN(new_n1062));
  OAI21_X1  g876(.A(G900), .B1(new_n1062), .B2(G227), .ZN(new_n1063));
  AOI22_X1  g877(.A1(new_n1059), .A2(new_n1061), .B1(new_n310), .B2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g878(.A1(new_n1051), .A2(new_n816), .A3(new_n820), .ZN(new_n1065));
  NAND2_X1  g879(.A1(new_n876), .A2(new_n883), .ZN(new_n1066));
  OAI21_X1  g880(.A(new_n1066), .B1(new_n836), .B2(new_n846), .ZN(new_n1067));
  INV_X1    g881(.A(new_n845), .ZN(new_n1068));
  AOI211_X1 g882(.A(new_n853), .B(new_n1065), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1069));
  OR3_X1    g883(.A1(new_n1069), .A2(new_n310), .A3(new_n1061), .ZN(new_n1070));
  NAND3_X1  g884(.A1(new_n1064), .A2(new_n1070), .A3(KEYINPUT125), .ZN(new_n1071));
  XOR2_X1   g885(.A(KEYINPUT126), .B(G900), .Z(new_n1072));
  AOI211_X1 g886(.A(new_n1061), .B(new_n1072), .C1(new_n1064), .C2(new_n1070), .ZN(new_n1073));
  INV_X1    g887(.A(G227), .ZN(new_n1074));
  OAI21_X1  g888(.A(new_n310), .B1(new_n1074), .B2(new_n714), .ZN(new_n1075));
  OAI21_X1  g889(.A(new_n1071), .B1(new_n1073), .B2(new_n1075), .ZN(G72));
  NAND2_X1  g890(.A1(G472), .A2(G902), .ZN(new_n1077));
  XOR2_X1   g891(.A(new_n1077), .B(KEYINPUT63), .Z(new_n1078));
  AND4_X1   g892(.A1(new_n597), .A2(new_n919), .A3(new_n737), .A4(new_n1078), .ZN(new_n1079));
  OR3_X1    g893(.A1(new_n1058), .A2(new_n895), .A3(new_n886), .ZN(new_n1080));
  AOI21_X1  g894(.A(new_n737), .B1(new_n1080), .B2(new_n1078), .ZN(new_n1081));
  INV_X1    g895(.A(new_n1078), .ZN(new_n1082));
  AOI21_X1  g896(.A(new_n1082), .B1(new_n1069), .B2(new_n1046), .ZN(new_n1083));
  OAI21_X1  g897(.A(new_n985), .B1(new_n1083), .B2(new_n597), .ZN(new_n1084));
  NAND2_X1  g898(.A1(new_n1084), .A2(KEYINPUT127), .ZN(new_n1085));
  INV_X1    g899(.A(KEYINPUT127), .ZN(new_n1086));
  OAI211_X1 g900(.A(new_n1086), .B(new_n985), .C1(new_n1083), .C2(new_n597), .ZN(new_n1087));
  AOI211_X1 g901(.A(new_n1079), .B(new_n1081), .C1(new_n1085), .C2(new_n1087), .ZN(G57));
endmodule


