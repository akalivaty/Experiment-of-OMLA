//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 0 0 0 1 0 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1307, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n202), .A2(G50), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n223));
  INV_X1    g0023(.A(G58), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  INV_X1    g0025(.A(G97), .ZN(new_n226));
  INV_X1    g0026(.A(G257), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n207), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n210), .B(new_n216), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT64), .Z(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G226), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT66), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(KEYINPUT7), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT3), .B(G33), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n250), .B1(new_n251), .B2(G20), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT72), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n214), .A2(KEYINPUT7), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n253), .B1(new_n251), .B2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT3), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n254), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n260), .A2(KEYINPUT72), .A3(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n252), .A2(new_n255), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G68), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n224), .A2(new_n218), .ZN(new_n265));
  OAI21_X1  g0065(.A(G20), .B1(new_n265), .B2(new_n201), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G20), .A2(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G159), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n264), .A2(KEYINPUT16), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT16), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT73), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n273), .B1(new_n258), .B2(G33), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n256), .A2(KEYINPUT73), .A3(KEYINPUT3), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(new_n259), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n261), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n218), .B1(new_n277), .B2(new_n252), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n272), .B1(new_n278), .B2(new_n269), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n213), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n271), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G13), .ZN(new_n283));
  NOR3_X1   g0083(.A1(new_n283), .A2(new_n214), .A3(G1), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(new_n281), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT8), .B(G58), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G1), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G20), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n283), .A2(G1), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G20), .ZN(new_n293));
  OAI22_X1  g0093(.A1(new_n286), .A2(new_n291), .B1(new_n293), .B2(new_n288), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT74), .ZN(new_n296));
  OR2_X1    g0096(.A1(G223), .A2(G1698), .ZN(new_n297));
  INV_X1    g0097(.A(G226), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G1698), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n257), .A2(new_n297), .A3(new_n259), .A4(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G87), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AND2_X1   g0104(.A1(G1), .A2(G13), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G41), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G41), .ZN(new_n308));
  INV_X1    g0108(.A(G45), .ZN(new_n309));
  AOI21_X1  g0109(.A(G1), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n307), .A2(G274), .A3(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n289), .B1(G41), .B2(G45), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n307), .A2(G232), .A3(new_n312), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(G200), .B1(new_n304), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n307), .B1(new_n300), .B2(new_n301), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n311), .A2(new_n313), .ZN(new_n317));
  NOR3_X1   g0117(.A1(new_n316), .A2(new_n317), .A3(G190), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n296), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G190), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n304), .A2(new_n314), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G200), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(new_n316), .B2(new_n317), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n321), .A2(new_n323), .A3(KEYINPUT74), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n282), .A2(new_n295), .A3(new_n319), .A4(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT17), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n281), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n269), .B1(new_n263), .B2(G68), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n328), .B1(new_n329), .B2(KEYINPUT16), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n294), .B1(new_n330), .B2(new_n279), .ZN(new_n331));
  INV_X1    g0131(.A(G169), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n332), .B1(new_n304), .B2(new_n314), .ZN(new_n333));
  INV_X1    g0133(.A(G179), .ZN(new_n334));
  NOR3_X1   g0134(.A1(new_n316), .A2(new_n317), .A3(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(KEYINPUT18), .B1(new_n331), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n282), .A2(new_n295), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT18), .ZN(new_n339));
  INV_X1    g0139(.A(new_n336), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AND3_X1   g0141(.A1(new_n321), .A2(KEYINPUT74), .A3(new_n323), .ZN(new_n342));
  AOI21_X1  g0142(.A(KEYINPUT74), .B1(new_n321), .B2(new_n323), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n331), .A2(new_n344), .A3(KEYINPUT17), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n327), .A2(new_n337), .A3(new_n341), .A4(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(G222), .A2(G1698), .ZN(new_n348));
  INV_X1    g0148(.A(G1698), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n349), .A2(G223), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n251), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n351), .B(new_n303), .C1(G77), .C2(new_n251), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n308), .A2(new_n309), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n289), .A2(new_n353), .B1(new_n305), .B2(new_n306), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G226), .ZN(new_n355));
  AND3_X1   g0155(.A1(new_n352), .A2(new_n311), .A3(new_n355), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n356), .A2(new_n334), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n214), .A2(G33), .ZN(new_n358));
  INV_X1    g0158(.A(G150), .ZN(new_n359));
  INV_X1    g0159(.A(new_n267), .ZN(new_n360));
  OAI22_X1  g0160(.A1(new_n287), .A2(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G50), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n214), .B1(new_n201), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n281), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n362), .B1(new_n289), .B2(G20), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n285), .A2(new_n365), .B1(new_n362), .B2(new_n284), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n356), .B2(G169), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n357), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n356), .A2(new_n322), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n370), .B1(G190), .B2(new_n356), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n367), .A2(KEYINPUT69), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n367), .A2(KEYINPUT69), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n373), .A2(KEYINPUT9), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT9), .ZN(new_n376));
  OR2_X1    g0176(.A1(new_n367), .A2(KEYINPUT69), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n376), .B1(new_n377), .B2(new_n372), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n371), .B1(new_n375), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT70), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT10), .B1(new_n370), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(KEYINPUT9), .B1(new_n373), .B2(new_n374), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n377), .A2(new_n376), .A3(new_n372), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n386), .A2(new_n381), .A3(new_n371), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n369), .B1(new_n383), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n298), .A2(new_n349), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n225), .A2(G1698), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n257), .A2(new_n389), .A3(new_n259), .A4(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G33), .A2(G97), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n303), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT13), .ZN(new_n395));
  INV_X1    g0195(.A(G274), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(new_n305), .B2(new_n306), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n354), .A2(G238), .B1(new_n397), .B2(new_n310), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n394), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n307), .B1(new_n391), .B2(new_n392), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n307), .A2(G238), .A3(new_n312), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n311), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(KEYINPUT13), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(G200), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n399), .A2(new_n403), .A3(G190), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n267), .A2(G50), .B1(G20), .B2(new_n218), .ZN(new_n407));
  INV_X1    g0207(.A(G77), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n407), .B1(new_n408), .B2(new_n358), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n409), .A2(KEYINPUT11), .A3(new_n281), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n285), .A2(G68), .A3(new_n290), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT12), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(new_n284), .B2(new_n218), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n293), .A2(KEYINPUT12), .A3(G68), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n410), .B(new_n411), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT11), .B1(new_n409), .B2(new_n281), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n405), .A2(new_n406), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT71), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n405), .A2(KEYINPUT71), .A3(new_n417), .A4(new_n406), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n417), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT14), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n404), .A2(new_n424), .A3(G169), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n334), .B2(new_n404), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n424), .B1(new_n404), .B2(G169), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n423), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n422), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n354), .A2(G244), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n311), .ZN(new_n432));
  OR2_X1    g0232(.A1(new_n432), .A2(KEYINPUT67), .ZN(new_n433));
  NOR2_X1   g0233(.A1(G232), .A2(G1698), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n349), .A2(G238), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n251), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n436), .B(new_n303), .C1(G107), .C2(new_n251), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n432), .A2(KEYINPUT67), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n433), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n439), .A2(G200), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n288), .A2(new_n267), .B1(G20), .B2(G77), .ZN(new_n441));
  XNOR2_X1  g0241(.A(KEYINPUT15), .B(G87), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n358), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n328), .B1(new_n441), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n285), .A2(G77), .A3(new_n290), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT68), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n293), .A2(new_n448), .A3(G77), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT68), .B1(new_n284), .B2(new_n408), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n447), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(new_n439), .B2(new_n320), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n440), .A2(new_n453), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n439), .A2(G179), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n452), .B1(new_n439), .B2(new_n332), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AND4_X1   g0257(.A1(new_n347), .A2(new_n388), .A3(new_n430), .A4(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(G250), .A2(G1698), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n460), .B1(new_n227), .B2(G1698), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n461), .A2(new_n251), .ZN(new_n462));
  INV_X1    g0262(.A(G294), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n256), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n303), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n309), .A2(G1), .ZN(new_n466));
  NAND2_X1  g0266(.A1(KEYINPUT5), .A2(G41), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n470), .A2(G264), .A3(new_n307), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT5), .B(G41), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n397), .A2(new_n466), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n465), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G169), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT80), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT80), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n474), .A2(new_n477), .A3(G169), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n476), .B(new_n478), .C1(new_n334), .C2(new_n474), .ZN(new_n479));
  INV_X1    g0279(.A(G107), .ZN(new_n480));
  AOI21_X1  g0280(.A(KEYINPUT79), .B1(new_n480), .B2(G20), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT23), .ZN(new_n482));
  OR2_X1    g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n482), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n483), .A2(new_n484), .B1(G116), .B2(new_n444), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n257), .A2(new_n259), .A3(new_n214), .A4(G87), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT22), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(new_n214), .A3(G87), .ZN(new_n488));
  OAI21_X1  g0288(.A(KEYINPUT77), .B1(new_n260), .B2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT77), .ZN(new_n490));
  NOR3_X1   g0290(.A1(new_n220), .A2(KEYINPUT22), .A3(G20), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n251), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  AOI221_X4 g0292(.A(KEYINPUT78), .B1(new_n486), .B2(KEYINPUT22), .C1(new_n489), .C2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT78), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n489), .A2(new_n492), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n486), .A2(KEYINPUT22), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n485), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT24), .ZN(new_n499));
  NOR3_X1   g0299(.A1(new_n260), .A2(KEYINPUT77), .A3(new_n488), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n490), .B1(new_n251), .B2(new_n491), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n496), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT78), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n495), .A2(new_n494), .A3(new_n496), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT24), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n505), .A2(new_n506), .A3(new_n485), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n328), .B1(new_n499), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n284), .A2(new_n480), .ZN(new_n509));
  OR2_X1    g0309(.A1(new_n509), .A2(KEYINPUT25), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n256), .A2(G1), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n284), .A2(new_n281), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G107), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n509), .A2(KEYINPUT25), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n510), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n479), .B1(new_n508), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n506), .B1(new_n505), .B2(new_n485), .ZN(new_n518));
  INV_X1    g0318(.A(new_n485), .ZN(new_n519));
  AOI211_X1 g0319(.A(KEYINPUT24), .B(new_n519), .C1(new_n503), .C2(new_n504), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n281), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  OR2_X1    g0321(.A1(new_n474), .A2(new_n320), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n474), .A2(G200), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n522), .A2(new_n515), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n517), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G250), .A2(G1698), .ZN(new_n527));
  NAND2_X1  g0327(.A1(KEYINPUT4), .A2(G244), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n527), .B1(new_n528), .B2(G1698), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n251), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G283), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(G244), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n533), .A2(G1698), .ZN(new_n534));
  AOI21_X1  g0334(.A(KEYINPUT4), .B1(new_n251), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n303), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n470), .A2(G257), .A3(new_n307), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n537), .A2(new_n473), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT75), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n251), .A2(new_n529), .B1(G33), .B2(G283), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n534), .A2(new_n257), .A3(new_n259), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT4), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n307), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n537), .A2(new_n473), .ZN(new_n546));
  OAI21_X1  g0346(.A(KEYINPUT75), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n540), .A2(new_n547), .A3(G200), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n293), .A2(G97), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n512), .B2(G97), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT6), .ZN(new_n552));
  AND2_X1   g0352(.A1(G97), .A2(G107), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n552), .B1(new_n553), .B2(new_n204), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n480), .A2(KEYINPUT6), .A3(G97), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n556), .A2(G20), .B1(G77), .B2(new_n267), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n260), .A2(new_n214), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n558), .A2(new_n250), .B1(new_n276), .B2(new_n261), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n557), .B1(new_n559), .B2(new_n480), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n551), .B1(new_n560), .B2(new_n281), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n536), .A2(new_n538), .A3(G190), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n548), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n219), .A2(new_n349), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n533), .A2(G1698), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n257), .A2(new_n564), .A3(new_n259), .A4(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(G33), .A2(G116), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n307), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n307), .A2(G274), .A3(new_n466), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n221), .B1(new_n289), .B2(G45), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n307), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n332), .B1(new_n568), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n397), .A2(new_n466), .B1(new_n307), .B2(new_n570), .ZN(new_n574));
  NOR2_X1   g0374(.A1(G238), .A2(G1698), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n575), .B1(new_n533), .B2(G1698), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n576), .A2(new_n251), .B1(G33), .B2(G116), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n334), .B(new_n574), .C1(new_n577), .C2(new_n307), .ZN(new_n578));
  AND2_X1   g0378(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n443), .A2(new_n293), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT19), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n214), .B1(new_n392), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(G87), .B2(new_n205), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n257), .A2(new_n259), .A3(new_n214), .A4(G68), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n581), .B1(new_n358), .B2(new_n226), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n580), .B1(new_n586), .B2(new_n281), .ZN(new_n587));
  INV_X1    g0387(.A(new_n512), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n587), .B1(new_n442), .B2(new_n588), .ZN(new_n589));
  AOI221_X4 g0389(.A(new_n580), .B1(new_n512), .B2(G87), .C1(new_n586), .C2(new_n281), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n322), .B1(new_n568), .B2(new_n572), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n320), .B(new_n574), .C1(new_n577), .C2(new_n307), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n579), .A2(new_n589), .B1(new_n590), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n267), .A2(G77), .ZN(new_n595));
  INV_X1    g0395(.A(new_n556), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n595), .B1(new_n596), .B2(new_n214), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n480), .B1(new_n277), .B2(new_n252), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n281), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n550), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n536), .A2(new_n538), .A3(G179), .ZN(new_n601));
  OAI21_X1  g0401(.A(G169), .B1(new_n545), .B2(new_n546), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n563), .A2(new_n594), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n470), .A2(G270), .A3(new_n307), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n606), .A2(new_n473), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT76), .ZN(new_n608));
  INV_X1    g0408(.A(G303), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n260), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n349), .A2(G264), .ZN(new_n611));
  NOR2_X1   g0411(.A1(G257), .A2(G1698), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n257), .B(new_n259), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  AND4_X1   g0413(.A1(new_n608), .A2(new_n610), .A3(new_n613), .A4(new_n303), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n307), .B1(new_n260), .B2(new_n609), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n608), .B1(new_n615), .B2(new_n613), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n607), .B(G179), .C1(new_n614), .C2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n606), .A2(new_n473), .ZN(new_n618));
  INV_X1    g0418(.A(new_n613), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n303), .B1(new_n251), .B2(G303), .ZN(new_n620));
  OAI21_X1  g0420(.A(KEYINPUT76), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n615), .A2(new_n608), .A3(new_n613), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n618), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(KEYINPUT21), .A2(G169), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n617), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(G116), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n512), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n284), .A2(G116), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n280), .A2(new_n213), .B1(G20), .B2(new_n626), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n531), .B(new_n214), .C1(G33), .C2(new_n226), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n629), .A2(KEYINPUT20), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT20), .B1(new_n629), .B2(new_n630), .ZN(new_n632));
  OAI22_X1  g0432(.A1(new_n627), .A2(new_n628), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n625), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n607), .B1(new_n614), .B2(new_n616), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n635), .A2(new_n633), .A3(G169), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT21), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n621), .A2(new_n622), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n639), .A2(G190), .A3(new_n607), .ZN(new_n640));
  INV_X1    g0440(.A(new_n633), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n640), .B(new_n641), .C1(new_n322), .C2(new_n623), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n634), .A2(new_n638), .A3(new_n642), .ZN(new_n643));
  NOR4_X1   g0443(.A1(new_n459), .A2(new_n526), .A3(new_n605), .A4(new_n643), .ZN(G372));
  NAND3_X1  g0444(.A1(new_n422), .A2(new_n455), .A3(new_n456), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n428), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(KEYINPUT83), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n647), .A2(new_n327), .A3(new_n345), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n646), .A2(KEYINPUT83), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n337), .B(new_n341), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n383), .A2(new_n387), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n369), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n579), .A2(new_n589), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n594), .A2(new_n600), .A3(new_n603), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT26), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n594), .A2(KEYINPUT26), .A3(new_n600), .A4(new_n603), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n657), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n563), .A2(new_n594), .A3(new_n604), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n525), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n635), .A2(KEYINPUT21), .A3(G169), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n641), .B1(new_n666), .B2(new_n617), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n332), .B1(new_n639), .B2(new_n607), .ZN(new_n668));
  AOI21_X1  g0468(.A(KEYINPUT21), .B1(new_n668), .B2(new_n633), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT82), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT82), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n634), .A2(new_n671), .A3(new_n638), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n665), .A2(KEYINPUT81), .B1(new_n673), .B2(new_n517), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT81), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n525), .A2(new_n675), .A3(new_n664), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n663), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n655), .B1(new_n459), .B2(new_n677), .ZN(G369));
  NAND2_X1  g0478(.A1(new_n292), .A2(new_n214), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G213), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(G343), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n641), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n643), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n670), .A2(new_n672), .A3(new_n686), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G330), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n684), .B1(new_n508), .B2(new_n516), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n691), .A2(new_n517), .A3(new_n525), .ZN(new_n692));
  INV_X1    g0492(.A(new_n517), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n684), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n690), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n693), .A2(new_n685), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n685), .B1(new_n667), .B2(new_n669), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n698), .A2(new_n517), .A3(new_n525), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n695), .A2(new_n700), .ZN(G399));
  INV_X1    g0501(.A(new_n208), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(G41), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n205), .A2(G87), .A3(G116), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(G1), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n211), .B2(new_n704), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT28), .ZN(new_n708));
  AOI22_X1  g0508(.A1(new_n461), .A2(new_n251), .B1(G33), .B2(G294), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n471), .B1(new_n709), .B2(new_n307), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n710), .A2(new_n568), .A3(new_n572), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT30), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n545), .A2(new_n546), .A3(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n711), .A2(G179), .A3(new_n713), .A4(new_n623), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n536), .A2(new_n538), .ZN(new_n715));
  INV_X1    g0515(.A(new_n568), .ZN(new_n716));
  AOI21_X1  g0516(.A(G179), .B1(new_n716), .B2(new_n574), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n635), .A2(new_n474), .A3(new_n715), .A4(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n465), .A2(new_n471), .A3(new_n716), .A4(new_n574), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n617), .A2(new_n719), .A3(new_n715), .ZN(new_n720));
  XOR2_X1   g0520(.A(KEYINPUT84), .B(KEYINPUT30), .Z(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  OAI211_X1 g0522(.A(new_n714), .B(new_n718), .C1(new_n720), .C2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n684), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT31), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n723), .A2(KEYINPUT31), .A3(new_n684), .ZN(new_n727));
  AND3_X1   g0527(.A1(new_n634), .A2(new_n638), .A3(new_n642), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n728), .A2(new_n664), .A3(new_n685), .ZN(new_n729));
  OAI211_X1 g0529(.A(new_n726), .B(new_n727), .C1(new_n526), .C2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G330), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(KEYINPUT85), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT85), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n730), .A2(new_n733), .A3(G330), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT29), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n673), .A2(new_n517), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n522), .A2(new_n515), .A3(new_n523), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n508), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(KEYINPUT81), .B1(new_n739), .B2(new_n605), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n737), .A2(new_n740), .A3(new_n676), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n662), .ZN(new_n742));
  AOI21_X1  g0542(.A(KEYINPUT86), .B1(new_n742), .B2(new_n685), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT86), .ZN(new_n744));
  AOI211_X1 g0544(.A(new_n744), .B(new_n684), .C1(new_n741), .C2(new_n662), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n736), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n667), .A2(new_n669), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n517), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n739), .A2(new_n605), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n657), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n660), .A2(KEYINPUT88), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n661), .A2(KEYINPUT87), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n661), .A2(KEYINPUT87), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT88), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n658), .A2(new_n754), .A3(new_n659), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n751), .A2(new_n752), .A3(new_n753), .A4(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n684), .B1(new_n750), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(KEYINPUT29), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n735), .B1(new_n746), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n708), .B1(new_n759), .B2(G1), .ZN(G364));
  NOR2_X1   g0560(.A1(new_n283), .A2(G20), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n289), .B1(new_n761), .B2(G45), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n703), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n214), .A2(new_n334), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G190), .A2(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n766), .A2(new_n320), .A3(G200), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n251), .B1(new_n768), .B2(new_n408), .C1(new_n218), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n766), .A2(G190), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G200), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n320), .A2(G179), .A3(G200), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n214), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n773), .A2(new_n224), .B1(new_n226), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n771), .A2(new_n322), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n362), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n214), .A2(G179), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n780), .A2(new_n320), .A3(G200), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n480), .ZN(new_n782));
  OR4_X1    g0582(.A1(new_n770), .A2(new_n776), .A3(new_n779), .A4(new_n782), .ZN(new_n783));
  XOR2_X1   g0583(.A(KEYINPUT92), .B(KEYINPUT32), .Z(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n780), .A2(new_n767), .ZN(new_n786));
  INV_X1    g0586(.A(G159), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n785), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n786), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n789), .A2(G159), .A3(new_n784), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n780), .A2(G190), .A3(G200), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G87), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n788), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(G322), .A2(new_n772), .B1(new_n777), .B2(G326), .ZN(new_n795));
  INV_X1    g0595(.A(G283), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n795), .B1(new_n796), .B2(new_n781), .ZN(new_n797));
  INV_X1    g0597(.A(new_n775), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n798), .A2(G294), .B1(new_n792), .B2(G303), .ZN(new_n799));
  INV_X1    g0599(.A(new_n769), .ZN(new_n800));
  XNOR2_X1  g0600(.A(KEYINPUT33), .B(G317), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n251), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n768), .ZN(new_n803));
  AOI22_X1  g0603(.A1(G311), .A2(new_n803), .B1(new_n789), .B2(G329), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n799), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n783), .A2(new_n794), .B1(new_n797), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n213), .B1(G20), .B2(new_n332), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n765), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT89), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n208), .B(new_n251), .C1(G355), .C2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(KEYINPUT89), .B1(new_n205), .B2(G87), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n810), .A2(new_n811), .B1(G116), .B2(new_n208), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT90), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n212), .A2(new_n309), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n702), .A2(new_n251), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n814), .B(new_n815), .C1(new_n248), .C2(new_n309), .ZN(new_n816));
  AOI21_X1  g0616(.A(KEYINPUT91), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n813), .A2(KEYINPUT91), .A3(new_n816), .ZN(new_n818));
  NOR2_X1   g0618(.A1(G13), .A2(G33), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(G20), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(new_n807), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n821), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n808), .B1(new_n817), .B2(new_n823), .C1(new_n689), .C2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n690), .A2(new_n765), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n689), .A2(G330), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT93), .ZN(G396));
  OAI21_X1  g0629(.A(new_n684), .B1(new_n446), .B2(new_n451), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n440), .B2(new_n453), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n455), .A2(new_n456), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n455), .A2(new_n456), .A3(new_n685), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n744), .B1(new_n677), .B2(new_n684), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n742), .A2(KEYINPUT86), .A3(new_n685), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n735), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT95), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n457), .A2(new_n685), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n841), .B1(new_n742), .B2(new_n843), .ZN(new_n844));
  AOI211_X1 g0644(.A(KEYINPUT95), .B(new_n842), .C1(new_n741), .C2(new_n662), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OR3_X1    g0646(.A1(new_n839), .A2(new_n840), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n840), .B1(new_n839), .B2(new_n846), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n847), .A2(new_n765), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n807), .A2(new_n819), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n765), .B1(new_n408), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n807), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n251), .B1(new_n789), .B2(G311), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n853), .B1(new_n626), .B2(new_n768), .C1(new_n796), .C2(new_n769), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n463), .A2(new_n773), .B1(new_n778), .B2(new_n609), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n781), .A2(new_n220), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n775), .A2(new_n226), .B1(new_n791), .B2(new_n480), .ZN(new_n857));
  NOR4_X1   g0657(.A1(new_n854), .A2(new_n855), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n781), .A2(new_n218), .ZN(new_n859));
  INV_X1    g0659(.A(G132), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n251), .B1(new_n786), .B2(new_n860), .C1(new_n362), .C2(new_n791), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n859), .B(new_n861), .C1(G58), .C2(new_n798), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT94), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n800), .A2(G150), .B1(new_n803), .B2(G159), .ZN(new_n864));
  INV_X1    g0664(.A(G137), .ZN(new_n865));
  INV_X1    g0665(.A(G143), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n864), .B1(new_n778), .B2(new_n865), .C1(new_n866), .C2(new_n773), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT34), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n858), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  OAI221_X1 g0669(.A(new_n851), .B1(new_n852), .B2(new_n869), .C1(new_n836), .C2(new_n820), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n849), .A2(new_n870), .ZN(G384));
  OR2_X1    g0671(.A1(new_n556), .A2(KEYINPUT35), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n556), .A2(KEYINPUT35), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n872), .A2(G116), .A3(new_n215), .A4(new_n873), .ZN(new_n874));
  XOR2_X1   g0674(.A(new_n874), .B(KEYINPUT36), .Z(new_n875));
  OR3_X1    g0675(.A1(new_n211), .A2(new_n408), .A3(new_n265), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n362), .A2(G68), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n289), .B(G13), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT96), .ZN(new_n880));
  INV_X1    g0680(.A(new_n834), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT95), .B1(new_n677), .B2(new_n842), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n742), .A2(new_n841), .A3(new_n843), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n423), .A2(new_n684), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n429), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n422), .A2(new_n428), .A3(new_n885), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n880), .B1(new_n884), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n834), .B1(new_n844), .B2(new_n845), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n892), .A2(KEYINPUT96), .A3(new_n889), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n329), .A2(KEYINPUT16), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n294), .B1(new_n894), .B2(new_n330), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n325), .B1(new_n895), .B2(new_n682), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n895), .A2(new_n336), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT37), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n338), .A2(new_n340), .ZN(new_n899));
  INV_X1    g0699(.A(new_n682), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n338), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT37), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n899), .A2(new_n901), .A3(new_n902), .A4(new_n325), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n898), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n895), .A2(new_n682), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n346), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT38), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n904), .A2(new_n906), .A3(KEYINPUT38), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n891), .A2(new_n893), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n900), .B1(new_n337), .B2(new_n341), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n909), .A2(KEYINPUT39), .A3(new_n910), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n903), .A2(new_n898), .B1(new_n346), .B2(new_n905), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n915), .A2(KEYINPUT97), .A3(KEYINPUT38), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT97), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n910), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n899), .A2(new_n901), .A3(new_n325), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(KEYINPUT37), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n903), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n346), .A2(new_n338), .A3(new_n900), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT38), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n916), .B1(new_n918), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n914), .B1(new_n924), .B2(KEYINPUT39), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  OR2_X1    g0726(.A1(new_n428), .A2(new_n684), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n913), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n912), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n459), .B1(KEYINPUT29), .B2(new_n757), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT98), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n746), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n932), .B1(new_n746), .B2(new_n931), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n655), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n930), .B(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n835), .B1(new_n887), .B2(new_n888), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n643), .A2(new_n605), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n939), .A2(new_n517), .A3(new_n525), .A4(new_n685), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n714), .A2(new_n718), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n711), .A2(G179), .A3(new_n623), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n721), .B1(new_n942), .B2(new_n715), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n685), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(KEYINPUT100), .B1(new_n944), .B2(KEYINPUT31), .ZN(new_n945));
  AOI21_X1  g0745(.A(KEYINPUT31), .B1(new_n723), .B2(new_n684), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT100), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n940), .A2(new_n945), .A3(new_n948), .A4(new_n727), .ZN(new_n949));
  AND3_X1   g0749(.A1(new_n904), .A2(KEYINPUT38), .A3(new_n906), .ZN(new_n950));
  AOI21_X1  g0750(.A(KEYINPUT38), .B1(new_n904), .B2(new_n906), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n938), .B(new_n949), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  AND3_X1   g0754(.A1(new_n952), .A2(KEYINPUT101), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(KEYINPUT101), .B1(new_n952), .B2(new_n954), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n949), .A2(new_n938), .A3(KEYINPUT40), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n955), .A2(new_n956), .B1(new_n924), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n458), .A2(new_n949), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(new_n959), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n960), .A2(G330), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n937), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n289), .B2(new_n761), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n937), .A2(new_n962), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n879), .B1(new_n964), .B2(new_n965), .ZN(G367));
  INV_X1    g0766(.A(new_n822), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(new_n702), .B2(new_n443), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n240), .A2(new_n815), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n765), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n685), .A2(new_n590), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n971), .A2(new_n656), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n594), .A2(new_n971), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n251), .B1(new_n786), .B2(new_n865), .C1(new_n778), .C2(new_n866), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT107), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n769), .A2(new_n787), .B1(new_n768), .B2(new_n362), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n976), .B2(new_n977), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n773), .A2(new_n359), .B1(new_n791), .B2(new_n224), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n775), .A2(new_n218), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n781), .A2(new_n408), .ZN(new_n982));
  NOR4_X1   g0782(.A1(new_n979), .A2(new_n980), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT108), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n781), .A2(new_n226), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n773), .A2(new_n609), .B1(new_n480), .B2(new_n775), .ZN(new_n986));
  AOI211_X1 g0786(.A(new_n985), .B(new_n986), .C1(G311), .C2(new_n777), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n769), .A2(new_n463), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n260), .B1(new_n768), .B2(new_n796), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n988), .B(new_n989), .C1(G317), .C2(new_n789), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT46), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n791), .B2(new_n626), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n792), .A2(KEYINPUT46), .A3(G116), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n987), .A2(new_n990), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n984), .A2(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT47), .Z(new_n996));
  OAI221_X1 g0796(.A(new_n970), .B1(new_n824), .B2(new_n974), .C1(new_n996), .C2(new_n852), .ZN(new_n997));
  INV_X1    g0797(.A(new_n974), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT43), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n600), .A2(new_n603), .A3(new_n684), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT102), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n563), .B(new_n604), .C1(new_n561), .C2(new_n685), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1006), .A2(new_n699), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT103), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1008), .A2(KEYINPUT42), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1005), .A2(new_n693), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n684), .B1(new_n1010), .B2(new_n604), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(new_n1008), .B2(KEYINPUT42), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1000), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(KEYINPUT43), .B2(new_n974), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n695), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1015), .A2(new_n1006), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1009), .A2(new_n1012), .A3(new_n999), .A4(new_n998), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n1019), .B(new_n1000), .C1(new_n1009), .C2(new_n1012), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1017), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n1020), .A2(new_n1021), .B1(new_n1015), .B2(new_n1006), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1018), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1005), .B1(new_n696), .B2(new_n699), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT44), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n696), .A2(new_n699), .A3(new_n1005), .ZN(new_n1026));
  XOR2_X1   g0826(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n1027));
  XNOR2_X1  g0827(.A(new_n1026), .B(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1015), .A2(KEYINPUT105), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n694), .A2(new_n692), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n699), .B1(new_n1034), .B2(new_n698), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT106), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n690), .A2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1035), .B(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n759), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n759), .B1(new_n1033), .B2(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n703), .B(KEYINPUT41), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n763), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n997), .B1(new_n1023), .B2(new_n1042), .ZN(G387));
  NAND2_X1  g0843(.A1(new_n1038), .A2(new_n763), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n251), .A2(new_n208), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n705), .A2(new_n1045), .B1(G107), .B2(new_n208), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n237), .A2(new_n309), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n815), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n705), .ZN(new_n1049));
  AOI211_X1 g0849(.A(G45), .B(new_n1049), .C1(G68), .C2(G77), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n287), .A2(G50), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT50), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1048), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1046), .B1(new_n1047), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n764), .B1(new_n1054), .B2(new_n967), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n769), .A2(new_n287), .B1(new_n768), .B2(new_n218), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT109), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n260), .B(new_n985), .C1(G150), .C2(new_n789), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n775), .A2(new_n442), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G159), .B2(new_n777), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n772), .A2(G50), .B1(new_n792), .B2(G77), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1057), .A2(new_n1058), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n772), .A2(G317), .B1(new_n803), .B2(G303), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1063), .A2(KEYINPUT111), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G322), .A2(new_n777), .B1(new_n800), .B2(G311), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(KEYINPUT111), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT48), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n775), .A2(new_n796), .B1(new_n791), .B2(new_n463), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT110), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1069), .A2(KEYINPUT49), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n251), .B1(new_n789), .B2(G326), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1073), .B(new_n1074), .C1(new_n626), .C2(new_n781), .ZN(new_n1075));
  AOI21_X1  g0875(.A(KEYINPUT49), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1062), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1055), .B1(new_n1077), .B2(new_n807), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n1034), .B2(new_n824), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1039), .A2(new_n703), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n759), .A2(new_n1038), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1044), .B(new_n1079), .C1(new_n1080), .C2(new_n1081), .ZN(G393));
  AND2_X1   g0882(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1039), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n704), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1029), .B(new_n695), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT115), .ZN(new_n1087));
  AND3_X1   g0887(.A1(new_n1086), .A2(new_n1087), .A3(new_n1039), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1087), .B1(new_n1086), .B2(new_n1039), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1085), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n245), .A2(new_n1048), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n822), .B1(new_n226), .B2(new_n208), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n764), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(G150), .A2(new_n777), .B1(new_n772), .B2(G159), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT51), .Z(new_n1095));
  OAI22_X1  g0895(.A1(new_n769), .A2(new_n362), .B1(new_n768), .B2(new_n287), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n775), .A2(new_n408), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  XOR2_X1   g0898(.A(new_n1098), .B(KEYINPUT112), .Z(new_n1099));
  OAI21_X1  g0899(.A(new_n251), .B1(new_n786), .B2(new_n866), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n856), .B(new_n1100), .C1(G68), .C2(new_n792), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1095), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT113), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(G311), .A2(new_n772), .B1(new_n777), .B2(G317), .ZN(new_n1105));
  XOR2_X1   g0905(.A(new_n1105), .B(KEYINPUT52), .Z(new_n1106));
  AOI21_X1  g0906(.A(new_n251), .B1(new_n800), .B2(G303), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G294), .A2(new_n803), .B1(new_n789), .B2(G322), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n791), .A2(new_n796), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n782), .B(new_n1109), .C1(G116), .C2(new_n798), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .A4(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1104), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1093), .B1(new_n1113), .B2(new_n807), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n1005), .B2(new_n824), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n1086), .B2(new_n762), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(KEYINPUT114), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT114), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1118), .B(new_n1115), .C1(new_n1086), .C2(new_n762), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1090), .A2(new_n1120), .ZN(G390));
  AND2_X1   g0921(.A1(new_n949), .A2(G330), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n458), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(KEYINPUT29), .B1(new_n837), .B2(new_n838), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n758), .A2(new_n458), .ZN(new_n1126));
  OAI21_X1  g0926(.A(KEYINPUT98), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n1124), .B(new_n654), .C1(new_n1127), .C2(new_n933), .ZN(new_n1128));
  INV_X1    g0928(.A(G330), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n727), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1130), .A2(new_n946), .ZN(new_n1131));
  AOI211_X1 g0931(.A(KEYINPUT85), .B(new_n1129), .C1(new_n1131), .C2(new_n940), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n733), .B1(new_n730), .B2(G330), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n938), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n881), .B1(new_n757), .B2(new_n833), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n949), .A2(G330), .A3(new_n836), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n890), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1134), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT117), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1134), .A2(KEYINPUT117), .A3(new_n1135), .A4(new_n1137), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n889), .B1(new_n735), .B2(new_n836), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n949), .A2(new_n938), .A3(G330), .ZN(new_n1144));
  OAI211_X1 g0944(.A(KEYINPUT116), .B(new_n892), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT116), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n836), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1144), .B1(new_n1147), .B2(new_n890), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1146), .B1(new_n1148), .B2(new_n884), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1142), .A2(new_n1145), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1128), .A2(new_n1150), .ZN(new_n1151));
  AND4_X1   g0951(.A1(KEYINPUT97), .A2(new_n904), .A3(KEYINPUT38), .A4(new_n906), .ZN(new_n1152));
  AOI21_X1  g0952(.A(KEYINPUT97), .B1(new_n915), .B2(KEYINPUT38), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n921), .A2(new_n922), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n908), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1152), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1156), .B(new_n927), .C1(new_n1135), .C2(new_n890), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n928), .B1(new_n892), .B2(new_n889), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1157), .B(new_n1134), .C1(new_n1158), .C2(new_n926), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n750), .A2(new_n756), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1160), .A2(new_n685), .A3(new_n833), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n890), .B1(new_n1161), .B2(new_n834), .ZN(new_n1162));
  NOR3_X1   g0962(.A1(new_n1162), .A2(new_n928), .A3(new_n924), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n927), .B1(new_n884), .B2(new_n890), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1163), .B1(new_n1164), .B2(new_n925), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1144), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1159), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  OR2_X1    g0967(.A1(new_n1151), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n704), .B1(new_n1151), .B2(new_n1167), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1159), .B(new_n763), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1171));
  INV_X1    g0971(.A(G128), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n778), .A2(new_n1172), .B1(new_n787), .B2(new_n775), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G132), .B2(new_n772), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n791), .A2(new_n359), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT53), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n789), .A2(G125), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(KEYINPUT54), .B(G143), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n800), .A2(G137), .B1(new_n803), .B2(new_n1179), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1174), .A2(new_n1176), .A3(new_n1177), .A4(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n251), .B1(new_n781), .B2(new_n362), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT118), .Z(new_n1183));
  OAI22_X1  g0983(.A1(new_n768), .A2(new_n226), .B1(new_n786), .B2(new_n463), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n251), .B(new_n1184), .C1(G107), .C2(new_n800), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1185), .B(new_n793), .C1(new_n218), .C2(new_n781), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1097), .B1(G116), .B2(new_n772), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n796), .B2(new_n778), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n1181), .A2(new_n1183), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n807), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n765), .B1(new_n287), .B2(new_n850), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1190), .B(new_n1191), .C1(new_n926), .C2(new_n820), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1171), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1170), .A2(new_n1194), .ZN(G378));
  AND3_X1   g0995(.A1(new_n1142), .A2(new_n1145), .A3(new_n1149), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1128), .B1(new_n1167), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n957), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1129), .B1(new_n1156), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT119), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n682), .B1(new_n377), .B2(new_n372), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n388), .A2(new_n1202), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n369), .B(new_n1201), .C1(new_n383), .C2(new_n387), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(new_n1203), .A2(new_n1204), .A3(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n387), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n381), .B1(new_n386), .B2(new_n371), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n653), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n1201), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n388), .A2(new_n1202), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1205), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1200), .B1(new_n1207), .B2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1206), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1211), .A2(new_n1212), .A3(new_n1205), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1215), .A2(new_n1216), .A3(KEYINPUT119), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1214), .A2(new_n1217), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1199), .B(new_n1218), .C1(new_n955), .C2(new_n956), .ZN(new_n1219));
  OAI21_X1  g1019(.A(G330), .B1(new_n924), .B2(new_n957), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT101), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n949), .A2(new_n938), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n910), .B2(new_n909), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1221), .B1(new_n1223), .B2(new_n953), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n952), .A2(KEYINPUT101), .A3(new_n954), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1220), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1219), .B(KEYINPUT120), .C1(new_n1226), .C2(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1199), .B1(new_n955), .B2(new_n956), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT120), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1229), .A2(new_n1230), .A3(new_n1216), .A4(new_n1215), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1228), .A2(new_n930), .A3(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n930), .B1(new_n1228), .B2(new_n1231), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1197), .B(KEYINPUT57), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n703), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1228), .A2(new_n1231), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n930), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1228), .A2(new_n930), .A3(new_n1231), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT57), .B1(new_n1240), .B2(new_n1197), .ZN(new_n1241));
  OR2_X1    g1041(.A1(new_n1235), .A2(new_n1241), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n769), .A2(new_n860), .B1(new_n768), .B2(new_n865), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(G150), .A2(new_n798), .B1(new_n777), .B2(G125), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n1172), .B2(new_n773), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1243), .B(new_n1245), .C1(new_n792), .C2(new_n1179), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT59), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(G33), .A2(G41), .ZN(new_n1250));
  INV_X1    g1050(.A(G124), .ZN(new_n1251));
  OAI221_X1 g1051(.A(new_n1250), .B1(new_n786), .B2(new_n1251), .C1(new_n787), .C2(new_n781), .ZN(new_n1252));
  NOR3_X1   g1052(.A1(new_n1248), .A2(new_n1249), .A3(new_n1252), .ZN(new_n1253));
  AOI211_X1 g1053(.A(G50), .B(new_n1250), .C1(new_n260), .C2(new_n308), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n773), .A2(new_n480), .B1(new_n781), .B2(new_n224), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(G116), .B2(new_n777), .ZN(new_n1256));
  AOI211_X1 g1056(.A(G41), .B(new_n251), .C1(new_n800), .C2(G97), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n443), .A2(new_n803), .B1(new_n789), .B2(G283), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n981), .B1(G77), .B2(new_n792), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .A4(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT58), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1254), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n1261), .B2(new_n1260), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n807), .B1(new_n1253), .B2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n765), .B1(new_n362), .B2(new_n850), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1264), .B(new_n1265), .C1(new_n1218), .C2(new_n820), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(new_n1240), .B2(new_n763), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1242), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(KEYINPUT121), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT121), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1242), .A2(new_n1271), .A3(new_n1268), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1270), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(G375));
  OAI21_X1  g1074(.A(KEYINPUT122), .B1(new_n1128), .B2(new_n1150), .ZN(new_n1275));
  AND2_X1   g1075(.A1(new_n1145), .A2(new_n1149), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n655), .B(new_n1123), .C1(new_n934), .C2(new_n935), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT122), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1276), .A2(new_n1277), .A3(new_n1278), .A4(new_n1142), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1275), .A2(new_n1279), .A3(new_n1041), .A4(new_n1151), .ZN(new_n1280));
  XOR2_X1   g1080(.A(new_n1280), .B(KEYINPUT123), .Z(new_n1281));
  NAND2_X1  g1081(.A1(new_n1150), .A2(new_n763), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n765), .B1(new_n218), .B2(new_n850), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(new_n800), .A2(G116), .B1(new_n789), .B2(G303), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n480), .B2(new_n768), .ZN(new_n1285));
  OAI22_X1  g1085(.A1(new_n778), .A2(new_n463), .B1(new_n791), .B2(new_n226), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n773), .A2(new_n796), .ZN(new_n1287));
  NOR4_X1   g1087(.A1(new_n1285), .A2(new_n1286), .A3(new_n1287), .A4(new_n1059), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n982), .A2(new_n251), .ZN(new_n1289));
  XOR2_X1   g1089(.A(new_n1289), .B(KEYINPUT124), .Z(new_n1290));
  OAI22_X1  g1090(.A1(new_n773), .A2(new_n865), .B1(new_n362), .B2(new_n775), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1291), .B1(G159), .B2(new_n792), .ZN(new_n1292));
  OAI22_X1  g1092(.A1(new_n778), .A2(new_n860), .B1(new_n781), .B2(new_n224), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n251), .B1(new_n769), .B2(new_n1178), .ZN(new_n1294));
  OAI22_X1  g1094(.A1(new_n768), .A2(new_n359), .B1(new_n786), .B2(new_n1172), .ZN(new_n1295));
  NOR3_X1   g1095(.A1(new_n1293), .A2(new_n1294), .A3(new_n1295), .ZN(new_n1296));
  AOI22_X1  g1096(.A1(new_n1288), .A2(new_n1290), .B1(new_n1292), .B2(new_n1296), .ZN(new_n1297));
  OAI221_X1 g1097(.A(new_n1283), .B1(new_n852), .B2(new_n1297), .C1(new_n889), .C2(new_n820), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1282), .A2(new_n1298), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1281), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(G381));
  AOI21_X1  g1101(.A(new_n1193), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1302));
  NOR3_X1   g1102(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(new_n1303), .B(KEYINPUT125), .ZN(new_n1304));
  NOR3_X1   g1104(.A1(new_n1304), .A2(G387), .A3(G390), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1273), .A2(new_n1302), .A3(new_n1300), .A4(new_n1305), .ZN(G407));
  NAND2_X1  g1106(.A1(new_n1273), .A2(new_n1302), .ZN(new_n1307));
  OAI211_X1 g1107(.A(G407), .B(G213), .C1(G343), .C2(new_n1307), .ZN(G409));
  OAI211_X1 g1108(.A(G390), .B(new_n997), .C1(new_n1042), .C2(new_n1023), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(G387), .A2(new_n1120), .A3(new_n1090), .ZN(new_n1310));
  XOR2_X1   g1110(.A(G393), .B(G396), .Z(new_n1311));
  AND3_X1   g1111(.A1(new_n1309), .A2(new_n1310), .A3(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1311), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  OAI211_X1 g1115(.A(G378), .B(new_n1268), .C1(new_n1235), .C2(new_n1241), .ZN(new_n1316));
  OAI211_X1 g1116(.A(new_n1197), .B(new_n1041), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n763), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1317), .A2(new_n1318), .A3(new_n1266), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n1302), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1316), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT62), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n683), .A2(G213), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1128), .A2(new_n1150), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n704), .B1(new_n1324), .B2(KEYINPUT60), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1275), .A2(new_n1279), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT60), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1327), .B1(new_n1128), .B2(new_n1150), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1325), .B1(new_n1326), .B2(new_n1328), .ZN(new_n1329));
  OAI211_X1 g1129(.A(new_n1282), .B(new_n1298), .C1(G384), .C2(KEYINPUT126), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1329), .A2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(G384), .A2(KEYINPUT126), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1332), .A2(new_n1334), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1329), .A2(new_n1331), .A3(new_n1333), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1321), .A2(new_n1322), .A3(new_n1323), .A4(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT61), .ZN(new_n1339));
  AOI22_X1  g1139(.A1(new_n1316), .A2(new_n1320), .B1(G213), .B2(new_n683), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n683), .A2(G213), .A3(G2897), .ZN(new_n1341));
  AND3_X1   g1141(.A1(new_n1329), .A2(new_n1331), .A3(new_n1333), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1333), .B1(new_n1329), .B2(new_n1331), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1341), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1341), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1335), .A2(new_n1336), .A3(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1344), .A2(new_n1346), .ZN(new_n1347));
  OAI211_X1 g1147(.A(new_n1338), .B(new_n1339), .C1(new_n1340), .C2(new_n1347), .ZN(new_n1348));
  XOR2_X1   g1148(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1349));
  AOI21_X1  g1149(.A(new_n1349), .B1(new_n1340), .B2(new_n1337), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1315), .B1(new_n1348), .B2(new_n1350), .ZN(new_n1351));
  AND2_X1   g1151(.A1(new_n1344), .A2(new_n1346), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1321), .A2(new_n1323), .ZN(new_n1353));
  AOI21_X1  g1153(.A(KEYINPUT61), .B1(new_n1352), .B2(new_n1353), .ZN(new_n1354));
  INV_X1    g1154(.A(KEYINPUT63), .ZN(new_n1355));
  INV_X1    g1155(.A(new_n1337), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1355), .B1(new_n1353), .B2(new_n1356), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1340), .A2(KEYINPUT63), .A3(new_n1337), .ZN(new_n1358));
  NAND4_X1  g1158(.A1(new_n1354), .A2(new_n1314), .A3(new_n1357), .A4(new_n1358), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1351), .A2(new_n1359), .ZN(G405));
  XNOR2_X1  g1160(.A(new_n1314), .B(new_n1337), .ZN(new_n1361));
  AOI21_X1  g1161(.A(G378), .B1(new_n1270), .B2(new_n1272), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1269), .A2(G378), .ZN(new_n1363));
  INV_X1    g1163(.A(new_n1363), .ZN(new_n1364));
  OAI21_X1  g1164(.A(new_n1361), .B1(new_n1362), .B2(new_n1364), .ZN(new_n1365));
  XNOR2_X1  g1165(.A(new_n1314), .B(new_n1356), .ZN(new_n1366));
  NAND3_X1  g1166(.A1(new_n1366), .A2(new_n1307), .A3(new_n1363), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1365), .A2(new_n1367), .ZN(G402));
endmodule


