//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0 1 0 1 0 0 1 1 0 0 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n565, new_n567, new_n568, new_n569, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n581, new_n582,
    new_n583, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n620, new_n621, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT67), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G221), .A3(G219), .A4(G218), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  XOR2_X1   g032(.A(G325), .B(KEYINPUT69), .Z(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT70), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n463), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n465), .A2(new_n467), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n466), .A2(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(new_n469), .A3(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n468), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n468), .A2(G2104), .ZN(new_n477));
  INV_X1    g052(.A(G101), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR3_X1   g054(.A1(new_n472), .A2(new_n476), .A3(new_n479), .ZN(G160));
  NAND4_X1  g055(.A1(new_n465), .A2(new_n467), .A3(G2105), .A4(new_n469), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(KEYINPUT71), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT71), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT72), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n488), .B(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n470), .ZN(new_n491));
  NOR2_X1   g066(.A1(G100), .A2(G2105), .ZN(new_n492));
  XNOR2_X1  g067(.A(new_n492), .B(KEYINPUT73), .ZN(new_n493));
  INV_X1    g068(.A(G112), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n464), .B1(new_n494), .B2(G2105), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n491), .A2(G136), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n490), .A2(new_n496), .ZN(G162));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n465), .A2(new_n467), .A3(new_n499), .A4(new_n469), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n473), .A2(new_n469), .ZN(new_n501));
  NOR3_X1   g076(.A1(new_n498), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n500), .A2(KEYINPUT4), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n505), .B1(G114), .B2(new_n468), .ZN(new_n506));
  INV_X1    g081(.A(G126), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n506), .B1(new_n481), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n503), .A2(new_n508), .ZN(G164));
  AND2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT74), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT74), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G651), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n514), .A2(new_n516), .A3(KEYINPUT6), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT75), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n518), .B1(new_n519), .B2(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT74), .B(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n522), .A2(new_n518), .A3(KEYINPUT6), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n512), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G88), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n521), .A2(new_n523), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n526), .A2(G50), .A3(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(G75), .A2(G543), .ZN(new_n528));
  INV_X1    g103(.A(G62), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n528), .B1(new_n512), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n522), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n525), .A2(new_n527), .A3(new_n532), .ZN(G303));
  INV_X1    g108(.A(G303), .ZN(G166));
  INV_X1    g109(.A(G51), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n526), .A2(G543), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(KEYINPUT76), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT76), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n526), .A2(new_n538), .A3(G543), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n535), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT7), .ZN(new_n542));
  INV_X1    g117(.A(new_n512), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n543), .A2(G63), .A3(G651), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n526), .A2(new_n543), .ZN(new_n545));
  INV_X1    g120(.A(G89), .ZN(new_n546));
  OAI211_X1 g121(.A(new_n542), .B(new_n544), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n540), .A2(new_n547), .ZN(G168));
  AOI22_X1  g123(.A1(new_n543), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(new_n522), .ZN(new_n550));
  INV_X1    g125(.A(G90), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n545), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n537), .A2(new_n539), .ZN(new_n553));
  XOR2_X1   g128(.A(KEYINPUT77), .B(G52), .Z(new_n554));
  AOI21_X1  g129(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(G171));
  NAND2_X1  g130(.A1(new_n553), .A2(G43), .ZN(new_n556));
  XNOR2_X1  g131(.A(KEYINPUT78), .B(G81), .ZN(new_n557));
  NAND2_X1  g132(.A1(G68), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G56), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n512), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n524), .A2(new_n557), .B1(new_n531), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n565));
  XOR2_X1   g140(.A(new_n565), .B(KEYINPUT79), .Z(G176));
  XOR2_X1   g141(.A(KEYINPUT80), .B(KEYINPUT8), .Z(new_n567));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NAND4_X1  g144(.A1(G319), .A2(G483), .A3(G661), .A4(new_n569), .ZN(G188));
  NAND2_X1  g145(.A1(G53), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n526), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT9), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G65), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n512), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n524), .A2(G91), .B1(G651), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n574), .A2(new_n578), .ZN(G299));
  INV_X1    g154(.A(G171), .ZN(G301));
  OR3_X1    g155(.A1(new_n540), .A2(KEYINPUT81), .A3(new_n547), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT81), .B1(new_n540), .B2(new_n547), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G286));
  OR2_X1    g159(.A1(new_n543), .A2(G74), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n524), .A2(G87), .B1(new_n585), .B2(G651), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n526), .A2(G49), .A3(G543), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G288));
  NAND2_X1  g163(.A1(new_n524), .A2(G86), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n526), .A2(G48), .A3(G543), .ZN(new_n590));
  AND2_X1   g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n543), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n522), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT82), .ZN(G305));
  NAND2_X1  g171(.A1(new_n553), .A2(G47), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n543), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT83), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n522), .B1(new_n598), .B2(new_n599), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n600), .A2(new_n601), .B1(new_n524), .B2(G85), .ZN(new_n602));
  AND2_X1   g177(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(new_n553), .A2(G54), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n543), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n606), .A2(new_n513), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  INV_X1    g183(.A(G92), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n545), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n524), .A2(KEYINPUT10), .A3(G92), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n605), .A2(new_n607), .A3(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(new_n614), .B2(G171), .ZN(G321));
  XOR2_X1   g191(.A(G321), .B(KEYINPUT84), .Z(G284));
  MUX2_X1   g192(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g193(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g194(.A(new_n613), .ZN(new_n620));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(G860), .ZN(G148));
  NOR2_X1   g197(.A1(new_n613), .A2(G559), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT85), .ZN(new_n624));
  MUX2_X1   g199(.A(new_n562), .B(new_n624), .S(G868), .Z(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g201(.A1(new_n473), .A2(new_n469), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n627), .A2(new_n477), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT13), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT87), .ZN(new_n632));
  INV_X1    g207(.A(G2100), .ZN(new_n633));
  OAI22_X1  g208(.A1(new_n630), .A2(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n634), .B1(new_n631), .B2(new_n630), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n632), .A2(new_n633), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n487), .A2(G123), .ZN(new_n638));
  INV_X1    g213(.A(G2096), .ZN(new_n639));
  OAI21_X1  g214(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n640));
  INV_X1    g215(.A(G111), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n640), .B1(new_n641), .B2(G2105), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(new_n491), .B2(G135), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n638), .A2(new_n639), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n638), .A2(new_n643), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(G2096), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n637), .A2(new_n644), .A3(new_n646), .ZN(G156));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2427), .B(G2430), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT14), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT88), .Z(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n649), .B2(new_n650), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2451), .B(G2454), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT89), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n658), .A2(new_n661), .ZN(new_n663));
  AND3_X1   g238(.A1(new_n662), .A2(G14), .A3(new_n663), .ZN(G401));
  INV_X1    g239(.A(KEYINPUT18), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(KEYINPUT17), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n666), .A2(new_n667), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n665), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(new_n633), .ZN(new_n672));
  XOR2_X1   g247(.A(G2072), .B(G2078), .Z(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n668), .B2(KEYINPUT18), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(new_n639), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n672), .B(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1956), .B(G2474), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1961), .B(G1966), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  NOR3_X1   g257(.A1(new_n678), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n678), .A2(new_n681), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT20), .Z(new_n685));
  AOI211_X1 g260(.A(new_n683), .B(new_n685), .C1(new_n678), .C2(new_n682), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT90), .ZN(new_n687));
  XOR2_X1   g262(.A(G1981), .B(G1986), .Z(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n687), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(G229));
  NOR2_X1   g269(.A1(G29), .A2(G35), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(G162), .B2(G29), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT100), .B(KEYINPUT29), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g275(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT26), .Z(new_n702));
  INV_X1    g277(.A(G105), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(new_n477), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(G141), .B2(new_n491), .ZN(new_n705));
  INV_X1    g280(.A(G129), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(new_n486), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT97), .ZN(new_n708));
  MUX2_X1   g283(.A(G32), .B(new_n708), .S(G29), .Z(new_n709));
  XOR2_X1   g284(.A(KEYINPUT27), .B(G1996), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G5), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G171), .B2(new_n712), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n714), .A2(G1961), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT24), .B(G34), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT96), .Z(new_n719));
  INV_X1    g294(.A(G160), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(new_n717), .ZN(new_n721));
  INV_X1    g296(.A(G2084), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AND3_X1   g298(.A1(new_n711), .A2(new_n715), .A3(new_n723), .ZN(new_n724));
  OAI22_X1  g299(.A1(new_n700), .A2(G2090), .B1(new_n724), .B2(KEYINPUT99), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n563), .A2(G16), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G16), .B2(G19), .ZN(new_n727));
  INV_X1    g302(.A(G1341), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G1966), .ZN(new_n730));
  NOR2_X1   g305(.A1(G168), .A2(new_n712), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n712), .B2(G21), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n729), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n727), .A2(new_n728), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT30), .B(G28), .ZN(new_n735));
  OR2_X1    g310(.A1(KEYINPUT31), .A2(G11), .ZN(new_n736));
  NAND2_X1  g311(.A1(KEYINPUT31), .A2(G11), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n735), .A2(new_n717), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n645), .B2(new_n717), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT98), .ZN(new_n740));
  NOR3_X1   g315(.A1(new_n733), .A2(new_n734), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n721), .A2(new_n722), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT25), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n501), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n745), .A2(new_n468), .ZN(new_n746));
  AOI211_X1 g321(.A(new_n744), .B(new_n746), .C1(G139), .C2(new_n491), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n747), .A2(new_n717), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n717), .B2(G33), .ZN(new_n749));
  INV_X1    g324(.A(G2072), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n742), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n717), .A2(G27), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G164), .B2(new_n717), .ZN(new_n753));
  INV_X1    g328(.A(G2078), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n751), .B(new_n755), .C1(new_n750), .C2(new_n749), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n730), .B2(new_n732), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n709), .A2(new_n710), .ZN(new_n758));
  NOR2_X1   g333(.A1(G4), .A2(G16), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n620), .B2(G16), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n760), .A2(G1348), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n760), .A2(G1348), .ZN(new_n762));
  NOR3_X1   g337(.A1(new_n758), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n712), .A2(G20), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT23), .Z(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G299), .B2(G16), .ZN(new_n766));
  INV_X1    g341(.A(G1956), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G1961), .B2(new_n714), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n741), .A2(new_n757), .A3(new_n763), .A4(new_n769), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n698), .A2(G2090), .A3(new_n699), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n491), .A2(G140), .ZN(new_n772));
  NOR2_X1   g347(.A1(G104), .A2(G2105), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT93), .Z(new_n774));
  OAI21_X1  g349(.A(G2104), .B1(new_n468), .B2(G116), .ZN(new_n775));
  INV_X1    g350(.A(G128), .ZN(new_n776));
  OAI221_X1 g351(.A(new_n772), .B1(new_n774), .B2(new_n775), .C1(new_n486), .C2(new_n776), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT94), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(G29), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT95), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n717), .A2(G26), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT28), .ZN(new_n782));
  AND3_X1   g357(.A1(new_n779), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n780), .B1(new_n779), .B2(new_n782), .ZN(new_n784));
  INV_X1    g359(.A(G2067), .ZN(new_n785));
  OR3_X1    g360(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(new_n783), .B2(new_n784), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n711), .A2(KEYINPUT99), .A3(new_n715), .A4(new_n723), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n771), .A2(new_n786), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  NOR3_X1   g364(.A1(new_n725), .A2(new_n770), .A3(new_n789), .ZN(new_n790));
  MUX2_X1   g365(.A(G6), .B(G305), .S(G16), .Z(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT32), .B(G1981), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n712), .A2(G23), .ZN(new_n794));
  INV_X1    g369(.A(G288), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(new_n712), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT33), .B(G1976), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n712), .A2(G22), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT91), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G303), .B2(G16), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G1971), .ZN(new_n802));
  AND2_X1   g377(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n791), .A2(new_n792), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n793), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n805), .A2(KEYINPUT34), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT34), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n793), .A2(new_n803), .A3(new_n807), .A4(new_n804), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n712), .A2(G24), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n603), .B2(new_n712), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1986), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n717), .A2(G25), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n487), .A2(G119), .ZN(new_n813));
  OAI21_X1  g388(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n814));
  INV_X1    g389(.A(G107), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n814), .B1(new_n815), .B2(G2105), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(new_n491), .B2(G131), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n812), .B1(new_n819), .B2(new_n717), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT35), .B(G1991), .Z(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n820), .B(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n811), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n806), .A2(new_n808), .A3(new_n824), .ZN(new_n825));
  AND2_X1   g400(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n826));
  NOR2_X1   g401(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n806), .A2(new_n826), .A3(new_n808), .A4(new_n824), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n790), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(G311));
  XNOR2_X1  g407(.A(new_n831), .B(KEYINPUT101), .ZN(G150));
  NAND2_X1  g408(.A1(new_n553), .A2(G55), .ZN(new_n834));
  NAND2_X1  g409(.A1(G80), .A2(G543), .ZN(new_n835));
  INV_X1    g410(.A(G67), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n835), .B1(new_n512), .B2(new_n836), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n524), .A2(G93), .B1(new_n531), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(KEYINPUT103), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT103), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n834), .A2(new_n841), .A3(new_n838), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  XOR2_X1   g419(.A(KEYINPUT104), .B(G860), .Z(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(KEYINPUT106), .B(KEYINPUT37), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n613), .A2(new_n621), .ZN(new_n849));
  XNOR2_X1  g424(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n563), .B1(new_n840), .B2(new_n842), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n839), .A2(new_n562), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n851), .B(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT39), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT105), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n856), .A2(new_n857), .A3(new_n845), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n857), .B1(new_n856), .B2(new_n845), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n848), .B1(new_n858), .B2(new_n859), .ZN(G145));
  XNOR2_X1  g435(.A(new_n645), .B(G160), .ZN(new_n861));
  XNOR2_X1  g436(.A(G162), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n818), .B(new_n630), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n491), .A2(G142), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT107), .Z(new_n865));
  NAND2_X1  g440(.A1(new_n487), .A2(G130), .ZN(new_n866));
  OR2_X1    g441(.A1(G106), .A2(G2105), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n867), .B(G2104), .C1(G118), .C2(new_n468), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n865), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n863), .B(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(G164), .ZN(new_n871));
  AND2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n870), .A2(new_n871), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n778), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n870), .A2(new_n871), .ZN(new_n875));
  INV_X1    g450(.A(new_n778), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n870), .A2(new_n871), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n747), .A2(new_n707), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n879), .B1(new_n708), .B2(new_n747), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n874), .A2(new_n878), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n881), .B1(new_n874), .B2(new_n878), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n862), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NOR3_X1   g459(.A1(new_n872), .A2(new_n873), .A3(new_n778), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n876), .B1(new_n875), .B2(new_n877), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n880), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n862), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n874), .A2(new_n878), .A3(new_n881), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(G37), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n884), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g468(.A(G305), .B(new_n603), .ZN(new_n894));
  XNOR2_X1  g469(.A(G288), .B(G303), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT42), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT42), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(new_n896), .B2(new_n897), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(KEYINPUT108), .A3(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n624), .B(new_n854), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n613), .A2(G299), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n613), .A2(G299), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n906), .B(KEYINPUT41), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n903), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n902), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT108), .B1(new_n899), .B2(new_n901), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n910), .A2(new_n614), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n902), .A2(new_n907), .A3(new_n909), .ZN(new_n913));
  AOI22_X1  g488(.A1(new_n912), .A2(new_n913), .B1(new_n614), .B2(new_n844), .ZN(G295));
  AOI22_X1  g489(.A1(new_n912), .A2(new_n913), .B1(new_n614), .B2(new_n844), .ZN(G331));
  INV_X1    g490(.A(KEYINPUT109), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n583), .A2(G171), .ZN(new_n917));
  INV_X1    g492(.A(G168), .ZN(new_n918));
  NAND2_X1  g493(.A1(G301), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n854), .A2(new_n920), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n917), .B(new_n919), .C1(new_n852), .C2(new_n853), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n908), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n906), .B1(new_n921), .B2(new_n922), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n916), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n921), .A2(new_n922), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n904), .A2(new_n905), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n923), .A2(new_n929), .A3(KEYINPUT109), .ZN(new_n930));
  INV_X1    g505(.A(new_n898), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n926), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n898), .A2(new_n929), .A3(new_n923), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n933), .A2(new_n891), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT43), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n931), .B1(new_n924), .B2(new_n925), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n934), .A2(KEYINPUT43), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT44), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n940), .B1(new_n932), .B2(new_n934), .ZN(new_n941));
  AND4_X1   g516(.A1(new_n940), .A2(new_n936), .A3(new_n933), .A4(new_n891), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n938), .A2(new_n943), .ZN(G397));
  INV_X1    g519(.A(G1384), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(new_n503), .B2(new_n508), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT45), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n476), .A2(new_n479), .ZN(new_n949));
  INV_X1    g524(.A(new_n472), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(new_n950), .A3(G40), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n778), .B(G2067), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n952), .B1(new_n953), .B2(new_n707), .ZN(new_n954));
  INV_X1    g529(.A(G1996), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n956), .B(KEYINPUT46), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(KEYINPUT47), .ZN(new_n959));
  INV_X1    g534(.A(new_n952), .ZN(new_n960));
  NOR3_X1   g535(.A1(G290), .A2(G1986), .A3(new_n960), .ZN(new_n961));
  XOR2_X1   g536(.A(new_n961), .B(KEYINPUT48), .Z(new_n962));
  NAND2_X1  g537(.A1(new_n707), .A2(G1996), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n963), .B1(new_n708), .B2(G1996), .ZN(new_n964));
  OR2_X1    g539(.A1(new_n953), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n818), .B(new_n822), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n962), .B1(new_n967), .B2(new_n960), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n819), .A2(new_n821), .ZN(new_n969));
  OAI22_X1  g544(.A1(new_n965), .A2(new_n969), .B1(G2067), .B2(new_n778), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n952), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n959), .A2(new_n968), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n948), .A2(KEYINPUT110), .ZN(new_n974));
  INV_X1    g549(.A(G40), .ZN(new_n975));
  NOR4_X1   g550(.A1(new_n472), .A2(new_n476), .A3(new_n975), .A4(new_n479), .ZN(new_n976));
  OAI211_X1 g551(.A(KEYINPUT45), .B(new_n945), .C1(new_n503), .C2(new_n508), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT110), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n946), .A2(new_n979), .A3(new_n947), .ZN(new_n980));
  XNOR2_X1  g555(.A(KEYINPUT56), .B(G2072), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n974), .A2(new_n978), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT116), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT57), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n573), .A2(KEYINPUT9), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT9), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n526), .B2(new_n572), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n578), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n983), .B(new_n986), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n976), .B1(new_n946), .B2(KEYINPUT50), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n946), .A2(KEYINPUT50), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n767), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n574), .A2(new_n984), .A3(new_n985), .A4(new_n578), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n982), .A2(new_n992), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n982), .A2(new_n995), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n998), .A2(KEYINPUT117), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n998), .A2(KEYINPUT117), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n992), .A2(new_n996), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G114), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n504), .B1(new_n1004), .B2(G2105), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1005), .B1(new_n482), .B2(G126), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n501), .A2(new_n502), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(G1384), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT50), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n951), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n946), .A2(new_n1013), .A3(KEYINPUT50), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1013), .B1(new_n946), .B2(KEYINPUT50), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1012), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G1348), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n951), .A2(new_n946), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n1016), .A2(new_n1017), .B1(new_n785), .B2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1019), .A2(new_n613), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n997), .B1(new_n1003), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n998), .A2(new_n1001), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n997), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT61), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n613), .A2(KEYINPUT60), .ZN(new_n1025));
  AOI22_X1  g600(.A1(new_n1023), .A2(new_n1024), .B1(new_n1019), .B2(new_n1025), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n1019), .A2(new_n613), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT60), .B1(new_n1027), .B2(new_n1020), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT59), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n974), .A2(new_n978), .A3(new_n955), .A4(new_n980), .ZN(new_n1030));
  XOR2_X1   g605(.A(KEYINPUT58), .B(G1341), .Z(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(new_n951), .B2(new_n946), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g608(.A(KEYINPUT118), .B(new_n1029), .C1(new_n1033), .C2(new_n562), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT118), .B1(new_n1033), .B2(new_n562), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n562), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1029), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1026), .A2(new_n1028), .A3(new_n1034), .A4(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT119), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1024), .B1(new_n997), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1042), .B1(new_n1041), .B2(new_n997), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1043), .A2(new_n1003), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1021), .B1(new_n1040), .B2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1012), .B(new_n722), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n948), .A2(new_n977), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n730), .B1(new_n1047), .B2(new_n951), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(G8), .ZN(new_n1050));
  OAI21_X1  g625(.A(G8), .B1(new_n540), .B2(new_n547), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT51), .B1(new_n1051), .B2(KEYINPUT120), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1050), .A2(new_n1053), .A3(new_n1051), .ZN(new_n1054));
  OAI211_X1 g629(.A(G8), .B(new_n1052), .C1(new_n1049), .C2(new_n918), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1049), .A2(G8), .A3(new_n918), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT112), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n1060));
  INV_X1    g635(.A(G8), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1060), .B1(G166), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT112), .ZN(new_n1063));
  NAND4_X1  g638(.A1(G303), .A2(new_n1063), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1059), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n974), .A2(new_n978), .A3(new_n980), .ZN(new_n1066));
  INV_X1    g641(.A(G1971), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n993), .A2(new_n994), .ZN(new_n1068));
  INV_X1    g643(.A(G2090), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1066), .A2(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1065), .B1(new_n1070), .B2(new_n1061), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1059), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1012), .B(new_n1069), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n979), .B1(new_n946), .B2(new_n947), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n976), .A2(new_n977), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(G1971), .B1(new_n1077), .B2(new_n980), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1072), .B(G8), .C1(new_n1074), .C2(new_n1078), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1071), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT49), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n589), .A2(new_n590), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT114), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n589), .A2(new_n1084), .A3(new_n590), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1083), .A2(new_n594), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1086), .A2(new_n1087), .A3(G1981), .ZN(new_n1088));
  INV_X1    g663(.A(G1981), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n591), .A2(new_n1089), .A3(new_n594), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1087), .B1(new_n1086), .B2(G1981), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1081), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n589), .A2(new_n1084), .A3(new_n590), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1084), .B1(new_n589), .B2(new_n590), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n1094), .A2(new_n1095), .A3(new_n593), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT115), .B1(new_n1096), .B2(new_n1089), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1097), .A2(KEYINPUT49), .A3(new_n1090), .A4(new_n1088), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1018), .A2(new_n1061), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1093), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G1976), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1099), .B1(G288), .B2(new_n1101), .ZN(new_n1102));
  AND2_X1   g677(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1102), .B(new_n1103), .ZN(new_n1104));
  OR3_X1    g679(.A1(new_n795), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1057), .A2(new_n1080), .A3(new_n1100), .A4(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n974), .A2(new_n978), .A3(new_n754), .A4(new_n980), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT53), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G1961), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1016), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1047), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n1114));
  AOI211_X1 g689(.A(new_n1109), .B(G2078), .C1(new_n951), .C2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(G160), .A2(KEYINPUT122), .A3(G40), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1113), .A2(new_n1115), .A3(KEYINPUT123), .A4(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT123), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n951), .A2(new_n1114), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1109), .A2(G2078), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1119), .A2(new_n1116), .A3(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1118), .B1(new_n1121), .B2(new_n1047), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1110), .A2(new_n1112), .A3(new_n1117), .A4(new_n1122), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1123), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT125), .B1(new_n1123), .B2(G171), .ZN(new_n1125));
  AND4_X1   g700(.A1(new_n948), .A2(new_n976), .A3(new_n977), .A4(new_n1120), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1126), .B1(new_n1016), .B2(new_n1111), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n1110), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT54), .B1(new_n1128), .B2(G171), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1124), .A2(new_n1125), .A3(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1107), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT124), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT54), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1134), .B1(new_n1128), .B2(G171), .ZN(new_n1135));
  AOI211_X1 g710(.A(KEYINPUT121), .B(G301), .C1(new_n1127), .C2(new_n1110), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1123), .A2(G171), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1132), .B(new_n1133), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1135), .A2(new_n1138), .A3(new_n1136), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT124), .B1(new_n1140), .B2(KEYINPUT54), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1045), .A2(new_n1131), .A3(new_n1139), .A4(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT126), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1100), .A2(new_n1106), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1074), .A2(new_n1078), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1065), .B1(new_n1145), .B2(new_n1061), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1050), .A2(G286), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(KEYINPUT63), .B1(new_n1144), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n795), .A2(new_n1101), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1099), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1097), .A2(new_n1090), .A3(new_n1088), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1151), .B1(new_n1152), .B2(new_n1081), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1150), .B1(new_n1153), .B2(new_n1098), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1090), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1099), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT63), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1147), .A2(new_n1071), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n1079), .ZN(new_n1159));
  AOI22_X1  g734(.A1(new_n1153), .A2(new_n1098), .B1(new_n1105), .B2(new_n1104), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1149), .A2(new_n1156), .A3(new_n1161), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n1142), .A2(new_n1143), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1143), .B1(new_n1142), .B2(new_n1162), .ZN(new_n1164));
  XOR2_X1   g739(.A(new_n1057), .B(KEYINPUT62), .Z(new_n1165));
  AND4_X1   g740(.A1(new_n1137), .A2(new_n1165), .A3(new_n1160), .A4(new_n1080), .ZN(new_n1166));
  NOR3_X1   g741(.A1(new_n1163), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n603), .B(G1986), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n960), .B1(new_n967), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n973), .B1(new_n1167), .B2(new_n1169), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g745(.A1(new_n461), .A2(G227), .ZN(new_n1172));
  OR2_X1    g746(.A1(new_n1172), .A2(KEYINPUT127), .ZN(new_n1173));
  NAND2_X1  g747(.A1(new_n1172), .A2(KEYINPUT127), .ZN(new_n1174));
  NAND3_X1  g748(.A1(new_n693), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  NOR2_X1   g749(.A1(G401), .A2(new_n1175), .ZN(new_n1176));
  OAI211_X1 g750(.A(new_n892), .B(new_n1176), .C1(new_n941), .C2(new_n942), .ZN(G225));
  INV_X1    g751(.A(G225), .ZN(G308));
endmodule


