

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757;

  XNOR2_X1 U368 ( .A(n442), .B(KEYINPUT108), .ZN(n756) );
  NOR2_X2 U369 ( .A1(n624), .A2(n625), .ZN(n434) );
  OR2_X2 U370 ( .A1(n722), .A2(G902), .ZN(n468) );
  NOR2_X2 U371 ( .A1(n677), .A2(n680), .ZN(n619) );
  XNOR2_X2 U372 ( .A(n440), .B(n348), .ZN(n584) );
  OR2_X2 U373 ( .A1(n718), .A2(G902), .ZN(n440) );
  XNOR2_X2 U374 ( .A(n534), .B(n730), .ZN(n536) );
  XNOR2_X2 U375 ( .A(n741), .B(n500), .ZN(n534) );
  INV_X1 U376 ( .A(n598), .ZN(n689) );
  INV_X1 U377 ( .A(G125), .ZN(n444) );
  NOR2_X1 U378 ( .A1(n754), .A2(n755), .ZN(n583) );
  XNOR2_X1 U379 ( .A(n570), .B(KEYINPUT99), .ZN(n660) );
  OR2_X2 U380 ( .A1(n569), .A2(n585), .ZN(n406) );
  AND2_X2 U381 ( .A1(n646), .A2(n647), .ZN(n720) );
  NAND2_X1 U382 ( .A1(n710), .A2(n639), .ZN(n647) );
  AND2_X1 U383 ( .A1(n371), .A2(n515), .ZN(n646) );
  AND2_X1 U384 ( .A1(n453), .A2(n452), .ZN(n451) );
  XNOR2_X1 U385 ( .A(n627), .B(KEYINPUT110), .ZN(n383) );
  XNOR2_X1 U386 ( .A(n433), .B(n621), .ZN(n757) );
  NAND2_X1 U387 ( .A1(n403), .A2(n401), .ZN(n627) );
  AND2_X1 U388 ( .A1(n398), .A2(n405), .ZN(n403) );
  AND2_X1 U389 ( .A1(n443), .A2(n485), .ZN(n409) );
  AND2_X1 U390 ( .A1(n612), .A2(n486), .ZN(n485) );
  NOR2_X2 U391 ( .A1(n660), .A2(n663), .ZN(n679) );
  XNOR2_X1 U392 ( .A(n619), .B(n618), .ZN(n375) );
  INV_X1 U393 ( .A(n599), .ZN(n347) );
  XNOR2_X1 U394 ( .A(n633), .B(KEYINPUT38), .ZN(n376) );
  XNOR2_X1 U395 ( .A(n584), .B(KEYINPUT97), .ZN(n569) );
  XOR2_X1 U396 ( .A(G478), .B(n554), .Z(n585) );
  XNOR2_X1 U397 ( .A(n415), .B(G116), .ZN(n548) );
  XNOR2_X1 U398 ( .A(n737), .B(G146), .ZN(n540) );
  INV_X1 U399 ( .A(KEYINPUT41), .ZN(n618) );
  INV_X2 U400 ( .A(G953), .ZN(n746) );
  XNOR2_X1 U401 ( .A(G131), .B(G134), .ZN(n737) );
  INV_X1 U402 ( .A(G143), .ZN(n445) );
  XNOR2_X2 U403 ( .A(n524), .B(n523), .ZN(n558) );
  XNOR2_X2 U404 ( .A(n444), .B(G146), .ZN(n524) );
  XNOR2_X2 U405 ( .A(n580), .B(n579), .ZN(n609) );
  XNOR2_X2 U406 ( .A(n411), .B(KEYINPUT45), .ZN(n724) );
  INV_X1 U407 ( .A(KEYINPUT10), .ZN(n523) );
  AND2_X1 U408 ( .A1(n459), .A2(n347), .ZN(n587) );
  XNOR2_X1 U409 ( .A(n586), .B(KEYINPUT104), .ZN(n459) );
  NAND2_X1 U410 ( .A1(n689), .A2(n688), .ZN(n685) );
  XNOR2_X1 U411 ( .A(n372), .B(n422), .ZN(n574) );
  INV_X1 U412 ( .A(KEYINPUT0), .ZN(n422) );
  XNOR2_X1 U413 ( .A(n489), .B(n488), .ZN(n487) );
  NAND2_X1 U414 ( .A1(n562), .A2(G210), .ZN(n488) );
  XNOR2_X1 U415 ( .A(n540), .B(n539), .ZN(n489) );
  XNOR2_X1 U416 ( .A(n368), .B(n552), .ZN(n719) );
  XNOR2_X1 U417 ( .A(n547), .B(n393), .ZN(n552) );
  XNOR2_X1 U418 ( .A(n551), .B(n553), .ZN(n368) );
  XNOR2_X1 U419 ( .A(n386), .B(n432), .ZN(n393) );
  XNOR2_X1 U420 ( .A(KEYINPUT65), .B(G101), .ZN(n500) );
  XNOR2_X1 U421 ( .A(n417), .B(n416), .ZN(n530) );
  XNOR2_X1 U422 ( .A(G104), .B(G107), .ZN(n416) );
  XNOR2_X1 U423 ( .A(n364), .B(G110), .ZN(n417) );
  INV_X1 U424 ( .A(KEYINPUT70), .ZN(n364) );
  XNOR2_X1 U425 ( .A(n622), .B(KEYINPUT39), .ZN(n637) );
  AND2_X1 U426 ( .A1(n485), .A2(n376), .ZN(n410) );
  INV_X1 U427 ( .A(KEYINPUT81), .ZN(n450) );
  NAND2_X1 U428 ( .A1(n638), .A2(KEYINPUT81), .ZN(n452) );
  NOR2_X1 U429 ( .A1(n589), .A2(n752), .ZN(n413) );
  XNOR2_X1 U430 ( .A(n545), .B(KEYINPUT92), .ZN(n365) );
  INV_X1 U431 ( .A(KEYINPUT18), .ZN(n495) );
  XNOR2_X1 U432 ( .A(n524), .B(n498), .ZN(n439) );
  XNOR2_X1 U433 ( .A(n370), .B(n369), .ZN(n635) );
  INV_X1 U434 ( .A(KEYINPUT48), .ZN(n369) );
  XNOR2_X1 U435 ( .A(n467), .B(KEYINPUT66), .ZN(n604) );
  NAND2_X1 U436 ( .A1(n598), .A2(n597), .ZN(n467) );
  NOR2_X1 U437 ( .A1(n686), .A2(n685), .ZN(n586) );
  XNOR2_X1 U438 ( .A(G113), .B(KEYINPUT3), .ZN(n501) );
  XNOR2_X1 U439 ( .A(n568), .B(n567), .ZN(n718) );
  XNOR2_X1 U440 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U441 ( .A(n395), .B(n561), .ZN(n568) );
  NOR2_X1 U442 ( .A1(n381), .A2(n686), .ZN(n380) );
  NOR2_X1 U443 ( .A1(n466), .A2(n465), .ZN(n381) );
  INV_X1 U444 ( .A(n633), .ZN(n474) );
  INV_X1 U445 ( .A(n611), .ZN(n486) );
  NAND2_X1 U446 ( .A1(n609), .A2(n675), .ZN(n484) );
  NOR2_X1 U447 ( .A1(G902), .A2(n719), .ZN(n554) );
  AND2_X1 U448 ( .A1(n392), .A2(n391), .ZN(n390) );
  NAND2_X1 U449 ( .A1(n541), .A2(n389), .ZN(n388) );
  XNOR2_X1 U450 ( .A(n575), .B(n374), .ZN(n373) );
  INV_X1 U451 ( .A(KEYINPUT22), .ZN(n374) );
  NAND2_X1 U452 ( .A1(n720), .A2(G472), .ZN(n651) );
  NAND2_X1 U453 ( .A1(n720), .A2(G478), .ZN(n427) );
  INV_X1 U454 ( .A(n719), .ZN(n430) );
  NAND2_X1 U455 ( .A1(n720), .A2(G475), .ZN(n493) );
  XNOR2_X1 U456 ( .A(n458), .B(n454), .ZN(n533) );
  XNOR2_X1 U457 ( .A(n457), .B(n455), .ZN(n454) );
  XNOR2_X1 U458 ( .A(n530), .B(n540), .ZN(n458) );
  AND2_X1 U459 ( .A1(n712), .A2(n356), .ZN(n714) );
  NAND2_X1 U460 ( .A1(G234), .A2(G237), .ZN(n508) );
  XOR2_X1 U461 ( .A(KEYINPUT69), .B(KEYINPUT14), .Z(n509) );
  NAND2_X1 U462 ( .A1(n604), .A2(KEYINPUT105), .ZN(n405) );
  NAND2_X1 U463 ( .A1(n474), .A2(n675), .ZN(n600) );
  XNOR2_X1 U464 ( .A(G116), .B(G137), .ZN(n537) );
  XNOR2_X1 U465 ( .A(n384), .B(KEYINPUT71), .ZN(n562) );
  NAND2_X1 U466 ( .A1(n746), .A2(n385), .ZN(n384) );
  INV_X1 U467 ( .A(G237), .ZN(n385) );
  INV_X1 U468 ( .A(G107), .ZN(n432) );
  XOR2_X1 U469 ( .A(G131), .B(G122), .Z(n564) );
  XNOR2_X1 U470 ( .A(G143), .B(G113), .ZN(n563) );
  XNOR2_X1 U471 ( .A(n558), .B(n557), .ZN(n395) );
  XNOR2_X1 U472 ( .A(G104), .B(G140), .ZN(n555) );
  XOR2_X1 U473 ( .A(KEYINPUT95), .B(KEYINPUT93), .Z(n556) );
  XNOR2_X1 U474 ( .A(KEYINPUT94), .B(KEYINPUT11), .ZN(n559) );
  XOR2_X1 U475 ( .A(KEYINPUT12), .B(KEYINPUT96), .Z(n560) );
  NAND2_X1 U476 ( .A1(n562), .A2(G214), .ZN(n566) );
  XNOR2_X1 U477 ( .A(KEYINPUT4), .B(KEYINPUT64), .ZN(n499) );
  XNOR2_X1 U478 ( .A(n456), .B(G140), .ZN(n531) );
  INV_X1 U479 ( .A(G137), .ZN(n456) );
  OR2_X1 U480 ( .A1(G902), .A2(G237), .ZN(n507) );
  NAND2_X1 U481 ( .A1(n376), .A2(n675), .ZN(n680) );
  INV_X1 U482 ( .A(n600), .ZN(n466) );
  XNOR2_X1 U483 ( .A(n600), .B(KEYINPUT19), .ZN(n607) );
  INV_X1 U484 ( .A(G902), .ZN(n389) );
  NAND2_X1 U485 ( .A1(n447), .A2(G902), .ZN(n391) );
  XNOR2_X1 U486 ( .A(n572), .B(n394), .ZN(n677) );
  INV_X1 U487 ( .A(KEYINPUT100), .ZN(n394) );
  NAND2_X1 U488 ( .A1(n448), .A2(n355), .ZN(n449) );
  INV_X1 U489 ( .A(G122), .ZN(n415) );
  XNOR2_X1 U490 ( .A(n462), .B(n461), .ZN(n460) );
  XNOR2_X1 U491 ( .A(KEYINPUT23), .B(KEYINPUT86), .ZN(n461) );
  XNOR2_X1 U492 ( .A(n463), .B(G110), .ZN(n462) );
  INV_X1 U493 ( .A(KEYINPUT85), .ZN(n463) );
  XNOR2_X1 U494 ( .A(n519), .B(n520), .ZN(n464) );
  XNOR2_X1 U495 ( .A(KEYINPUT24), .B(KEYINPUT67), .ZN(n520) );
  XNOR2_X1 U496 ( .A(n436), .B(n435), .ZN(n546) );
  INV_X1 U497 ( .A(KEYINPUT8), .ZN(n435) );
  NAND2_X1 U498 ( .A1(n746), .A2(G234), .ZN(n436) );
  XOR2_X1 U499 ( .A(G902), .B(KEYINPUT15), .Z(n515) );
  INV_X1 U500 ( .A(n531), .ZN(n455) );
  XNOR2_X1 U501 ( .A(n532), .B(KEYINPUT72), .ZN(n457) );
  XNOR2_X1 U502 ( .A(n497), .B(n439), .ZN(n473) );
  NOR2_X1 U503 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U504 ( .A(n397), .B(n396), .ZN(n605) );
  INV_X1 U505 ( .A(KEYINPUT28), .ZN(n396) );
  NOR2_X1 U506 ( .A1(n603), .A2(n604), .ZN(n397) );
  INV_X1 U507 ( .A(KEYINPUT6), .ZN(n446) );
  XNOR2_X1 U508 ( .A(n530), .B(n414), .ZN(n731) );
  XNOR2_X1 U509 ( .A(n548), .B(KEYINPUT16), .ZN(n414) );
  NAND2_X1 U510 ( .A1(n637), .A2(n663), .ZN(n623) );
  NAND2_X1 U511 ( .A1(n379), .A2(n377), .ZN(n601) );
  NAND2_X1 U512 ( .A1(n378), .A2(KEYINPUT36), .ZN(n377) );
  AND2_X1 U513 ( .A1(n382), .A2(n380), .ZN(n379) );
  XNOR2_X1 U514 ( .A(n469), .B(KEYINPUT35), .ZN(n752) );
  XNOR2_X1 U515 ( .A(n472), .B(n471), .ZN(n470) );
  INV_X1 U516 ( .A(KEYINPUT34), .ZN(n471) );
  XNOR2_X1 U517 ( .A(n419), .B(n418), .ZN(n755) );
  INV_X1 U518 ( .A(KEYINPUT32), .ZN(n418) );
  XNOR2_X1 U519 ( .A(n542), .B(n366), .ZN(n668) );
  XNOR2_X1 U520 ( .A(n367), .B(KEYINPUT91), .ZN(n366) );
  INV_X1 U521 ( .A(KEYINPUT31), .ZN(n367) );
  XNOR2_X1 U522 ( .A(n421), .B(n420), .ZN(n754) );
  INV_X1 U523 ( .A(KEYINPUT103), .ZN(n420) );
  AND2_X1 U524 ( .A1(n373), .A2(n358), .ZN(n421) );
  NAND2_X1 U525 ( .A1(n652), .A2(n428), .ZN(n653) );
  XNOR2_X1 U526 ( .A(n651), .B(n360), .ZN(n652) );
  XNOR2_X1 U527 ( .A(n722), .B(n721), .ZN(n479) );
  INV_X1 U528 ( .A(KEYINPUT122), .ZN(n423) );
  NAND2_X1 U529 ( .A1(n429), .A2(n428), .ZN(n424) );
  XNOR2_X1 U530 ( .A(n427), .B(n430), .ZN(n429) );
  INV_X1 U531 ( .A(KEYINPUT60), .ZN(n490) );
  NAND2_X1 U532 ( .A1(n492), .A2(n428), .ZN(n491) );
  XNOR2_X1 U533 ( .A(n493), .B(n361), .ZN(n492) );
  XNOR2_X1 U534 ( .A(n717), .B(n716), .ZN(n476) );
  INV_X1 U535 ( .A(KEYINPUT56), .ZN(n425) );
  INV_X1 U536 ( .A(KEYINPUT53), .ZN(n437) );
  XOR2_X1 U537 ( .A(KEYINPUT13), .B(G475), .Z(n348) );
  AND2_X1 U538 ( .A1(G210), .A2(n507), .ZN(n349) );
  AND2_X1 U539 ( .A1(n373), .A2(n686), .ZN(n350) );
  AND2_X1 U540 ( .A1(n608), .A2(n664), .ZN(n351) );
  INV_X1 U541 ( .A(n541), .ZN(n447) );
  NOR2_X1 U542 ( .A1(n689), .A2(n609), .ZN(n352) );
  AND2_X1 U543 ( .A1(n585), .A2(n584), .ZN(n353) );
  AND2_X1 U544 ( .A1(n708), .A2(n375), .ZN(n354) );
  AND2_X1 U545 ( .A1(n673), .A2(n450), .ZN(n355) );
  NOR2_X1 U546 ( .A1(n713), .A2(n354), .ZN(n356) );
  AND2_X1 U547 ( .A1(n466), .A2(n465), .ZN(n357) );
  AND2_X1 U548 ( .A1(n686), .A2(n352), .ZN(n358) );
  XNOR2_X1 U549 ( .A(KEYINPUT74), .B(n582), .ZN(n359) );
  INV_X1 U550 ( .A(KEYINPUT36), .ZN(n465) );
  INV_X1 U551 ( .A(KEYINPUT105), .ZN(n408) );
  XOR2_X1 U552 ( .A(n650), .B(KEYINPUT62), .Z(n360) );
  XOR2_X1 U553 ( .A(n718), .B(n494), .Z(n361) );
  XOR2_X1 U554 ( .A(n504), .B(n503), .Z(n362) );
  NOR2_X1 U555 ( .A1(G952), .A2(n746), .ZN(n723) );
  INV_X1 U556 ( .A(n723), .ZN(n428) );
  XNOR2_X1 U557 ( .A(n363), .B(KEYINPUT46), .ZN(n624) );
  NAND2_X1 U558 ( .A1(n482), .A2(n757), .ZN(n363) );
  NAND2_X1 U559 ( .A1(n412), .A2(n590), .ZN(n411) );
  NAND2_X1 U560 ( .A1(n679), .A2(KEYINPUT47), .ZN(n441) );
  OR2_X1 U561 ( .A1(n707), .A2(n588), .ZN(n472) );
  NAND2_X1 U562 ( .A1(n470), .A2(n353), .ZN(n469) );
  NAND2_X1 U563 ( .A1(n365), .A2(n571), .ZN(n578) );
  NAND2_X1 U564 ( .A1(n483), .A2(n409), .ZN(n442) );
  NAND2_X1 U565 ( .A1(n626), .A2(n434), .ZN(n370) );
  AND2_X1 U566 ( .A1(n353), .A2(n474), .ZN(n443) );
  NAND2_X1 U567 ( .A1(n644), .A2(n724), .ZN(n371) );
  NAND2_X1 U568 ( .A1(n711), .A2(n371), .ZN(n712) );
  NAND2_X1 U569 ( .A1(n607), .A2(n514), .ZN(n372) );
  NAND2_X1 U570 ( .A1(n373), .A2(n359), .ZN(n419) );
  NAND2_X1 U571 ( .A1(n620), .A2(n375), .ZN(n433) );
  NAND2_X1 U572 ( .A1(n699), .A2(n375), .ZN(n700) );
  NOR2_X1 U573 ( .A1(n376), .A2(n675), .ZN(n676) );
  INV_X1 U574 ( .A(n383), .ZN(n378) );
  NAND2_X1 U575 ( .A1(n383), .A2(n357), .ZN(n382) );
  XNOR2_X2 U576 ( .A(n386), .B(n499), .ZN(n741) );
  XNOR2_X2 U577 ( .A(n445), .B(G128), .ZN(n386) );
  NAND2_X4 U578 ( .A1(n390), .A2(n387), .ZN(n580) );
  OR2_X1 U579 ( .A1(n649), .A2(n388), .ZN(n387) );
  NAND2_X1 U580 ( .A1(n649), .A2(n447), .ZN(n392) );
  NOR2_X1 U581 ( .A1(n585), .A2(n584), .ZN(n572) );
  NOR2_X1 U582 ( .A1(n406), .A2(n400), .ZN(n402) );
  NAND2_X1 U583 ( .A1(n399), .A2(KEYINPUT105), .ZN(n398) );
  NAND2_X1 U584 ( .A1(n404), .A2(n347), .ZN(n399) );
  NAND2_X1 U585 ( .A1(n347), .A2(n408), .ZN(n400) );
  XNOR2_X2 U586 ( .A(n580), .B(n446), .ZN(n599) );
  NAND2_X1 U587 ( .A1(n402), .A2(n407), .ZN(n401) );
  INV_X1 U588 ( .A(n406), .ZN(n404) );
  INV_X1 U589 ( .A(n406), .ZN(n663) );
  INV_X1 U590 ( .A(n604), .ZN(n407) );
  NAND2_X1 U591 ( .A1(n483), .A2(n410), .ZN(n622) );
  XNOR2_X1 U592 ( .A(n413), .B(KEYINPUT44), .ZN(n412) );
  INV_X1 U593 ( .A(n574), .ZN(n588) );
  XNOR2_X1 U594 ( .A(n424), .B(n423), .ZN(G63) );
  XNOR2_X1 U595 ( .A(n426), .B(n425), .ZN(G51) );
  NAND2_X1 U596 ( .A1(n431), .A2(n428), .ZN(n426) );
  NAND2_X1 U597 ( .A1(n546), .A2(G217), .ZN(n547) );
  XNOR2_X1 U598 ( .A(n536), .B(n487), .ZN(n649) );
  XNOR2_X1 U599 ( .A(n648), .B(n362), .ZN(n431) );
  XNOR2_X1 U600 ( .A(n464), .B(n460), .ZN(n522) );
  NOR2_X2 U601 ( .A1(n606), .A2(n685), .ZN(n612) );
  XNOR2_X1 U602 ( .A(n438), .B(n437), .ZN(G75) );
  NAND2_X1 U603 ( .A1(n715), .A2(n746), .ZN(n438) );
  NAND2_X1 U604 ( .A1(n640), .A2(KEYINPUT81), .ZN(n453) );
  NAND2_X1 U605 ( .A1(n756), .A2(n441), .ZN(n613) );
  INV_X1 U606 ( .A(n640), .ZN(n448) );
  NAND2_X2 U607 ( .A1(n451), .A2(n449), .ZN(n481) );
  NAND2_X1 U608 ( .A1(n481), .A2(n724), .ZN(n710) );
  NOR2_X1 U609 ( .A1(n505), .A2(n515), .ZN(n506) );
  XNOR2_X1 U610 ( .A(n473), .B(n731), .ZN(n502) );
  XNOR2_X2 U611 ( .A(n606), .B(KEYINPUT1), .ZN(n686) );
  XNOR2_X2 U612 ( .A(n468), .B(n526), .ZN(n598) );
  XNOR2_X2 U613 ( .A(n506), .B(n349), .ZN(n633) );
  NOR2_X1 U614 ( .A1(n475), .A2(n723), .ZN(G54) );
  XNOR2_X1 U615 ( .A(n477), .B(n476), .ZN(n475) );
  NAND2_X1 U616 ( .A1(n720), .A2(G469), .ZN(n477) );
  NOR2_X1 U617 ( .A1(n478), .A2(n723), .ZN(G66) );
  XNOR2_X1 U618 ( .A(n480), .B(n479), .ZN(n478) );
  NAND2_X1 U619 ( .A1(n720), .A2(G217), .ZN(n480) );
  XNOR2_X1 U620 ( .A(n481), .B(n745), .ZN(n747) );
  XNOR2_X1 U621 ( .A(n482), .B(G131), .ZN(G33) );
  XNOR2_X2 U622 ( .A(n623), .B(KEYINPUT40), .ZN(n482) );
  XNOR2_X2 U623 ( .A(n484), .B(n610), .ZN(n483) );
  XNOR2_X1 U624 ( .A(n491), .B(n490), .ZN(G60) );
  XNOR2_X2 U625 ( .A(G469), .B(n535), .ZN(n606) );
  XNOR2_X1 U626 ( .A(KEYINPUT121), .B(KEYINPUT59), .ZN(n494) );
  XNOR2_X1 U627 ( .A(n496), .B(n495), .ZN(n497) );
  INV_X1 U628 ( .A(KEYINPUT9), .ZN(n549) );
  XNOR2_X1 U629 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U630 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n504) );
  XOR2_X1 U631 ( .A(KEYINPUT73), .B(KEYINPUT17), .Z(n496) );
  NAND2_X1 U632 ( .A1(G224), .A2(n746), .ZN(n498) );
  XNOR2_X1 U633 ( .A(n501), .B(G119), .ZN(n730) );
  XNOR2_X1 U634 ( .A(n536), .B(n502), .ZN(n505) );
  XNOR2_X1 U635 ( .A(n505), .B(KEYINPUT78), .ZN(n503) );
  NAND2_X1 U636 ( .A1(G214), .A2(n507), .ZN(n675) );
  XNOR2_X1 U637 ( .A(n509), .B(n508), .ZN(n511) );
  NAND2_X1 U638 ( .A1(G952), .A2(n511), .ZN(n510) );
  XNOR2_X1 U639 ( .A(n510), .B(KEYINPUT84), .ZN(n706) );
  OR2_X1 U640 ( .A1(G953), .A2(n706), .ZN(n593) );
  NAND2_X1 U641 ( .A1(G902), .A2(n511), .ZN(n591) );
  INV_X1 U642 ( .A(n591), .ZN(n512) );
  NOR2_X1 U643 ( .A1(G898), .A2(n746), .ZN(n734) );
  NAND2_X1 U644 ( .A1(n512), .A2(n734), .ZN(n513) );
  NAND2_X1 U645 ( .A1(n593), .A2(n513), .ZN(n514) );
  XOR2_X1 U646 ( .A(KEYINPUT87), .B(KEYINPUT25), .Z(n518) );
  INV_X1 U647 ( .A(n515), .ZN(n645) );
  NAND2_X1 U648 ( .A1(G234), .A2(n645), .ZN(n516) );
  XNOR2_X1 U649 ( .A(KEYINPUT20), .B(n516), .ZN(n527) );
  NAND2_X1 U650 ( .A1(n527), .A2(G217), .ZN(n517) );
  XNOR2_X1 U651 ( .A(n518), .B(n517), .ZN(n526) );
  XNOR2_X1 U652 ( .A(G128), .B(G119), .ZN(n519) );
  NAND2_X1 U653 ( .A1(G221), .A2(n546), .ZN(n521) );
  XNOR2_X1 U654 ( .A(n522), .B(n521), .ZN(n525) );
  XNOR2_X1 U655 ( .A(n558), .B(n531), .ZN(n739) );
  XNOR2_X1 U656 ( .A(n525), .B(n739), .ZN(n722) );
  NAND2_X1 U657 ( .A1(n527), .A2(G221), .ZN(n528) );
  XNOR2_X1 U658 ( .A(n528), .B(KEYINPUT21), .ZN(n529) );
  XNOR2_X1 U659 ( .A(KEYINPUT88), .B(n529), .ZN(n596) );
  INV_X1 U660 ( .A(n596), .ZN(n688) );
  NAND2_X1 U661 ( .A1(G227), .A2(n746), .ZN(n532) );
  XNOR2_X1 U662 ( .A(n534), .B(n533), .ZN(n717) );
  NOR2_X1 U663 ( .A1(G902), .A2(n717), .ZN(n535) );
  XOR2_X1 U664 ( .A(KEYINPUT5), .B(KEYINPUT89), .Z(n538) );
  XNOR2_X1 U665 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U666 ( .A(KEYINPUT90), .B(G472), .ZN(n541) );
  INV_X1 U667 ( .A(n580), .ZN(n692) );
  NAND2_X1 U668 ( .A1(n586), .A2(n692), .ZN(n695) );
  NOR2_X1 U669 ( .A1(n588), .A2(n695), .ZN(n542) );
  INV_X1 U670 ( .A(n612), .ZN(n543) );
  NOR2_X1 U671 ( .A1(n588), .A2(n543), .ZN(n544) );
  NAND2_X1 U672 ( .A1(n580), .A2(n544), .ZN(n657) );
  NAND2_X1 U673 ( .A1(n668), .A2(n657), .ZN(n545) );
  XNOR2_X1 U674 ( .A(KEYINPUT98), .B(KEYINPUT7), .ZN(n553) );
  XNOR2_X1 U675 ( .A(n548), .B(G134), .ZN(n550) );
  XNOR2_X1 U676 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U677 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U678 ( .A(n564), .B(n563), .ZN(n565) );
  NAND2_X1 U679 ( .A1(n569), .A2(n585), .ZN(n570) );
  INV_X1 U680 ( .A(n679), .ZN(n571) );
  NOR2_X1 U681 ( .A1(n677), .A2(n596), .ZN(n573) );
  NAND2_X1 U682 ( .A1(n574), .A2(n573), .ZN(n575) );
  INV_X1 U683 ( .A(n686), .ZN(n630) );
  NAND2_X1 U684 ( .A1(n599), .A2(n350), .ZN(n576) );
  NOR2_X1 U685 ( .A1(n576), .A2(n598), .ZN(n577) );
  XNOR2_X1 U686 ( .A(n577), .B(KEYINPUT101), .ZN(n753) );
  AND2_X1 U687 ( .A1(n578), .A2(n753), .ZN(n590) );
  INV_X1 U688 ( .A(KEYINPUT102), .ZN(n579) );
  NAND2_X1 U689 ( .A1(n598), .A2(n599), .ZN(n581) );
  NOR2_X1 U690 ( .A1(n686), .A2(n581), .ZN(n582) );
  XNOR2_X1 U691 ( .A(n583), .B(KEYINPUT83), .ZN(n589) );
  XNOR2_X1 U692 ( .A(KEYINPUT33), .B(n587), .ZN(n707) );
  NOR2_X1 U693 ( .A1(G900), .A2(n591), .ZN(n592) );
  NAND2_X1 U694 ( .A1(G953), .A2(n592), .ZN(n594) );
  NAND2_X1 U695 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U696 ( .A(KEYINPUT75), .B(n595), .ZN(n611) );
  NOR2_X1 U697 ( .A1(n596), .A2(n611), .ZN(n597) );
  XNOR2_X1 U698 ( .A(n601), .B(KEYINPUT111), .ZN(n750) );
  NOR2_X1 U699 ( .A1(KEYINPUT47), .A2(n679), .ZN(n602) );
  XNOR2_X1 U700 ( .A(KEYINPUT68), .B(n602), .ZN(n608) );
  INV_X1 U701 ( .A(n609), .ZN(n603) );
  NOR2_X1 U702 ( .A1(n606), .A2(n605), .ZN(n620) );
  NAND2_X1 U703 ( .A1(n620), .A2(n607), .ZN(n614) );
  INV_X1 U704 ( .A(n614), .ZN(n664) );
  NOR2_X1 U705 ( .A1(n750), .A2(n351), .ZN(n626) );
  INV_X1 U706 ( .A(KEYINPUT30), .ZN(n610) );
  XNOR2_X1 U707 ( .A(n613), .B(KEYINPUT77), .ZN(n616) );
  NAND2_X1 U708 ( .A1(KEYINPUT47), .A2(n614), .ZN(n615) );
  NAND2_X1 U709 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U710 ( .A(n617), .B(KEYINPUT80), .ZN(n625) );
  XOR2_X1 U711 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n621) );
  NAND2_X1 U712 ( .A1(n627), .A2(n675), .ZN(n628) );
  XNOR2_X1 U713 ( .A(KEYINPUT106), .B(n628), .ZN(n629) );
  NOR2_X1 U714 ( .A1(n630), .A2(n629), .ZN(n632) );
  XNOR2_X1 U715 ( .A(KEYINPUT43), .B(KEYINPUT107), .ZN(n631) );
  XNOR2_X1 U716 ( .A(n632), .B(n631), .ZN(n634) );
  NAND2_X1 U717 ( .A1(n634), .A2(n633), .ZN(n674) );
  NAND2_X1 U718 ( .A1(n635), .A2(n674), .ZN(n636) );
  XNOR2_X2 U719 ( .A(n636), .B(KEYINPUT82), .ZN(n640) );
  NAND2_X1 U720 ( .A1(n637), .A2(n660), .ZN(n673) );
  INV_X1 U721 ( .A(n673), .ZN(n638) );
  INV_X1 U722 ( .A(KEYINPUT2), .ZN(n639) );
  BUF_X1 U723 ( .A(n640), .Z(n643) );
  NAND2_X1 U724 ( .A1(KEYINPUT2), .A2(n673), .ZN(n641) );
  XNOR2_X1 U725 ( .A(KEYINPUT76), .B(n641), .ZN(n642) );
  NAND2_X1 U726 ( .A1(n720), .A2(G210), .ZN(n648) );
  BUF_X1 U727 ( .A(n649), .Z(n650) );
  XNOR2_X1 U728 ( .A(n653), .B(KEYINPUT63), .ZN(G57) );
  INV_X1 U729 ( .A(n663), .ZN(n666) );
  NOR2_X1 U730 ( .A1(n666), .A2(n657), .ZN(n654) );
  XOR2_X1 U731 ( .A(G104), .B(n654), .Z(G6) );
  XOR2_X1 U732 ( .A(KEYINPUT112), .B(KEYINPUT26), .Z(n656) );
  XNOR2_X1 U733 ( .A(G107), .B(KEYINPUT27), .ZN(n655) );
  XNOR2_X1 U734 ( .A(n656), .B(n655), .ZN(n659) );
  INV_X1 U735 ( .A(n660), .ZN(n669) );
  NOR2_X1 U736 ( .A1(n669), .A2(n657), .ZN(n658) );
  XOR2_X1 U737 ( .A(n659), .B(n658), .Z(G9) );
  XOR2_X1 U738 ( .A(G128), .B(KEYINPUT29), .Z(n662) );
  NAND2_X1 U739 ( .A1(n660), .A2(n664), .ZN(n661) );
  XNOR2_X1 U740 ( .A(n662), .B(n661), .ZN(G30) );
  NAND2_X1 U741 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U742 ( .A(n665), .B(G146), .ZN(G48) );
  NOR2_X1 U743 ( .A1(n666), .A2(n668), .ZN(n667) );
  XOR2_X1 U744 ( .A(G113), .B(n667), .Z(G15) );
  NOR2_X1 U745 ( .A1(n669), .A2(n668), .ZN(n671) );
  XNOR2_X1 U746 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n670) );
  XNOR2_X1 U747 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U748 ( .A(G116), .B(n672), .ZN(G18) );
  XNOR2_X1 U749 ( .A(G134), .B(n673), .ZN(G36) );
  XNOR2_X1 U750 ( .A(G140), .B(n674), .ZN(G42) );
  NOR2_X1 U751 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U752 ( .A(n678), .B(KEYINPUT116), .ZN(n682) );
  NOR2_X1 U753 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U754 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U755 ( .A1(n683), .A2(n707), .ZN(n684) );
  XNOR2_X1 U756 ( .A(KEYINPUT117), .B(n684), .ZN(n701) );
  NAND2_X1 U757 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U758 ( .A(n687), .B(KEYINPUT50), .ZN(n694) );
  NOR2_X1 U759 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U760 ( .A(KEYINPUT49), .B(n690), .Z(n691) );
  NOR2_X1 U761 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U762 ( .A1(n694), .A2(n693), .ZN(n696) );
  NAND2_X1 U763 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U764 ( .A(n697), .B(KEYINPUT115), .ZN(n698) );
  XNOR2_X1 U765 ( .A(n698), .B(KEYINPUT51), .ZN(n699) );
  NAND2_X1 U766 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U767 ( .A(n702), .B(KEYINPUT119), .ZN(n704) );
  XNOR2_X1 U768 ( .A(KEYINPUT52), .B(KEYINPUT118), .ZN(n703) );
  XNOR2_X1 U769 ( .A(n704), .B(n703), .ZN(n705) );
  NOR2_X1 U770 ( .A1(n706), .A2(n705), .ZN(n713) );
  INV_X1 U771 ( .A(n707), .ZN(n708) );
  XNOR2_X1 U772 ( .A(KEYINPUT79), .B(KEYINPUT2), .ZN(n709) );
  NAND2_X1 U773 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U774 ( .A(n714), .B(KEYINPUT120), .ZN(n715) );
  XOR2_X1 U775 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n716) );
  XOR2_X1 U776 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n721) );
  NAND2_X1 U777 ( .A1(n746), .A2(n724), .ZN(n728) );
  NAND2_X1 U778 ( .A1(G953), .A2(G224), .ZN(n725) );
  XNOR2_X1 U779 ( .A(KEYINPUT61), .B(n725), .ZN(n726) );
  NAND2_X1 U780 ( .A1(n726), .A2(G898), .ZN(n727) );
  NAND2_X1 U781 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U782 ( .A(n729), .B(KEYINPUT125), .ZN(n736) );
  XNOR2_X1 U783 ( .A(G101), .B(n730), .ZN(n732) );
  XNOR2_X1 U784 ( .A(n732), .B(n731), .ZN(n733) );
  NOR2_X1 U785 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U786 ( .A(n736), .B(n735), .Z(G69) );
  XOR2_X1 U787 ( .A(KEYINPUT126), .B(n737), .Z(n738) );
  XNOR2_X1 U788 ( .A(n739), .B(n738), .ZN(n740) );
  XOR2_X1 U789 ( .A(n741), .B(n740), .Z(n745) );
  XOR2_X1 U790 ( .A(G227), .B(n745), .Z(n742) );
  NAND2_X1 U791 ( .A1(n742), .A2(G900), .ZN(n743) );
  NAND2_X1 U792 ( .A1(n743), .A2(G953), .ZN(n744) );
  XOR2_X1 U793 ( .A(KEYINPUT127), .B(n744), .Z(n749) );
  NAND2_X1 U794 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U795 ( .A1(n749), .A2(n748), .ZN(G72) );
  XNOR2_X1 U796 ( .A(n750), .B(G125), .ZN(n751) );
  XNOR2_X1 U797 ( .A(n751), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U798 ( .A(G122), .B(n752), .Z(G24) );
  XNOR2_X1 U799 ( .A(G101), .B(n753), .ZN(G3) );
  XOR2_X1 U800 ( .A(n754), .B(G110), .Z(G12) );
  XOR2_X1 U801 ( .A(G119), .B(n755), .Z(G21) );
  XNOR2_X1 U802 ( .A(G143), .B(n756), .ZN(G45) );
  XNOR2_X1 U803 ( .A(n757), .B(G137), .ZN(G39) );
endmodule

