//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 1 1 1 1 1 1 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n820, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924;
  OR3_X1    g000(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n202));
  OAI21_X1  g001(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n203));
  AOI22_X1  g002(.A1(new_n202), .A2(new_n203), .B1(G29gat), .B2(G36gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(G43gat), .B(G50gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n204), .B1(KEYINPUT15), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(KEYINPUT15), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n208), .A2(KEYINPUT17), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(KEYINPUT17), .ZN(new_n210));
  NAND2_X1  g009(.A1(G85gat), .A2(G92gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n211), .B(KEYINPUT7), .ZN(new_n212));
  INV_X1    g011(.A(G99gat), .ZN(new_n213));
  INV_X1    g012(.A(G106gat), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT8), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n212), .B(new_n215), .C1(G85gat), .C2(G92gat), .ZN(new_n216));
  XOR2_X1   g015(.A(G99gat), .B(G106gat), .Z(new_n217));
  XOR2_X1   g016(.A(new_n216), .B(new_n217), .Z(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n209), .A2(new_n210), .A3(new_n219), .ZN(new_n220));
  AND2_X1   g019(.A1(G232gat), .A2(G233gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT41), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n220), .B(new_n222), .C1(new_n208), .C2(new_n219), .ZN(new_n223));
  XOR2_X1   g022(.A(G190gat), .B(G218gat), .Z(new_n224));
  XNOR2_X1  g023(.A(new_n223), .B(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(G134gat), .B(G162gat), .Z(new_n226));
  NOR2_X1   g025(.A1(new_n221), .A2(KEYINPUT41), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g027(.A(new_n225), .B(new_n228), .Z(new_n229));
  XNOR2_X1  g028(.A(G57gat), .B(G64gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT96), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT9), .ZN(new_n232));
  INV_X1    g031(.A(G71gat), .ZN(new_n233));
  INV_X1    g032(.A(G78gat), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n230), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G71gat), .B(G78gat), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n236), .B(new_n237), .C1(new_n231), .C2(new_n235), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(KEYINPUT97), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n237), .B(KEYINPUT95), .ZN(new_n240));
  INV_X1    g039(.A(new_n235), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n240), .B1(new_n241), .B2(new_n230), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  XOR2_X1   g042(.A(KEYINPUT98), .B(KEYINPUT21), .Z(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G127gat), .B(G155gat), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n245), .B(new_n246), .Z(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G15gat), .B(G22gat), .ZN(new_n249));
  INV_X1    g048(.A(G1gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(KEYINPUT16), .A3(new_n250), .ZN(new_n251));
  OAI221_X1 g050(.A(new_n251), .B1(KEYINPUT92), .B2(G8gat), .C1(new_n250), .C2(new_n249), .ZN(new_n252));
  NAND2_X1  g051(.A1(KEYINPUT92), .A2(G8gat), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n252), .B(new_n253), .Z(new_n254));
  INV_X1    g053(.A(KEYINPUT21), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n254), .B1(new_n243), .B2(new_n255), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n256), .B(KEYINPUT99), .Z(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n258));
  OR2_X1    g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n258), .ZN(new_n260));
  XNOR2_X1  g059(.A(G183gat), .B(G211gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(G231gat), .A2(G233gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n259), .A2(new_n260), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n264), .B1(new_n259), .B2(new_n260), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n248), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n259), .A2(new_n260), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(new_n263), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n259), .A2(new_n260), .A3(new_n264), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(new_n247), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n229), .B1(new_n267), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT102), .ZN(new_n273));
  NAND2_X1  g072(.A1(G230gat), .A2(G233gat), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n243), .B(new_n218), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT10), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n239), .A2(new_n218), .A3(KEYINPUT10), .A4(new_n242), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n275), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OR2_X1    g079(.A1(new_n276), .A2(new_n274), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n280), .B1(KEYINPUT100), .B2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G120gat), .B(G148gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT101), .ZN(new_n285));
  XNOR2_X1  g084(.A(G176gat), .B(G204gat), .ZN(new_n286));
  XOR2_X1   g085(.A(new_n285), .B(new_n286), .Z(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n283), .B(new_n288), .C1(KEYINPUT100), .C2(new_n282), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n287), .B1(new_n282), .B2(new_n280), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n272), .A2(new_n273), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n273), .B1(new_n272), .B2(new_n292), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n296));
  NOR2_X1   g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT26), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(KEYINPUT70), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G169gat), .A2(G176gat), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n301), .B1(new_n297), .B2(new_n298), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT70), .B1(new_n297), .B2(new_n298), .ZN(new_n303));
  NOR3_X1   g102(.A1(new_n300), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G183gat), .A2(G190gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n296), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n303), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(new_n299), .ZN(new_n309));
  OAI211_X1 g108(.A(KEYINPUT71), .B(new_n305), .C1(new_n309), .C2(new_n302), .ZN(new_n310));
  XOR2_X1   g109(.A(KEYINPUT67), .B(G190gat), .Z(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT27), .B(G183gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(KEYINPUT69), .A2(KEYINPUT28), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n313), .B1(new_n311), .B2(new_n312), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n307), .A2(new_n310), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n297), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT23), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n297), .A2(KEYINPUT23), .ZN(new_n321));
  INV_X1    g120(.A(new_n301), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n322), .A2(KEYINPUT66), .ZN(new_n323));
  AND3_X1   g122(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n320), .B(new_n321), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT67), .B(G190gat), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT68), .B1(new_n327), .B2(G183gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n305), .B(KEYINPUT24), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT68), .ZN(new_n330));
  INV_X1    g129(.A(G183gat), .ZN(new_n331));
  INV_X1    g130(.A(G190gat), .ZN(new_n332));
  AND2_X1   g131(.A1(new_n332), .A2(KEYINPUT67), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(KEYINPUT67), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n330), .B(new_n331), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n328), .A2(new_n329), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n326), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT25), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT65), .ZN(new_n339));
  INV_X1    g138(.A(G176gat), .ZN(new_n340));
  INV_X1    g139(.A(G169gat), .ZN(new_n341));
  AND2_X1   g140(.A1(new_n341), .A2(KEYINPUT64), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(KEYINPUT64), .ZN(new_n343));
  OAI211_X1 g142(.A(KEYINPUT23), .B(new_n340), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n322), .B1(new_n318), .B2(new_n319), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n339), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT25), .B1(new_n329), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n344), .A2(new_n339), .A3(new_n345), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n347), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G127gat), .B(G134gat), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT1), .ZN(new_n353));
  INV_X1    g152(.A(G113gat), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(KEYINPUT72), .A3(G120gat), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G113gat), .B(G120gat), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT72), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  XOR2_X1   g158(.A(G113gat), .B(G120gat), .Z(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n353), .ZN(new_n361));
  INV_X1    g160(.A(new_n352), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n356), .A2(new_n359), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n317), .A2(new_n338), .A3(new_n351), .A4(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT73), .ZN(new_n365));
  AND3_X1   g164(.A1(new_n344), .A2(new_n339), .A3(new_n345), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n366), .A2(new_n346), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n367), .A2(new_n349), .B1(new_n337), .B2(KEYINPUT25), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT73), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n368), .A2(new_n369), .A3(new_n363), .A4(new_n317), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n317), .A2(new_n338), .A3(new_n351), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n361), .A2(new_n362), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n359), .A2(new_n353), .A3(new_n352), .A4(new_n355), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(G227gat), .A2(G233gat), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n365), .A2(new_n370), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  AND2_X1   g176(.A1(KEYINPUT75), .A2(KEYINPUT34), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT75), .B(KEYINPUT34), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n379), .B1(new_n377), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT32), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n365), .A2(new_n370), .A3(new_n375), .ZN(new_n383));
  INV_X1    g182(.A(new_n376), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT33), .B1(new_n383), .B2(new_n384), .ZN(new_n386));
  XNOR2_X1  g185(.A(G15gat), .B(G43gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(KEYINPUT74), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n388), .B(G71gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n389), .B(new_n213), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NOR3_X1   g190(.A1(new_n385), .A2(new_n386), .A3(new_n391), .ZN(new_n392));
  AOI221_X4 g191(.A(new_n382), .B1(KEYINPUT33), .B2(new_n390), .C1(new_n383), .C2(new_n384), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n381), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n383), .A2(new_n384), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT33), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n391), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n385), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n393), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n377), .A2(new_n380), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n401), .B1(new_n377), .B2(new_n378), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n399), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n394), .A2(new_n403), .ZN(new_n404));
  AND2_X1   g203(.A1(KEYINPUT76), .A2(KEYINPUT36), .ZN(new_n405));
  NOR2_X1   g204(.A1(KEYINPUT76), .A2(KEYINPUT36), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n394), .A2(new_n403), .A3(new_n405), .ZN(new_n409));
  XOR2_X1   g208(.A(KEYINPUT80), .B(KEYINPUT81), .Z(new_n410));
  XNOR2_X1  g209(.A(G8gat), .B(G36gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G64gat), .B(G92gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT79), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT29), .B1(new_n368), .B2(new_n317), .ZN(new_n416));
  NAND2_X1  g215(.A1(G226gat), .A2(G233gat), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n415), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT29), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n371), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n421), .A2(KEYINPUT79), .A3(new_n417), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n371), .A2(new_n418), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT78), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT77), .B(G218gat), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT22), .B1(new_n425), .B2(G211gat), .ZN(new_n426));
  XOR2_X1   g225(.A(G197gat), .B(G204gat), .Z(new_n427));
  OAI21_X1  g226(.A(new_n424), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(G218gat), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT77), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT77), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(G218gat), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n430), .A2(new_n432), .A3(G211gat), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT22), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n427), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n436), .A3(KEYINPUT78), .ZN(new_n437));
  XNOR2_X1  g236(.A(G211gat), .B(G218gat), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n428), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n438), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n435), .A2(new_n436), .A3(KEYINPUT78), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n419), .A2(new_n422), .A3(new_n423), .A4(new_n443), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n416), .A2(new_n418), .ZN(new_n445));
  INV_X1    g244(.A(new_n423), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n442), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n414), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n444), .A2(new_n447), .A3(new_n414), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(KEYINPUT30), .A3(new_n450), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n444), .A2(new_n447), .A3(new_n414), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT30), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n452), .B1(new_n448), .B2(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(G1gat), .B(G29gat), .ZN(new_n455));
  INV_X1    g254(.A(G85gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n455), .B(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(KEYINPUT0), .B(G57gat), .ZN(new_n458));
  XOR2_X1   g257(.A(new_n457), .B(new_n458), .Z(new_n459));
  INV_X1    g258(.A(G141gat), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n460), .A2(G148gat), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  AND2_X1   g261(.A1(KEYINPUT83), .A2(G148gat), .ZN(new_n463));
  NOR2_X1   g262(.A1(KEYINPUT83), .A2(G148gat), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n462), .B1(new_n465), .B2(new_n460), .ZN(new_n466));
  INV_X1    g265(.A(G155gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT84), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT84), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(G155gat), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n470), .A3(G162gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT2), .ZN(new_n472));
  XNOR2_X1  g271(.A(G155gat), .B(G162gat), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n466), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT82), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT2), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n460), .A2(G148gat), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n476), .B1(new_n461), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(G155gat), .A2(G162gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n479), .B(new_n475), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n478), .B(new_n480), .C1(G155gat), .C2(G162gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n474), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n374), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n363), .A2(new_n474), .A3(new_n481), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT86), .ZN(new_n485));
  NAND2_X1  g284(.A1(G225gat), .A2(G233gat), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT86), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n482), .A2(new_n488), .A3(new_n374), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT5), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n482), .A2(KEYINPUT3), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT3), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n474), .A2(new_n481), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n492), .A2(new_n374), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT85), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n492), .A2(KEYINPUT85), .A3(new_n374), .A4(new_n494), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n482), .A2(new_n374), .A3(KEYINPUT4), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n484), .A2(KEYINPUT4), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n487), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n491), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT87), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n502), .B1(new_n500), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n484), .A2(KEYINPUT87), .A3(KEYINPUT4), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n487), .A2(KEYINPUT5), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n508), .A2(new_n499), .A3(new_n509), .ZN(new_n510));
  OAI211_X1 g309(.A(KEYINPUT6), .B(new_n459), .C1(new_n504), .C2(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n459), .B1(new_n504), .B2(new_n510), .ZN(new_n512));
  INV_X1    g311(.A(new_n459), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n508), .A2(new_n499), .A3(new_n509), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n499), .A2(new_n503), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n513), .B(new_n514), .C1(new_n515), .C2(new_n491), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT6), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n512), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AOI22_X1  g317(.A1(new_n451), .A2(new_n454), .B1(new_n511), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(G22gat), .ZN(new_n520));
  INV_X1    g319(.A(new_n482), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n439), .A2(new_n420), .A3(new_n441), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n521), .B1(new_n522), .B2(new_n493), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n494), .A2(new_n420), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT89), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n494), .A2(KEYINPUT89), .A3(new_n420), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(new_n442), .A3(new_n528), .ZN(new_n529));
  AND2_X1   g328(.A1(G228gat), .A2(G233gat), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n524), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT88), .ZN(new_n532));
  AND3_X1   g331(.A1(new_n442), .A2(new_n525), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n532), .B1(new_n442), .B2(new_n525), .ZN(new_n534));
  NOR3_X1   g333(.A1(new_n533), .A2(new_n523), .A3(new_n534), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n520), .B(new_n531), .C1(new_n535), .C2(new_n530), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT90), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G78gat), .B(G106gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT31), .B(G50gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n531), .B1(new_n535), .B2(new_n530), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(G22gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(new_n536), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n544), .A2(KEYINPUT90), .A3(new_n536), .A4(new_n541), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n408), .B(new_n409), .C1(new_n519), .C2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(KEYINPUT91), .B(KEYINPUT38), .Z(new_n551));
  INV_X1    g350(.A(new_n414), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n552), .A2(KEYINPUT37), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n448), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n444), .A2(new_n447), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n555), .A2(KEYINPUT37), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n551), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n518), .A2(new_n511), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n419), .A2(new_n422), .A3(new_n423), .A4(new_n442), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n443), .B1(new_n445), .B2(new_n446), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n559), .A2(KEYINPUT37), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n551), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n561), .B(new_n562), .C1(new_n448), .C2(new_n553), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n557), .A2(new_n558), .A3(new_n450), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n508), .A2(new_n499), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(new_n487), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n485), .A2(new_n489), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(new_n486), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(KEYINPUT39), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT39), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n565), .A2(new_n570), .A3(new_n487), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n569), .A2(new_n513), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT40), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n512), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n575), .B1(new_n572), .B2(new_n573), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n574), .A2(new_n576), .A3(new_n454), .A4(new_n451), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n564), .A2(new_n548), .A3(new_n577), .ZN(new_n578));
  NOR3_X1   g377(.A1(new_n392), .A2(new_n381), .A3(new_n393), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n402), .B1(new_n399), .B2(new_n400), .ZN(new_n580));
  INV_X1    g379(.A(new_n547), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n538), .A2(new_n541), .B1(new_n544), .B2(new_n536), .ZN(new_n582));
  OAI22_X1  g381(.A1(new_n579), .A2(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n518), .A2(new_n511), .ZN(new_n584));
  NOR3_X1   g383(.A1(new_n452), .A2(new_n448), .A3(new_n453), .ZN(new_n585));
  NOR3_X1   g384(.A1(new_n555), .A2(KEYINPUT30), .A3(new_n552), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT35), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n403), .A2(new_n394), .B1(new_n546), .B2(new_n547), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT35), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n589), .A2(new_n590), .A3(new_n519), .ZN(new_n591));
  AOI22_X1  g390(.A1(new_n550), .A2(new_n578), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n295), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n209), .A2(new_n254), .A3(new_n210), .ZN(new_n594));
  OR2_X1    g393(.A1(new_n254), .A2(new_n208), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G229gat), .A2(G233gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT93), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT18), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n254), .A2(new_n208), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n595), .A2(KEYINPUT94), .A3(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n597), .B(KEYINPUT13), .Z(new_n603));
  INV_X1    g402(.A(KEYINPUT94), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n254), .A2(new_n604), .A3(new_n208), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n602), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT18), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n598), .A2(KEYINPUT93), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n600), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G113gat), .B(G141gat), .ZN(new_n610));
  INV_X1    g409(.A(G197gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(KEYINPUT11), .B(G169gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n614), .B(KEYINPUT12), .Z(new_n615));
  NAND2_X1  g414(.A1(new_n609), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n615), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n600), .A2(new_n606), .A3(new_n608), .A4(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n593), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n620), .A2(new_n584), .ZN(new_n621));
  XOR2_X1   g420(.A(KEYINPUT103), .B(G1gat), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(G1324gat));
  INV_X1    g422(.A(new_n620), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n585), .A2(new_n586), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT42), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT16), .B(G8gat), .ZN(new_n628));
  OR3_X1    g427(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(G8gat), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n627), .B1(new_n626), .B2(new_n628), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(G1325gat));
  AOI21_X1  g431(.A(G15gat), .B1(new_n624), .B2(new_n404), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n408), .A2(new_n409), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n634), .A2(KEYINPUT104), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(KEYINPUT104), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n620), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n633), .B1(G15gat), .B2(new_n639), .ZN(G1326gat));
  INV_X1    g439(.A(new_n548), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n624), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT105), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT43), .B(G22gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(G1327gat));
  AND3_X1   g444(.A1(new_n564), .A2(new_n548), .A3(new_n577), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n590), .B1(new_n589), .B2(new_n519), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n583), .A2(new_n587), .A3(KEYINPUT35), .ZN(new_n648));
  OAI22_X1  g447(.A1(new_n646), .A2(new_n549), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n267), .A2(new_n271), .ZN(new_n650));
  INV_X1    g449(.A(new_n619), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n650), .A2(new_n651), .A3(new_n291), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n649), .A2(new_n652), .A3(new_n229), .ZN(new_n653));
  INV_X1    g452(.A(G29gat), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n653), .A2(new_n654), .A3(new_n558), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT45), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n550), .A2(new_n578), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT106), .ZN(new_n658));
  AND3_X1   g457(.A1(new_n588), .A2(new_n658), .A3(new_n591), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n658), .B1(new_n588), .B2(new_n591), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT44), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n661), .A2(new_n662), .A3(new_n229), .ZN(new_n663));
  INV_X1    g462(.A(new_n229), .ZN(new_n664));
  OAI21_X1  g463(.A(KEYINPUT44), .B1(new_n592), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n666), .A2(new_n652), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n667), .A2(new_n558), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n656), .B1(new_n668), .B2(new_n654), .ZN(G1328gat));
  INV_X1    g468(.A(G36gat), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n653), .A2(new_n670), .A3(new_n625), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n671), .B(KEYINPUT46), .Z(new_n672));
  AND2_X1   g471(.A1(new_n667), .A2(new_n625), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n672), .B1(new_n673), .B2(new_n670), .ZN(G1329gat));
  INV_X1    g473(.A(G43gat), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n653), .A2(new_n675), .A3(new_n404), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n667), .A2(KEYINPUT107), .A3(new_n634), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(G43gat), .ZN(new_n678));
  AOI21_X1  g477(.A(KEYINPUT107), .B1(new_n667), .B2(new_n634), .ZN(new_n679));
  OAI211_X1 g478(.A(KEYINPUT47), .B(new_n676), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n676), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n667), .A2(new_n637), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n681), .B1(new_n682), .B2(G43gat), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n680), .B1(KEYINPUT47), .B2(new_n683), .ZN(G1330gat));
  INV_X1    g483(.A(KEYINPUT109), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n667), .A2(new_n641), .ZN(new_n686));
  INV_X1    g485(.A(G50gat), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n641), .A2(KEYINPUT108), .A3(new_n687), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT108), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(new_n548), .B2(G50gat), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n653), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n692), .B1(new_n686), .B2(new_n687), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT48), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n688), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  OAI221_X1 g494(.A(new_n692), .B1(new_n685), .B2(KEYINPUT48), .C1(new_n686), .C2(new_n687), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(G1331gat));
  AND2_X1   g496(.A1(new_n272), .A2(new_n651), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n661), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(new_n291), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n584), .B(KEYINPUT110), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(G57gat), .ZN(G1332gat));
  INV_X1    g504(.A(new_n625), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n700), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n708));
  AND2_X1   g507(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n707), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n710), .B1(new_n707), .B2(new_n708), .ZN(G1333gat));
  AND3_X1   g510(.A1(new_n699), .A2(new_n404), .A3(new_n291), .ZN(new_n712));
  OR2_X1    g511(.A1(new_n712), .A2(KEYINPUT111), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(KEYINPUT111), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n713), .A2(new_n233), .A3(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n701), .A2(G71gat), .A3(new_n637), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1334gat));
  NOR2_X1   g518(.A1(new_n700), .A2(new_n548), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(new_n234), .ZN(G1335gat));
  INV_X1    g520(.A(KEYINPUT114), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n650), .A2(new_n619), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n291), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT113), .B1(new_n666), .B2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT113), .ZN(new_n727));
  AOI211_X1 g526(.A(new_n727), .B(new_n724), .C1(new_n663), .C2(new_n665), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n722), .B1(new_n729), .B2(new_n584), .ZN(new_n730));
  OAI211_X1 g529(.A(KEYINPUT114), .B(new_n558), .C1(new_n726), .C2(new_n728), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n730), .A2(G85gat), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n661), .A2(new_n229), .A3(new_n723), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(KEYINPUT51), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT51), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n661), .A2(new_n735), .A3(new_n229), .A4(new_n723), .ZN(new_n736));
  AND3_X1   g535(.A1(new_n734), .A2(new_n291), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n737), .A2(new_n456), .A3(new_n558), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n732), .A2(new_n738), .ZN(G1336gat));
  AOI21_X1  g538(.A(new_n662), .B1(new_n649), .B2(new_n229), .ZN(new_n740));
  OAI21_X1  g539(.A(KEYINPUT106), .B1(new_n648), .B2(new_n647), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n588), .A2(new_n591), .A3(new_n658), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n664), .B1(new_n743), .B2(new_n657), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n740), .B1(new_n744), .B2(new_n662), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n727), .B1(new_n745), .B2(new_n724), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n666), .A2(KEYINPUT113), .A3(new_n725), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n706), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(G92gat), .ZN(new_n749));
  OAI21_X1  g548(.A(KEYINPUT115), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n737), .A2(new_n749), .A3(new_n625), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n625), .B1(new_n726), .B2(new_n728), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT115), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n752), .A2(new_n753), .A3(G92gat), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n750), .A2(new_n751), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(KEYINPUT52), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n745), .A2(new_n706), .A3(new_n724), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n751), .B(new_n757), .C1(new_n749), .C2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n756), .A2(new_n759), .ZN(G1337gat));
  OAI21_X1  g559(.A(G99gat), .B1(new_n729), .B2(new_n638), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n737), .A2(new_n213), .A3(new_n404), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(G1338gat));
  NAND3_X1  g562(.A1(new_n737), .A2(new_n214), .A3(new_n641), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT53), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n745), .A2(new_n548), .A3(new_n724), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n764), .B(new_n765), .C1(new_n214), .C2(new_n766), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n734), .A2(new_n641), .A3(new_n291), .A4(new_n736), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n768), .A2(G106gat), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n641), .B1(new_n726), .B2(new_n728), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n769), .B1(new_n770), .B2(G106gat), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT116), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n771), .A2(new_n772), .A3(new_n765), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n548), .B1(new_n746), .B2(new_n747), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n764), .B1(new_n774), .B2(new_n214), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT116), .B1(new_n775), .B2(KEYINPUT53), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n767), .B1(new_n773), .B2(new_n776), .ZN(G1339gat));
  INV_X1    g576(.A(new_n650), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n278), .A2(new_n279), .A3(new_n275), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT117), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n280), .B2(new_n780), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n278), .A2(KEYINPUT117), .A3(new_n279), .A4(new_n275), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n781), .A2(KEYINPUT54), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n288), .B1(new_n280), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n783), .A2(KEYINPUT55), .A3(new_n785), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n788), .A2(new_n619), .A3(new_n289), .A4(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n596), .A2(new_n597), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n603), .B1(new_n602), .B2(new_n605), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n614), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OR2_X1    g594(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n291), .A2(new_n618), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n229), .B1(new_n790), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n788), .A2(new_n289), .A3(new_n789), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n796), .A2(new_n618), .A3(new_n795), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n799), .A2(new_n664), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n778), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n698), .A2(new_n292), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR4_X1   g603(.A1(new_n804), .A2(new_n625), .A3(new_n583), .A4(new_n702), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n805), .A2(new_n354), .A3(new_n619), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT119), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n625), .A2(new_n584), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n804), .A2(new_n583), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n619), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n807), .B1(new_n811), .B2(G113gat), .ZN(new_n812));
  AOI211_X1 g611(.A(KEYINPUT119), .B(new_n354), .C1(new_n810), .C2(new_n619), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n806), .B1(new_n812), .B2(new_n813), .ZN(G1340gat));
  INV_X1    g613(.A(new_n810), .ZN(new_n815));
  OAI21_X1  g614(.A(G120gat), .B1(new_n815), .B2(new_n292), .ZN(new_n816));
  INV_X1    g615(.A(G120gat), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n805), .A2(new_n817), .A3(new_n291), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(G1341gat));
  AOI21_X1  g618(.A(G127gat), .B1(new_n805), .B2(new_n650), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n650), .A2(G127gat), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n820), .B1(new_n810), .B2(new_n821), .ZN(G1342gat));
  INV_X1    g621(.A(G134gat), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n805), .A2(new_n823), .A3(new_n229), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n824), .A2(KEYINPUT56), .ZN(new_n825));
  OAI21_X1  g624(.A(G134gat), .B1(new_n815), .B2(new_n664), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(KEYINPUT56), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(G1343gat));
  NOR2_X1   g627(.A1(new_n809), .A2(new_n634), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n802), .A2(new_n803), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT57), .B1(new_n830), .B2(new_n641), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832));
  AOI211_X1 g631(.A(new_n832), .B(new_n548), .C1(new_n802), .C2(new_n803), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n619), .B(new_n829), .C1(new_n831), .C2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(G141gat), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(KEYINPUT58), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n638), .A2(new_n641), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n804), .B1(KEYINPUT120), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n838), .A2(KEYINPUT120), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n840), .A2(new_n625), .A3(new_n702), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n839), .A2(new_n460), .A3(new_n841), .A4(new_n619), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n835), .A2(new_n837), .A3(new_n842), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n836), .A2(KEYINPUT58), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n843), .B(new_n844), .ZN(G1344gat));
  AND2_X1   g644(.A1(new_n839), .A2(new_n841), .ZN(new_n846));
  INV_X1    g645(.A(new_n465), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(new_n847), .A3(new_n291), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n291), .B(new_n829), .C1(new_n831), .C2(new_n833), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n847), .A2(KEYINPUT59), .ZN(new_n850));
  AND3_X1   g649(.A1(new_n849), .A2(KEYINPUT122), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(KEYINPUT122), .B1(new_n849), .B2(new_n850), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n802), .B1(new_n295), .B2(new_n619), .ZN(new_n855));
  AOI21_X1  g654(.A(KEYINPUT57), .B1(new_n855), .B2(new_n641), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n856), .A2(new_n833), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(new_n291), .A3(new_n829), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n854), .B1(new_n858), .B2(G148gat), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n848), .B1(new_n853), .B2(new_n859), .ZN(G1345gat));
  NAND2_X1  g659(.A1(new_n846), .A2(new_n650), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n468), .A2(new_n470), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n831), .A2(new_n833), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n863), .A2(new_n634), .A3(new_n809), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n778), .A2(new_n862), .ZN(new_n865));
  XOR2_X1   g664(.A(new_n865), .B(KEYINPUT123), .Z(new_n866));
  AOI22_X1  g665(.A1(new_n861), .A2(new_n862), .B1(new_n864), .B2(new_n866), .ZN(G1346gat));
  AOI21_X1  g666(.A(G162gat), .B1(new_n846), .B2(new_n229), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n229), .A2(G162gat), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n868), .B1(new_n864), .B2(new_n869), .ZN(G1347gat));
  NOR4_X1   g669(.A1(new_n804), .A2(new_n558), .A3(new_n706), .A4(new_n583), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n871), .B(new_n619), .C1(new_n342), .C2(new_n343), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n804), .A2(new_n583), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n703), .A2(new_n706), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(G169gat), .B1(new_n875), .B2(new_n651), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n872), .A2(new_n876), .ZN(G1348gat));
  NOR3_X1   g676(.A1(new_n875), .A2(new_n340), .A3(new_n292), .ZN(new_n878));
  AOI21_X1  g677(.A(G176gat), .B1(new_n871), .B2(new_n291), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(G1349gat));
  INV_X1    g679(.A(new_n875), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n331), .B1(new_n881), .B2(new_n650), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n873), .A2(new_n584), .A3(new_n625), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n650), .A2(new_n312), .ZN(new_n884));
  OAI21_X1  g683(.A(KEYINPUT124), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OR3_X1    g684(.A1(new_n882), .A2(new_n885), .A3(KEYINPUT60), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT60), .B1(new_n882), .B2(new_n885), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(G1350gat));
  NAND3_X1  g687(.A1(new_n871), .A2(new_n311), .A3(new_n229), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n881), .A2(new_n229), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n890), .B1(new_n891), .B2(G190gat), .ZN(new_n892));
  AOI211_X1 g691(.A(KEYINPUT61), .B(new_n332), .C1(new_n881), .C2(new_n229), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n889), .B1(new_n892), .B2(new_n893), .ZN(G1351gat));
  NAND3_X1  g693(.A1(new_n638), .A2(new_n625), .A3(new_n641), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n830), .B(new_n584), .C1(KEYINPUT125), .C2(new_n895), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n895), .A2(KEYINPUT125), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n611), .A3(new_n619), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n856), .A2(new_n833), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n638), .A2(new_n874), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n619), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n899), .B1(new_n904), .B2(new_n611), .ZN(G1352gat));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n896), .A2(G204gat), .A3(new_n897), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(new_n907), .B2(new_n291), .ZN(new_n908));
  INV_X1    g707(.A(new_n901), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n857), .A2(new_n291), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n908), .B1(G204gat), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n907), .A2(new_n906), .A3(new_n291), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n912), .A2(KEYINPUT126), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(KEYINPUT126), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n911), .A2(new_n913), .A3(new_n914), .ZN(G1353gat));
  INV_X1    g714(.A(G211gat), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n898), .A2(new_n916), .A3(new_n650), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n857), .A2(new_n650), .A3(new_n909), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n918), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n919));
  AOI21_X1  g718(.A(KEYINPUT63), .B1(new_n918), .B2(G211gat), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n917), .B1(new_n919), .B2(new_n920), .ZN(G1354gat));
  AOI21_X1  g720(.A(G218gat), .B1(new_n898), .B2(new_n229), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n229), .A2(new_n425), .ZN(new_n923));
  XOR2_X1   g722(.A(new_n923), .B(KEYINPUT127), .Z(new_n924));
  AOI21_X1  g723(.A(new_n922), .B1(new_n902), .B2(new_n924), .ZN(G1355gat));
endmodule


