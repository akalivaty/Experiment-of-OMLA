//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 1 1 1 1 1 1 0 0 1 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n814, new_n816, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n986, new_n987, new_n988, new_n989, new_n990, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G43gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G71gat), .B(G99gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G169gat), .ZN(new_n206));
  INV_X1    g005(.A(G176gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT23), .ZN(new_n208));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT65), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n211), .A2(G169gat), .A3(G176gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n208), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT66), .ZN(new_n214));
  NOR2_X1   g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215));
  AOI22_X1  g014(.A1(new_n215), .A2(KEYINPUT23), .B1(new_n209), .B2(KEYINPUT65), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(new_n217), .A3(new_n212), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n214), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT24), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n220), .A2(G183gat), .A3(G190gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(G183gat), .B(G190gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n221), .B1(new_n222), .B2(new_n220), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n207), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT25), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n223), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G190gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n229), .A2(G183gat), .ZN(new_n230));
  INV_X1    g029(.A(G183gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n231), .A2(G190gat), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT24), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  AND2_X1   g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n234), .B1(KEYINPUT23), .B2(new_n215), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n233), .A2(new_n221), .A3(new_n235), .A4(new_n226), .ZN(new_n236));
  XOR2_X1   g035(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n237));
  AOI22_X1  g036(.A1(new_n219), .A2(new_n228), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n224), .A2(KEYINPUT26), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT26), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n209), .B1(new_n215), .B2(new_n240), .ZN(new_n241));
  OAI22_X1  g040(.A1(new_n239), .A2(new_n241), .B1(new_n231), .B2(new_n229), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT27), .B(G183gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT28), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n244), .A2(G190gat), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT69), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT27), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT27), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(G183gat), .ZN(new_n249));
  AND4_X1   g048(.A1(KEYINPUT69), .A2(new_n245), .A3(new_n247), .A4(new_n249), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(KEYINPUT68), .B1(new_n231), .B2(KEYINPUT27), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n253), .A2(new_n248), .A3(G183gat), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(new_n231), .A3(KEYINPUT27), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n252), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n248), .A2(G183gat), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n229), .B1(new_n258), .B2(new_n255), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n244), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n242), .B1(new_n251), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT71), .B1(new_n238), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G120gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(G113gat), .ZN(new_n264));
  INV_X1    g063(.A(G113gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G120gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT1), .ZN(new_n268));
  XNOR2_X1  g067(.A(G127gat), .B(G134gat), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT70), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n267), .B(new_n268), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(G134gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(G127gat), .ZN(new_n273));
  INV_X1    g072(.A(G127gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(G134gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n270), .A2(new_n268), .ZN(new_n277));
  XNOR2_X1  g076(.A(G113gat), .B(G120gat), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n276), .B(new_n277), .C1(new_n278), .C2(KEYINPUT1), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n271), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n226), .A2(new_n209), .A3(new_n208), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n237), .B1(new_n223), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n217), .B1(new_n216), .B2(new_n212), .ZN(new_n283));
  AND4_X1   g082(.A1(new_n217), .A2(new_n208), .A3(new_n210), .A4(new_n212), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n233), .A2(KEYINPUT25), .A3(new_n221), .A4(new_n226), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n282), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n288));
  INV_X1    g087(.A(new_n242), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n252), .A2(new_n254), .A3(new_n256), .ZN(new_n290));
  AOI21_X1  g089(.A(G190gat), .B1(new_n247), .B2(KEYINPUT67), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT28), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n245), .A2(new_n247), .A3(new_n249), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT69), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n243), .A2(KEYINPUT69), .A3(new_n245), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n289), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n287), .A2(new_n288), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n262), .A2(new_n280), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G227gat), .A2(G233gat), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n271), .A2(new_n279), .ZN(new_n303));
  OAI211_X1 g102(.A(KEYINPUT71), .B(new_n303), .C1(new_n238), .C2(new_n261), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n300), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n205), .B1(new_n305), .B2(KEYINPUT32), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT33), .ZN(new_n307));
  AND3_X1   g106(.A1(new_n305), .A2(KEYINPUT72), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT72), .B1(new_n305), .B2(new_n307), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n306), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT34), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n311), .B1(new_n301), .B2(KEYINPUT73), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n300), .A2(new_n304), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n313), .B1(new_n314), .B2(new_n301), .ZN(new_n315));
  AOI211_X1 g114(.A(new_n302), .B(new_n312), .C1(new_n300), .C2(new_n304), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n305), .B(KEYINPUT32), .C1(new_n307), .C2(new_n205), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n310), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n317), .B1(new_n310), .B2(new_n318), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n202), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n318), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n305), .A2(new_n307), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT72), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n305), .A2(KEYINPUT72), .A3(new_n307), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n323), .B1(new_n328), .B2(new_n306), .ZN(new_n329));
  INV_X1    g128(.A(new_n315), .ZN(new_n330));
  INV_X1    g129(.A(new_n316), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT74), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT74), .B1(new_n315), .B2(new_n316), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n319), .B(KEYINPUT36), .C1(new_n329), .C2(new_n335), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n322), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT85), .ZN(new_n338));
  XOR2_X1   g137(.A(G155gat), .B(G162gat), .Z(new_n339));
  XNOR2_X1  g138(.A(G141gat), .B(G148gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(KEYINPUT78), .B(KEYINPUT2), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AND2_X1   g141(.A1(G141gat), .A2(G148gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(G141gat), .A2(G148gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G155gat), .B(G162gat), .ZN(new_n346));
  INV_X1    g145(.A(G155gat), .ZN(new_n347));
  INV_X1    g146(.A(G162gat), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT2), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n345), .A2(new_n346), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n342), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT29), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G197gat), .B(G204gat), .ZN(new_n355));
  INV_X1    g154(.A(G211gat), .ZN(new_n356));
  INV_X1    g155(.A(G218gat), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n355), .B1(KEYINPUT22), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G211gat), .B(G218gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n360), .B(new_n355), .C1(KEYINPUT22), .C2(new_n358), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n354), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G228gat), .A2(G233gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT3), .B1(new_n364), .B2(new_n353), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n342), .A2(new_n350), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n366), .B(new_n368), .C1(new_n369), .C2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n364), .B1(new_n353), .B2(new_n352), .ZN(new_n373));
  NOR2_X1   g172(.A1(G211gat), .A2(G218gat), .ZN(new_n374));
  AOI211_X1 g173(.A(new_n374), .B(new_n358), .C1(new_n355), .C2(KEYINPUT22), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT29), .B1(new_n375), .B2(KEYINPUT84), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT84), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n362), .A2(new_n377), .A3(new_n363), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(new_n351), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n345), .A2(new_n346), .A3(new_n349), .ZN(new_n381));
  AND2_X1   g180(.A1(KEYINPUT78), .A2(KEYINPUT2), .ZN(new_n382));
  NOR2_X1   g181(.A1(KEYINPUT78), .A2(KEYINPUT2), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n346), .B1(new_n345), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT79), .B1(new_n381), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT79), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n342), .A2(new_n350), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n373), .B1(new_n380), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n372), .B1(new_n390), .B2(new_n368), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(G22gat), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT3), .B1(new_n376), .B2(new_n378), .ZN(new_n393));
  INV_X1    g192(.A(new_n389), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n366), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OR2_X1    g194(.A1(new_n369), .A2(new_n371), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n373), .A2(new_n367), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n395), .A2(new_n367), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(G22gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(G50gat), .ZN(new_n402));
  XOR2_X1   g201(.A(G78gat), .B(G106gat), .Z(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  AND4_X1   g203(.A1(new_n338), .A2(new_n392), .A3(new_n400), .A4(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT85), .B1(new_n398), .B2(new_n399), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n406), .A2(new_n404), .B1(new_n392), .B2(new_n400), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n353), .B1(new_n238), .B2(new_n261), .ZN(new_n409));
  NAND2_X1  g208(.A1(G226gat), .A2(G233gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n410), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n412), .B1(new_n238), .B2(new_n261), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT75), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT75), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n415), .B1(new_n409), .B2(new_n410), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n364), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT88), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT37), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n410), .B1(new_n287), .B2(new_n298), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n420), .B1(new_n410), .B2(new_n409), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n419), .B1(new_n421), .B2(new_n365), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n417), .A2(new_n418), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n418), .B1(new_n417), .B2(new_n422), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT38), .ZN(new_n426));
  XNOR2_X1  g225(.A(G8gat), .B(G36gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(G64gat), .B(G92gat), .ZN(new_n428));
  XOR2_X1   g227(.A(new_n427), .B(new_n428), .Z(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n365), .B1(new_n414), .B2(new_n416), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT29), .B1(new_n287), .B2(new_n298), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n364), .B(new_n413), .C1(new_n432), .C2(new_n412), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT76), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT76), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n411), .A2(new_n435), .A3(new_n364), .A4(new_n413), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n431), .A2(new_n437), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n426), .B(new_n430), .C1(new_n438), .C2(KEYINPUT37), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n425), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n411), .A2(KEYINPUT75), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n441), .B1(new_n421), .B2(KEYINPUT75), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n442), .A2(new_n365), .B1(new_n434), .B2(new_n436), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n429), .B1(new_n443), .B2(new_n419), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n438), .A2(KEYINPUT37), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n426), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n431), .A2(new_n437), .A3(new_n429), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT77), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT80), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT4), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n386), .A2(new_n303), .A3(new_n450), .A4(new_n388), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT4), .B1(new_n280), .B2(new_n370), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT5), .ZN(new_n454));
  NAND2_X1  g253(.A1(G225gat), .A2(G233gat), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n352), .A2(new_n280), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n351), .B1(new_n342), .B2(new_n350), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n454), .B(new_n455), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n449), .B1(new_n453), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n458), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n451), .A2(new_n452), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(KEYINPUT80), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n456), .ZN(new_n463));
  INV_X1    g262(.A(new_n457), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n386), .A2(new_n303), .A3(KEYINPUT4), .A4(new_n388), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n450), .B1(new_n280), .B2(new_n370), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n465), .A2(new_n466), .A3(new_n455), .A4(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n280), .B(new_n370), .ZN(new_n469));
  INV_X1    g268(.A(new_n455), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n454), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI22_X1  g270(.A1(new_n459), .A2(new_n462), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(G1gat), .B(G29gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(KEYINPUT0), .ZN(new_n474));
  XNOR2_X1  g273(.A(G57gat), .B(G85gat), .ZN(new_n475));
  XOR2_X1   g274(.A(new_n474), .B(new_n475), .Z(new_n476));
  AOI21_X1  g275(.A(KEYINPUT6), .B1(new_n472), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n468), .A2(new_n471), .ZN(new_n478));
  NOR3_X1   g277(.A1(new_n453), .A2(new_n449), .A3(new_n458), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT80), .B1(new_n460), .B2(new_n461), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n476), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n481), .A2(KEYINPUT6), .A3(new_n482), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT77), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n431), .A2(new_n437), .A3(new_n486), .A4(new_n429), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n448), .A2(new_n484), .A3(new_n485), .A4(new_n487), .ZN(new_n488));
  NOR3_X1   g287(.A1(new_n440), .A2(new_n446), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n461), .A2(new_n465), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(new_n470), .ZN(new_n491));
  OR3_X1    g290(.A1(new_n469), .A2(KEYINPUT87), .A3(new_n470), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT87), .B1(new_n469), .B2(new_n470), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT39), .A4(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(KEYINPUT86), .B(KEYINPUT39), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n490), .A2(new_n470), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n494), .A2(new_n476), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT40), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n498), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(new_n483), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT30), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n448), .A2(new_n502), .A3(new_n487), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n429), .B1(new_n431), .B2(new_n437), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n431), .A2(new_n437), .A3(new_n429), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n504), .B1(new_n505), .B2(KEYINPUT30), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n501), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n408), .B1(new_n489), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT81), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n509), .B1(new_n472), .B2(new_n476), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n481), .A2(KEYINPUT81), .A3(new_n482), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n510), .A2(new_n477), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(new_n485), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n513), .A2(new_n503), .A3(new_n506), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT82), .ZN(new_n515));
  INV_X1    g314(.A(new_n408), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT82), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n513), .A2(new_n503), .A3(new_n517), .A4(new_n506), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n515), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n337), .B1(new_n508), .B2(new_n519), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n408), .B(new_n319), .C1(new_n329), .C2(new_n335), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n515), .A2(new_n518), .A3(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n320), .A2(new_n321), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n503), .A2(new_n506), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT35), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n408), .A2(new_n526), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n484), .A2(new_n485), .ZN(new_n528));
  NOR3_X1   g327(.A1(new_n525), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI22_X1  g328(.A1(new_n523), .A2(KEYINPUT35), .B1(new_n524), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n520), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G229gat), .A2(G233gat), .ZN(new_n532));
  XOR2_X1   g331(.A(new_n532), .B(KEYINPUT13), .Z(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(G15gat), .B(G22gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT93), .ZN(new_n536));
  INV_X1    g335(.A(G1gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT16), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n535), .A2(KEYINPUT93), .A3(G1gat), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n538), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(G8gat), .ZN(new_n543));
  OAI21_X1  g342(.A(KEYINPUT94), .B1(new_n535), .B2(G1gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n543), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n546), .A2(new_n538), .A3(new_n540), .A4(new_n541), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(G50gat), .ZN(new_n549));
  AND2_X1   g348(.A1(KEYINPUT90), .A2(G43gat), .ZN(new_n550));
  NOR2_X1   g349(.A1(KEYINPUT90), .A2(G43gat), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT91), .B1(new_n549), .B2(G43gat), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT15), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT91), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n557), .B(new_n549), .C1(new_n550), .C2(new_n551), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n555), .A2(KEYINPUT92), .A3(new_n556), .A4(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G29gat), .A2(G36gat), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT89), .B1(G29gat), .B2(G36gat), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n560), .B1(new_n561), .B2(KEYINPUT14), .ZN(new_n562));
  INV_X1    g361(.A(new_n561), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT14), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OR3_X1    g364(.A1(KEYINPUT89), .A2(G29gat), .A3(G36gat), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n562), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n559), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n549), .A2(G43gat), .ZN(new_n569));
  INV_X1    g368(.A(G43gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(G50gat), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n569), .A2(new_n571), .A3(KEYINPUT15), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT90), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(new_n570), .ZN(new_n575));
  NAND2_X1  g374(.A1(KEYINPUT90), .A2(G43gat), .ZN(new_n576));
  AOI21_X1  g375(.A(G50gat), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT15), .B1(new_n577), .B2(new_n557), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT92), .B1(new_n578), .B2(new_n555), .ZN(new_n579));
  INV_X1    g378(.A(new_n572), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n567), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n548), .A2(new_n573), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n573), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n545), .A2(new_n547), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n534), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n581), .A2(new_n573), .A3(KEYINPUT17), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT17), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n565), .A2(new_n566), .ZN(new_n589));
  INV_X1    g388(.A(new_n562), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT92), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n558), .A2(new_n556), .ZN(new_n593));
  XNOR2_X1  g392(.A(KEYINPUT90), .B(G43gat), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n553), .B1(new_n594), .B2(new_n549), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n592), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n591), .B1(new_n596), .B2(new_n572), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n580), .B1(new_n559), .B2(new_n567), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n588), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n548), .B1(new_n587), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n583), .A2(new_n584), .ZN(new_n601));
  INV_X1    g400(.A(new_n532), .ZN(new_n602));
  NOR3_X1   g401(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n586), .B1(new_n603), .B2(KEYINPUT18), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n599), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n601), .B1(new_n584), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(new_n532), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT18), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G113gat), .B(G141gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(G197gat), .ZN(new_n611));
  XOR2_X1   g410(.A(KEYINPUT11), .B(G169gat), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n604), .B(new_n609), .C1(KEYINPUT95), .C2(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(KEYINPUT17), .B1(new_n581), .B2(new_n573), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n597), .A2(new_n598), .A3(new_n588), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n584), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n618), .A2(KEYINPUT18), .A3(new_n582), .A4(new_n532), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n582), .A2(new_n585), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(new_n533), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n619), .A2(KEYINPUT95), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n614), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n619), .A2(new_n621), .ZN(new_n624));
  AOI21_X1  g423(.A(KEYINPUT18), .B1(new_n606), .B2(new_n532), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n622), .B(new_n623), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n615), .A2(KEYINPUT96), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT96), .B1(new_n615), .B2(new_n626), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n531), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(G85gat), .A2(G92gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(KEYINPUT7), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT7), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n634), .A2(G85gat), .A3(G92gat), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(G99gat), .A2(G106gat), .ZN(new_n637));
  INV_X1    g436(.A(G85gat), .ZN(new_n638));
  INV_X1    g437(.A(G92gat), .ZN(new_n639));
  AOI22_X1  g438(.A1(KEYINPUT8), .A2(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G99gat), .B(G106gat), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n636), .A2(new_n640), .A3(new_n642), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n644), .A2(KEYINPUT101), .A3(new_n645), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT103), .ZN(new_n652));
  XNOR2_X1  g451(.A(G190gat), .B(G218gat), .ZN(new_n653));
  AOI22_X1  g452(.A1(new_n605), .A2(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n650), .A2(new_n573), .A3(new_n581), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT102), .ZN(new_n656));
  NAND2_X1  g455(.A1(G232gat), .A2(G233gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT100), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(KEYINPUT41), .ZN(new_n660));
  AND3_X1   g459(.A1(new_n655), .A2(new_n656), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n656), .B1(new_n655), .B2(new_n660), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n654), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n653), .A2(new_n652), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI221_X1 g464(.A(new_n654), .B1(new_n652), .B2(new_n653), .C1(new_n661), .C2(new_n662), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n659), .A2(KEYINPUT41), .ZN(new_n667));
  XNOR2_X1  g466(.A(G134gat), .B(G162gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n665), .A2(new_n666), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n669), .B1(new_n665), .B2(new_n666), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(G71gat), .A2(G78gat), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(G71gat), .A2(G78gat), .ZN(new_n675));
  AND2_X1   g474(.A1(G57gat), .A2(G64gat), .ZN(new_n676));
  OAI21_X1  g475(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n677));
  OAI211_X1 g476(.A(new_n674), .B(new_n675), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(G64gat), .ZN(new_n679));
  INV_X1    g478(.A(G57gat), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n679), .B1(new_n680), .B2(KEYINPUT98), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT9), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n675), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n675), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n681), .B(new_n683), .C1(new_n684), .C2(new_n673), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT97), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT98), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n686), .A2(new_n687), .A3(G57gat), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n680), .A2(KEYINPUT97), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n679), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n678), .B1(new_n685), .B2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT21), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(G231gat), .A2(G233gat), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XOR2_X1   g494(.A(G127gat), .B(G155gat), .Z(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT20), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n695), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g497(.A(G183gat), .B(G211gat), .Z(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n584), .B1(new_n692), .B2(new_n691), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT99), .B(KEYINPUT19), .Z(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n700), .A2(new_n703), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(G230gat), .A2(G233gat), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT104), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT105), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n710), .B1(new_n636), .B2(new_n640), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n709), .B1(new_n691), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n646), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n646), .B(new_n709), .C1(new_n691), .C2(new_n711), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT10), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n691), .A2(new_n709), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n714), .A2(new_n715), .A3(new_n716), .A4(new_n717), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n691), .A2(new_n716), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n650), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n708), .B1(new_n718), .B2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n714), .A2(new_n715), .A3(new_n717), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n722), .B1(new_n708), .B2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(G120gat), .B(G148gat), .ZN(new_n725));
  XNOR2_X1  g524(.A(G176gat), .B(G204gat), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n725), .B(new_n726), .Z(new_n727));
  OR2_X1    g526(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n724), .A2(new_n727), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n672), .A2(new_n706), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n631), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n733), .A2(new_n513), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(new_n537), .ZN(G1324gat));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n736));
  INV_X1    g535(.A(new_n525), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n733), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n736), .B1(new_n738), .B2(new_n543), .ZN(new_n739));
  OAI211_X1 g538(.A(KEYINPUT106), .B(G8gat), .C1(new_n733), .C2(new_n737), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT42), .ZN(new_n741));
  XOR2_X1   g540(.A(KEYINPUT16), .B(G8gat), .Z(new_n742));
  AND3_X1   g541(.A1(new_n738), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n741), .B1(new_n738), .B2(new_n742), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n739), .B(new_n740), .C1(new_n743), .C2(new_n744), .ZN(G1325gat));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n322), .A2(new_n746), .A3(new_n336), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n746), .B1(new_n322), .B2(new_n336), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(G15gat), .B1(new_n733), .B2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n524), .ZN(new_n751));
  OR2_X1    g550(.A1(new_n751), .A2(G15gat), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n733), .B2(new_n752), .ZN(G1326gat));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n733), .B2(new_n408), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n631), .A2(KEYINPUT108), .A3(new_n516), .A4(new_n732), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(KEYINPUT43), .B(G22gat), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(G1327gat));
  INV_X1    g558(.A(new_n672), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n706), .A2(new_n730), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n629), .B(new_n762), .C1(new_n520), .C2(new_n530), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n763), .A2(G29gat), .A3(new_n513), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n764), .B(KEYINPUT45), .Z(new_n765));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n508), .A2(new_n519), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n523), .A2(KEYINPUT35), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n529), .A2(new_n524), .ZN(new_n769));
  AOI22_X1  g568(.A1(new_n767), .A2(new_n749), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n766), .B1(new_n770), .B2(new_n760), .ZN(new_n771));
  OAI211_X1 g570(.A(KEYINPUT44), .B(new_n672), .C1(new_n520), .C2(new_n530), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n615), .A2(new_n626), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n761), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n771), .A2(new_n772), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(G29gat), .B1(new_n776), .B2(new_n513), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n765), .A2(new_n777), .ZN(G1328gat));
  NOR3_X1   g577(.A1(new_n763), .A2(G36gat), .A3(new_n737), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT46), .ZN(new_n780));
  OAI21_X1  g579(.A(G36gat), .B1(new_n776), .B2(new_n737), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(G1329gat));
  INV_X1    g581(.A(new_n749), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n594), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n763), .A2(new_n751), .ZN(new_n785));
  OAI22_X1  g584(.A1(new_n776), .A2(new_n784), .B1(new_n594), .B2(new_n785), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g586(.A(KEYINPUT109), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n771), .A2(new_n516), .A3(new_n772), .A4(new_n775), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n788), .B1(new_n789), .B2(G50gat), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n763), .A2(G50gat), .A3(new_n408), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n791), .B1(new_n789), .B2(G50gat), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT48), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n790), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  AOI221_X4 g593(.A(new_n791), .B1(new_n788), .B2(KEYINPUT48), .C1(new_n789), .C2(G50gat), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n794), .A2(new_n795), .ZN(G1331gat));
  INV_X1    g595(.A(new_n706), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n760), .A2(new_n797), .A3(new_n774), .A4(new_n731), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n770), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n513), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n686), .A2(G57gat), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n689), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n801), .B(new_n803), .ZN(G1332gat));
  INV_X1    g603(.A(KEYINPUT49), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n525), .B1(new_n805), .B2(new_n679), .ZN(new_n806));
  XOR2_X1   g605(.A(new_n806), .B(KEYINPUT110), .Z(new_n807));
  NAND2_X1  g606(.A1(new_n799), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n805), .A2(new_n679), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n808), .B(new_n809), .ZN(G1333gat));
  NAND2_X1  g609(.A1(new_n799), .A2(new_n783), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n751), .A2(G71gat), .ZN(new_n812));
  AOI22_X1  g611(.A1(new_n811), .A2(G71gat), .B1(new_n799), .B2(new_n812), .ZN(new_n813));
  XNOR2_X1  g612(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n813), .B(new_n814), .ZN(G1334gat));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n516), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g616(.A1(new_n767), .A2(new_n749), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n768), .A2(new_n769), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n760), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n797), .A2(new_n773), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n820), .A2(KEYINPUT51), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT51), .B1(new_n820), .B2(new_n821), .ZN(new_n823));
  OR2_X1    g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n824), .A2(new_n638), .A3(new_n800), .A4(new_n731), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n821), .A2(new_n731), .ZN(new_n826));
  XOR2_X1   g625(.A(new_n826), .B(KEYINPUT112), .Z(new_n827));
  NAND3_X1  g626(.A1(new_n771), .A2(new_n772), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(G85gat), .B1(new_n828), .B2(new_n513), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n825), .A2(new_n829), .ZN(G1336gat));
  OAI21_X1  g629(.A(G92gat), .B1(new_n828), .B2(new_n737), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n737), .A2(G92gat), .A3(new_n730), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n832), .B1(new_n822), .B2(new_n823), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT113), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(new_n836), .A3(KEYINPUT52), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n831), .B(new_n833), .C1(new_n835), .C2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(G1337gat));
  NOR3_X1   g639(.A1(new_n751), .A2(G99gat), .A3(new_n730), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n824), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(G99gat), .B1(new_n828), .B2(new_n749), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(G1338gat));
  OAI21_X1  g643(.A(G106gat), .B1(new_n828), .B2(new_n408), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n408), .A2(new_n730), .A3(G106gat), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n846), .B1(new_n822), .B2(new_n823), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n847), .A3(KEYINPUT114), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT53), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n845), .A2(new_n847), .A3(KEYINPUT114), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n851), .ZN(G1339gat));
  NAND3_X1  g651(.A1(new_n718), .A2(new_n708), .A3(new_n721), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n718), .A2(new_n721), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n707), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n718), .A2(KEYINPUT115), .A3(new_n721), .A4(new_n708), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n855), .A2(new_n857), .A3(KEYINPUT54), .A4(new_n858), .ZN(new_n859));
  XNOR2_X1  g658(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n727), .B1(new_n722), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n859), .A2(KEYINPUT55), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(KEYINPUT117), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n859), .A2(new_n864), .A3(KEYINPUT55), .A4(new_n861), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n863), .A2(new_n729), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(KEYINPUT118), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n863), .A2(new_n868), .A3(new_n729), .A4(new_n865), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n859), .A2(new_n861), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT55), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n867), .A2(new_n773), .A3(new_n869), .A4(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n604), .A2(new_n609), .A3(new_n614), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n606), .A2(new_n532), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n620), .A2(new_n533), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n613), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(new_n730), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n672), .B1(new_n873), .B2(new_n880), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n878), .A2(new_n670), .A3(new_n671), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n882), .A2(new_n867), .A3(new_n869), .A4(new_n872), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n706), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n732), .A2(new_n774), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n525), .A2(new_n513), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n751), .A2(new_n516), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n890), .A2(new_n265), .A3(new_n630), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n887), .A2(new_n800), .A3(new_n522), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n513), .B1(new_n885), .B2(new_n886), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(KEYINPUT119), .A3(new_n522), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n525), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n773), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n891), .B1(new_n898), .B2(new_n265), .ZN(G1340gat));
  NOR3_X1   g698(.A1(new_n890), .A2(new_n263), .A3(new_n730), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n897), .A2(new_n731), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n900), .B1(new_n901), .B2(new_n263), .ZN(G1341gat));
  NAND3_X1  g701(.A1(new_n897), .A2(new_n274), .A3(new_n797), .ZN(new_n903));
  OAI21_X1  g702(.A(G127gat), .B1(new_n890), .B2(new_n706), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(G1342gat));
  NOR3_X1   g704(.A1(new_n760), .A2(new_n525), .A3(G134gat), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n907), .B1(new_n894), .B2(new_n896), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT56), .ZN(new_n909));
  OR3_X1    g708(.A1(new_n908), .A2(KEYINPUT120), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT120), .B1(new_n908), .B2(new_n909), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n908), .A2(new_n909), .ZN(new_n912));
  OAI21_X1  g711(.A(G134gat), .B1(new_n890), .B2(new_n760), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n910), .A2(new_n911), .A3(new_n912), .A4(new_n913), .ZN(G1343gat));
  AND2_X1   g713(.A1(new_n749), .A2(new_n888), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n408), .B1(new_n885), .B2(new_n886), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n916), .A2(KEYINPUT57), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT57), .ZN(new_n918));
  AND4_X1   g717(.A1(new_n729), .A2(new_n863), .A3(new_n865), .A4(new_n872), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT96), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n773), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n615), .A2(new_n626), .A3(KEYINPUT96), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n919), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n672), .B1(new_n923), .B2(new_n880), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n706), .B1(new_n924), .B2(new_n884), .ZN(new_n925));
  AOI211_X1 g724(.A(new_n918), .B(new_n408), .C1(new_n925), .C2(new_n886), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n915), .B1(new_n917), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(G141gat), .B1(new_n927), .B2(new_n630), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n783), .A2(new_n408), .A3(new_n525), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n895), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n630), .A2(G141gat), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT58), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n773), .B(new_n915), .C1(new_n917), .C2(new_n926), .ZN(new_n934));
  AOI22_X1  g733(.A1(new_n934), .A2(G141gat), .B1(new_n930), .B2(new_n931), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT58), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(G1344gat));
  NOR3_X1   g736(.A1(new_n927), .A2(KEYINPUT59), .A3(new_n730), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n930), .A2(new_n731), .ZN(new_n939));
  AOI21_X1  g738(.A(G148gat), .B1(new_n939), .B2(KEYINPUT59), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n630), .A2(new_n732), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n408), .B1(new_n925), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g742(.A(KEYINPUT121), .B1(new_n943), .B2(KEYINPUT57), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT121), .ZN(new_n945));
  INV_X1    g744(.A(new_n942), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n879), .B1(new_n629), .B2(new_n919), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n883), .B1(new_n947), .B2(new_n672), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n948), .B2(new_n706), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n945), .B(new_n918), .C1(new_n949), .C2(new_n408), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n887), .A2(KEYINPUT57), .A3(new_n516), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n944), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n952), .A2(new_n731), .A3(new_n915), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n953), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n941), .A2(new_n954), .ZN(G1345gat));
  OAI21_X1  g754(.A(G155gat), .B1(new_n927), .B2(new_n706), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n930), .A2(new_n347), .A3(new_n797), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(G1346gat));
  OAI21_X1  g757(.A(G162gat), .B1(new_n927), .B2(new_n760), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n930), .A2(new_n348), .A3(new_n672), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(G1347gat));
  NOR2_X1   g760(.A1(new_n737), .A2(new_n800), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n887), .A2(new_n889), .A3(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT122), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND4_X1  g764(.A1(new_n887), .A2(KEYINPUT122), .A3(new_n889), .A4(new_n962), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n630), .A2(new_n206), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(new_n962), .ZN(new_n969));
  AOI211_X1 g768(.A(new_n521), .B(new_n969), .C1(new_n885), .C2(new_n886), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n970), .A2(new_n773), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n968), .B1(new_n971), .B2(G169gat), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT123), .ZN(new_n973));
  XNOR2_X1  g772(.A(new_n972), .B(new_n973), .ZN(G1348gat));
  NAND3_X1  g773(.A1(new_n965), .A2(new_n731), .A3(new_n966), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(G176gat), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n970), .A2(new_n207), .A3(new_n731), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(G1349gat));
  NAND3_X1  g777(.A1(new_n965), .A2(new_n797), .A3(new_n966), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(G183gat), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n970), .A2(new_n243), .A3(new_n797), .ZN(new_n981));
  XNOR2_X1  g780(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n982));
  AND3_X1   g781(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n982), .B1(new_n980), .B2(new_n981), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n983), .A2(new_n984), .ZN(G1350gat));
  NAND3_X1  g784(.A1(new_n970), .A2(new_n229), .A3(new_n672), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n965), .A2(new_n672), .A3(new_n966), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT61), .ZN(new_n988));
  AND3_X1   g787(.A1(new_n987), .A2(new_n988), .A3(G190gat), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n988), .B1(new_n987), .B2(G190gat), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n986), .B1(new_n989), .B2(new_n990), .ZN(G1351gat));
  NOR2_X1   g790(.A1(new_n783), .A2(new_n969), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n916), .A2(new_n992), .ZN(new_n993));
  NOR3_X1   g792(.A1(new_n993), .A2(G197gat), .A3(new_n774), .ZN(new_n994));
  XNOR2_X1  g793(.A(new_n994), .B(KEYINPUT125), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n952), .A2(new_n992), .ZN(new_n996));
  OAI21_X1  g795(.A(G197gat), .B1(new_n996), .B2(new_n630), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n995), .A2(new_n997), .ZN(G1352gat));
  XOR2_X1   g797(.A(KEYINPUT126), .B(G204gat), .Z(new_n999));
  NOR3_X1   g798(.A1(new_n993), .A2(new_n730), .A3(new_n999), .ZN(new_n1000));
  XNOR2_X1  g799(.A(new_n1000), .B(KEYINPUT62), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n999), .B1(new_n996), .B2(new_n730), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1001), .A2(new_n1002), .ZN(G1353gat));
  INV_X1    g802(.A(new_n993), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n1004), .A2(new_n356), .A3(new_n797), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n952), .A2(new_n797), .A3(new_n992), .ZN(new_n1006));
  AND3_X1   g805(.A1(new_n1006), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1007));
  AOI21_X1  g806(.A(KEYINPUT63), .B1(new_n1006), .B2(G211gat), .ZN(new_n1008));
  OAI21_X1  g807(.A(new_n1005), .B1(new_n1007), .B2(new_n1008), .ZN(G1354gat));
  OAI21_X1  g808(.A(G218gat), .B1(new_n996), .B2(new_n760), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n1004), .A2(new_n357), .A3(new_n672), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1010), .A2(new_n1011), .ZN(G1355gat));
endmodule


