//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 1 1 0 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n538, new_n539, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n555,
    new_n556, new_n557, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n589, new_n590, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT65), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n455), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT66), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n461), .A2(new_n463), .A3(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(G137), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n461), .A2(new_n463), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n466), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n470), .B1(G2105), .B2(new_n475), .ZN(G160));
  INV_X1    g051(.A(new_n466), .ZN(new_n477));
  XNOR2_X1  g052(.A(KEYINPUT66), .B(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n477), .B1(new_n478), .B2(KEYINPUT3), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT67), .ZN(new_n483));
  INV_X1    g058(.A(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  NOR2_X1   g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(new_n484), .B2(G112), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n483), .B(new_n487), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  XOR2_X1   g065(.A(new_n490), .B(KEYINPUT68), .Z(G162));
  NAND2_X1  g066(.A1(new_n484), .A2(G138), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n464), .A2(new_n494), .A3(new_n466), .ZN(new_n495));
  AND2_X1   g070(.A1(G126), .A2(G2105), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n464), .A2(new_n466), .A3(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n493), .B1(new_n473), .B2(new_n492), .ZN(new_n498));
  OR2_X1    g073(.A1(G102), .A2(G2105), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n499), .B(G2104), .C1(G114), .C2(new_n484), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n495), .A2(new_n497), .A3(new_n498), .A4(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  XNOR2_X1  g077(.A(KEYINPUT6), .B(G651), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT5), .B(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G88), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n503), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G50), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n505), .A2(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n509), .A2(new_n512), .ZN(G166));
  INV_X1    g088(.A(new_n505), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT7), .ZN(new_n515));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n514), .A2(G89), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  XOR2_X1   g092(.A(KEYINPUT69), .B(G51), .Z(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n507), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n504), .A2(G63), .ZN(new_n520));
  NAND3_X1  g095(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n511), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n519), .A2(new_n522), .ZN(G168));
  INV_X1    g098(.A(G90), .ZN(new_n524));
  INV_X1    g099(.A(G52), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n505), .A2(new_n524), .B1(new_n507), .B2(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(new_n511), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n526), .A2(new_n528), .ZN(G171));
  INV_X1    g104(.A(G81), .ZN(new_n530));
  INV_X1    g105(.A(G43), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n505), .A2(new_n530), .B1(new_n507), .B2(new_n531), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n504), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n511), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G860), .ZN(G153));
  NAND4_X1  g111(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g112(.A1(G1), .A2(G3), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT8), .ZN(new_n539));
  NAND4_X1  g114(.A1(G319), .A2(G483), .A3(G661), .A4(new_n539), .ZN(G188));
  INV_X1    g115(.A(new_n507), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G53), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT9), .ZN(new_n543));
  NAND2_X1  g118(.A1(G78), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(new_n504), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT71), .B(G65), .Z(new_n546));
  OAI21_X1  g121(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G651), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n505), .B(KEYINPUT70), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G91), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n543), .A2(new_n548), .A3(new_n550), .ZN(G299));
  INV_X1    g126(.A(G171), .ZN(G301));
  OR2_X1    g127(.A1(new_n519), .A2(new_n522), .ZN(G286));
  INV_X1    g128(.A(G166), .ZN(G303));
  NAND2_X1  g129(.A1(new_n549), .A2(G87), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n504), .A2(G74), .ZN(new_n556));
  AOI22_X1  g131(.A1(G49), .A2(new_n541), .B1(new_n556), .B2(G651), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(G288));
  NAND2_X1  g133(.A1(new_n549), .A2(G86), .ZN(new_n559));
  NAND2_X1  g134(.A1(G73), .A2(G543), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT72), .ZN(new_n561));
  INV_X1    g136(.A(G61), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n545), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n563), .A2(G651), .B1(new_n541), .B2(G48), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT73), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n559), .A2(KEYINPUT73), .A3(new_n564), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(G305));
  NAND2_X1  g144(.A1(G72), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G60), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n545), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n511), .B1(new_n572), .B2(KEYINPUT74), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n573), .B1(KEYINPUT74), .B2(new_n572), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n541), .A2(G47), .ZN(new_n575));
  XOR2_X1   g150(.A(KEYINPUT75), .B(G85), .Z(new_n576));
  OAI211_X1 g151(.A(new_n574), .B(new_n575), .C1(new_n505), .C2(new_n576), .ZN(G290));
  NAND2_X1  g152(.A1(G301), .A2(G868), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n504), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G54), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n579), .A2(new_n511), .B1(new_n507), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n549), .A2(G92), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT10), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n549), .A2(KEYINPUT10), .A3(G92), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n581), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n578), .B1(new_n586), .B2(G868), .ZN(G284));
  OAI21_X1  g162(.A(new_n578), .B1(new_n586), .B2(G868), .ZN(G321));
  INV_X1    g163(.A(G868), .ZN(new_n589));
  NAND2_X1  g164(.A1(G299), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n590), .B1(new_n589), .B2(G168), .ZN(G297));
  OAI21_X1  g166(.A(new_n590), .B1(new_n589), .B2(G168), .ZN(G280));
  INV_X1    g167(.A(G559), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n586), .B1(new_n593), .B2(G860), .ZN(G148));
  INV_X1    g169(.A(new_n535), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(new_n589), .ZN(new_n596));
  INV_X1    g171(.A(new_n586), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(G559), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n596), .B1(new_n598), .B2(new_n589), .ZN(G323));
  XNOR2_X1  g174(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g175(.A1(new_n478), .A2(G2105), .ZN(new_n601));
  XNOR2_X1  g176(.A(KEYINPUT3), .B(G2104), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT12), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT13), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(G2100), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n486), .A2(G135), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n481), .A2(G123), .ZN(new_n608));
  NOR2_X1   g183(.A1(G99), .A2(G2105), .ZN(new_n609));
  OAI21_X1  g184(.A(G2104), .B1(new_n484), .B2(G111), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n607), .B(new_n608), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G2096), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n606), .A2(new_n613), .ZN(G156));
  XOR2_X1   g189(.A(G2451), .B(G2454), .Z(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT16), .ZN(new_n616));
  XNOR2_X1  g191(.A(G1341), .B(G1348), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(G2443), .B(G2446), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(G2427), .B(G2438), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2430), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2435), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n624), .A2(new_n625), .A3(KEYINPUT14), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n620), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n620), .A2(new_n626), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n627), .A2(G14), .A3(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(KEYINPUT76), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT77), .Z(G401));
  XOR2_X1   g207(.A(G2084), .B(G2090), .Z(new_n633));
  XNOR2_X1  g208(.A(G2067), .B(G2678), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT78), .Z(new_n635));
  NOR2_X1   g210(.A1(G2072), .A2(G2078), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n444), .A2(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n633), .B1(new_n635), .B2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n637), .B(KEYINPUT17), .Z(new_n640));
  OAI21_X1  g215(.A(new_n639), .B1(new_n640), .B2(new_n635), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n637), .A2(new_n634), .A3(new_n633), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT18), .Z(new_n643));
  NAND3_X1  g218(.A1(new_n640), .A2(new_n635), .A3(new_n633), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n641), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(new_n612), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(G2100), .Z(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(G227));
  XOR2_X1   g223(.A(G1961), .B(G1966), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT79), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1956), .B(G2474), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n650), .A2(new_n652), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT80), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1971), .B(G1976), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n654), .A2(new_n658), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT20), .Z(new_n661));
  OAI211_X1 g236(.A(new_n659), .B(new_n661), .C1(new_n658), .C2(new_n653), .ZN(new_n662));
  INV_X1    g237(.A(G1986), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1991), .B(G1996), .ZN(new_n667));
  INV_X1    g242(.A(G1981), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n666), .A2(new_n669), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(G229));
  NOR2_X1   g247(.A1(KEYINPUT86), .A2(KEYINPUT36), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT32), .B(G1981), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(G16), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n567), .B2(new_n568), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n676), .A2(G6), .ZN(new_n678));
  OAI21_X1  g253(.A(KEYINPUT82), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NOR3_X1   g255(.A1(new_n677), .A2(KEYINPUT82), .A3(new_n678), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n675), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n681), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n683), .A2(new_n674), .A3(new_n679), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT83), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n682), .A2(new_n684), .A3(KEYINPUT83), .ZN(new_n688));
  NOR2_X1   g263(.A1(G16), .A2(G23), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT84), .Z(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G288), .B2(new_n676), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT33), .B(G1976), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n676), .A2(G22), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G166), .B2(new_n676), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G1971), .ZN(new_n697));
  NOR3_X1   g272(.A1(new_n693), .A2(new_n694), .A3(new_n697), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n687), .A2(new_n688), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(KEYINPUT85), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT85), .ZN(new_n701));
  NAND4_X1  g276(.A1(new_n687), .A2(new_n701), .A3(new_n688), .A4(new_n698), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n700), .A2(KEYINPUT34), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(KEYINPUT86), .A2(KEYINPUT36), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n676), .A2(G24), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G290), .B2(G16), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n704), .B1(new_n706), .B2(new_n663), .ZN(new_n707));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G25), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n481), .A2(G119), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n486), .A2(G131), .ZN(new_n711));
  OAI21_X1  g286(.A(KEYINPUT81), .B1(G95), .B2(G2105), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  NOR3_X1   g288(.A1(KEYINPUT81), .A2(G95), .A3(G2105), .ZN(new_n714));
  OAI221_X1 g289(.A(G2104), .B1(G107), .B2(new_n484), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n710), .A2(new_n711), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n709), .B1(new_n717), .B2(new_n708), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT35), .B(G1991), .Z(new_n719));
  XOR2_X1   g294(.A(new_n718), .B(new_n719), .Z(new_n720));
  AOI211_X1 g295(.A(new_n707), .B(new_n720), .C1(new_n663), .C2(new_n706), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n703), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(KEYINPUT34), .B1(new_n700), .B2(new_n702), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n673), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n723), .ZN(new_n725));
  INV_X1    g300(.A(new_n673), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n725), .A2(new_n726), .A3(new_n703), .A4(new_n721), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n708), .A2(G35), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G162), .B2(new_n708), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT29), .B(G2090), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n484), .A2(G103), .A3(G2104), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT25), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n602), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n734), .A2(new_n484), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT89), .Z(new_n736));
  AOI211_X1 g311(.A(new_n733), .B(new_n736), .C1(G139), .C2(new_n486), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(new_n708), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n708), .B2(G33), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(new_n442), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT24), .ZN(new_n741));
  INV_X1    g316(.A(G34), .ZN(new_n742));
  AOI21_X1  g317(.A(G29), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n741), .B2(new_n742), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G160), .B2(new_n708), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n740), .B1(G2084), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n739), .A2(new_n442), .ZN(new_n747));
  NAND3_X1  g322(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT26), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n748), .A2(new_n749), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n601), .A2(G105), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G129), .ZN(new_n753));
  INV_X1    g328(.A(G141), .ZN(new_n754));
  OAI221_X1 g329(.A(new_n752), .B1(new_n480), .B2(new_n753), .C1(new_n754), .C2(new_n485), .ZN(new_n755));
  MUX2_X1   g330(.A(G32), .B(new_n755), .S(G29), .Z(new_n756));
  XOR2_X1   g331(.A(KEYINPUT27), .B(G1996), .Z(new_n757));
  NOR2_X1   g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT90), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n676), .A2(G20), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT23), .ZN(new_n761));
  AND3_X1   g336(.A1(new_n543), .A2(new_n548), .A3(new_n550), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n762), .B2(new_n676), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT92), .B(G1956), .Z(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR4_X1   g340(.A1(new_n746), .A2(new_n747), .A3(new_n759), .A4(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(G168), .A2(new_n676), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n676), .B2(G21), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G164), .A2(new_n708), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G27), .B2(new_n708), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n769), .A2(G1966), .B1(new_n443), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n443), .B2(new_n771), .ZN(new_n773));
  INV_X1    g348(.A(G28), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n774), .A2(KEYINPUT30), .ZN(new_n775));
  AOI21_X1  g350(.A(G29), .B1(new_n774), .B2(KEYINPUT30), .ZN(new_n776));
  OR2_X1    g351(.A1(KEYINPUT31), .A2(G11), .ZN(new_n777));
  NAND2_X1  g352(.A1(KEYINPUT31), .A2(G11), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n775), .A2(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI221_X1 g354(.A(new_n779), .B1(new_n708), .B2(new_n611), .C1(new_n769), .C2(G1966), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n676), .A2(G5), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G171), .B2(new_n676), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT91), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(G1961), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n756), .A2(new_n757), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n763), .A2(new_n764), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n745), .A2(G2084), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n784), .A2(new_n785), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n783), .A2(G1961), .ZN(new_n789));
  NOR4_X1   g364(.A1(new_n773), .A2(new_n780), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n676), .A2(G4), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n586), .B2(new_n676), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(G1348), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n676), .A2(G19), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n535), .B2(new_n676), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(G1341), .Z(new_n796));
  OR2_X1    g371(.A1(G104), .A2(G2105), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n797), .B(G2104), .C1(G116), .C2(new_n484), .ZN(new_n798));
  INV_X1    g373(.A(G128), .ZN(new_n799));
  INV_X1    g374(.A(G140), .ZN(new_n800));
  OAI221_X1 g375(.A(new_n798), .B1(new_n480), .B2(new_n799), .C1(new_n800), .C2(new_n485), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(G29), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n708), .A2(G26), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT87), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT28), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(G2067), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n792), .A2(G1348), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n793), .A2(new_n796), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT88), .ZN(new_n811));
  AND4_X1   g386(.A1(new_n731), .A2(new_n766), .A3(new_n790), .A4(new_n811), .ZN(new_n812));
  AND3_X1   g387(.A1(new_n724), .A2(new_n727), .A3(new_n812), .ZN(G311));
  NAND3_X1  g388(.A1(new_n724), .A2(new_n727), .A3(new_n812), .ZN(G150));
  AND2_X1   g389(.A1(G80), .A2(G543), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n504), .B2(G67), .ZN(new_n816));
  OR3_X1    g391(.A1(new_n816), .A2(KEYINPUT93), .A3(new_n511), .ZN(new_n817));
  OAI21_X1  g392(.A(KEYINPUT93), .B1(new_n816), .B2(new_n511), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n541), .A2(G55), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n514), .A2(G93), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n817), .A2(new_n818), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(new_n595), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n595), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT38), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n586), .A2(G559), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  AND2_X1   g402(.A1(new_n827), .A2(KEYINPUT39), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n827), .A2(KEYINPUT39), .ZN(new_n829));
  NOR3_X1   g404(.A1(new_n828), .A2(new_n829), .A3(G860), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n821), .A2(G860), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT37), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n830), .A2(new_n832), .ZN(G145));
  INV_X1    g408(.A(G37), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n611), .B(G160), .Z(new_n835));
  XNOR2_X1  g410(.A(G162), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n497), .A2(new_n500), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(KEYINPUT94), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n495), .A2(new_n498), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT94), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n497), .A2(new_n841), .A3(new_n500), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n838), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n801), .B(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n755), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT95), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n737), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n845), .B(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(G130), .ZN(new_n849));
  NOR2_X1   g424(.A1(G106), .A2(G2105), .ZN(new_n850));
  OAI21_X1  g425(.A(G2104), .B1(new_n484), .B2(G118), .ZN(new_n851));
  OAI22_X1  g426(.A1(new_n480), .A2(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(G142), .B2(new_n486), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n604), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n717), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n848), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n848), .A2(new_n855), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(KEYINPUT96), .ZN(new_n859));
  INV_X1    g434(.A(new_n857), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n859), .A2(new_n860), .A3(new_n836), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n856), .A2(KEYINPUT96), .ZN(new_n862));
  OAI221_X1 g437(.A(new_n834), .B1(new_n836), .B2(new_n858), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g439(.A1(new_n821), .A2(new_n589), .ZN(new_n865));
  XOR2_X1   g440(.A(G290), .B(G288), .Z(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(KEYINPUT100), .ZN(new_n867));
  XNOR2_X1  g442(.A(G290), .B(G288), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT100), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(G305), .A2(G303), .ZN(new_n871));
  AOI21_X1  g446(.A(G166), .B1(new_n567), .B2(new_n568), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n867), .A2(new_n870), .A3(new_n873), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n866), .B(KEYINPUT100), .C1(new_n872), .C2(new_n871), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n876), .A2(KEYINPUT101), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT42), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n824), .B(KEYINPUT97), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n598), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n762), .A2(KEYINPUT98), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT98), .ZN(new_n882));
  NAND2_X1  g457(.A1(G299), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n881), .A2(new_n586), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n597), .A2(new_n882), .A3(G299), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n880), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(KEYINPUT99), .B(KEYINPUT41), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT41), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n884), .A2(new_n885), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n887), .B1(new_n880), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n878), .B(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n865), .B1(new_n895), .B2(new_n589), .ZN(G295));
  OAI21_X1  g471(.A(new_n865), .B1(new_n895), .B2(new_n589), .ZN(G331));
  INV_X1    g472(.A(KEYINPUT43), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n874), .A2(new_n875), .ZN(new_n899));
  NAND2_X1  g474(.A1(G286), .A2(G171), .ZN(new_n900));
  NAND2_X1  g475(.A1(G168), .A2(G301), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(new_n824), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n903), .B1(new_n890), .B2(new_n892), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n822), .A2(new_n823), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n902), .B(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n906), .A2(new_n886), .ZN(new_n907));
  NOR3_X1   g482(.A1(new_n899), .A2(new_n904), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n899), .B1(new_n904), .B2(new_n907), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n834), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n908), .B1(new_n910), .B2(KEYINPUT102), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT102), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n909), .A2(new_n912), .A3(new_n834), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n898), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n904), .A2(new_n907), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n834), .B1(new_n915), .B2(new_n899), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n886), .A2(new_n891), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n884), .A2(new_n885), .A3(new_n889), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(new_n906), .A3(new_n918), .ZN(new_n919));
  OR2_X1    g494(.A1(new_n919), .A2(KEYINPUT103), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n907), .B1(new_n919), .B2(KEYINPUT103), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n876), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n916), .A2(new_n922), .A3(KEYINPUT43), .ZN(new_n923));
  NOR3_X1   g498(.A1(new_n914), .A2(new_n923), .A3(KEYINPUT44), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n916), .A2(new_n922), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n925), .B1(new_n926), .B2(new_n898), .ZN(new_n927));
  OAI211_X1 g502(.A(KEYINPUT104), .B(KEYINPUT43), .C1(new_n916), .C2(new_n922), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n911), .A2(new_n898), .A3(new_n913), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n924), .B1(KEYINPUT44), .B2(new_n930), .ZN(G397));
  INV_X1    g506(.A(G1384), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT45), .B1(new_n843), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(G40), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n935), .B1(new_n475), .B2(G2105), .ZN(new_n936));
  INV_X1    g511(.A(G101), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n478), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n938), .B1(new_n479), .B2(G137), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n936), .B(KEYINPUT105), .C1(new_n939), .C2(G2105), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT105), .ZN(new_n941));
  INV_X1    g516(.A(new_n471), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n942), .B1(new_n602), .B2(G125), .ZN(new_n943));
  OAI21_X1  g518(.A(G40), .B1(new_n943), .B2(new_n484), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n941), .B1(new_n470), .B2(new_n944), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n940), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n934), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n801), .B(new_n807), .ZN(new_n948));
  OR2_X1    g523(.A1(new_n717), .A2(new_n719), .ZN(new_n949));
  INV_X1    g524(.A(G1996), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n755), .B(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n717), .A2(new_n719), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n948), .A2(new_n949), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(G290), .B(G1986), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n947), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT123), .ZN(new_n956));
  XOR2_X1   g531(.A(KEYINPUT109), .B(G8), .Z(new_n957));
  NOR2_X1   g532(.A1(G168), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n958), .A2(KEYINPUT51), .ZN(new_n959));
  INV_X1    g534(.A(G2084), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n940), .A2(new_n945), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT50), .B1(new_n843), .B2(new_n932), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n501), .A2(new_n932), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT50), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n960), .B(new_n961), .C1(new_n962), .C2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT111), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n968), .B1(new_n933), .B2(new_n946), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n932), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n839), .B1(KEYINPUT94), .B2(new_n837), .ZN(new_n971));
  AOI21_X1  g546(.A(G1384), .B1(new_n971), .B2(new_n842), .ZN(new_n972));
  OAI211_X1 g547(.A(KEYINPUT111), .B(new_n961), .C1(new_n972), .C2(KEYINPUT45), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n969), .A2(new_n970), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G1966), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n967), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n959), .B1(new_n976), .B2(new_n957), .ZN(new_n977));
  INV_X1    g552(.A(G8), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n958), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT51), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  AOI211_X1 g555(.A(new_n958), .B(new_n967), .C1(new_n974), .C2(new_n975), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n977), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT120), .ZN(new_n984));
  NAND3_X1  g559(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT107), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g562(.A1(G303), .A2(KEYINPUT107), .A3(KEYINPUT55), .A4(G8), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n989), .B1(G166), .B2(new_n978), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n987), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n843), .A2(new_n932), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n965), .B1(new_n992), .B2(new_n964), .ZN(new_n993));
  XNOR2_X1  g568(.A(KEYINPUT106), .B(G2090), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n961), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n997));
  AOI22_X1  g572(.A1(new_n940), .A2(new_n945), .B1(new_n963), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n843), .A2(KEYINPUT45), .A3(new_n932), .ZN(new_n999));
  AOI21_X1  g574(.A(G1971), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  OAI211_X1 g575(.A(G8), .B(new_n991), .C1(new_n996), .C2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT108), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n998), .A2(new_n999), .ZN(new_n1003));
  OAI22_X1  g578(.A1(new_n1003), .A2(G1971), .B1(new_n993), .B2(new_n995), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT108), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1004), .A2(new_n1005), .A3(G8), .A4(new_n991), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n957), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n555), .A2(new_n557), .A3(G1976), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1008), .B(new_n1009), .C1(new_n946), .C2(new_n992), .ZN(new_n1010));
  NAND2_X1  g585(.A1(KEYINPUT110), .A2(KEYINPUT52), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n957), .B1(new_n972), .B2(new_n961), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1011), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1013), .A2(new_n1009), .A3(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(KEYINPUT52), .A2(G1976), .ZN(new_n1016));
  NAND2_X1  g591(.A1(G288), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1012), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G86), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n564), .B1(new_n1019), .B2(new_n505), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(G1981), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n559), .A2(new_n668), .A3(new_n564), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT49), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1021), .A2(KEYINPUT49), .A3(new_n1022), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(new_n1013), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n998), .A2(new_n999), .ZN(new_n1028));
  INV_X1    g603(.A(G1971), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n992), .A2(KEYINPUT50), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n501), .A2(new_n964), .A3(new_n932), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1031), .A2(new_n961), .A3(new_n994), .A4(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n957), .B1(new_n1030), .B2(new_n1033), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1018), .B(new_n1027), .C1(new_n1034), .C2(new_n991), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n984), .B1(new_n1007), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1038), .A2(G2078), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n969), .A2(new_n970), .A3(new_n973), .A4(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g615(.A(KEYINPUT117), .B(G1961), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(new_n993), .B2(new_n946), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n998), .A2(new_n443), .A3(new_n999), .ZN(new_n1043));
  XOR2_X1   g618(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1040), .A2(new_n1042), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(G171), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(G171), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1049));
  XOR2_X1   g624(.A(KEYINPUT119), .B(G2078), .Z(new_n1050));
  NOR4_X1   g625(.A1(new_n470), .A2(new_n944), .A3(new_n1038), .A4(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n934), .A2(new_n1051), .A3(new_n999), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1049), .A2(new_n1042), .A3(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1037), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1018), .A2(new_n1027), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n991), .B1(new_n1056), .B2(new_n1008), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1058), .A2(KEYINPUT120), .A3(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n983), .A2(new_n1036), .A3(new_n1054), .A4(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1040), .A2(new_n1042), .A3(new_n1049), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT121), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1040), .A2(KEYINPUT121), .A3(new_n1049), .A4(new_n1042), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1042), .A2(new_n1045), .A3(new_n1052), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1037), .B1(new_n1067), .B2(G171), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n1066), .A2(KEYINPUT122), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT122), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n956), .B1(new_n1061), .B2(new_n1071), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1058), .A2(KEYINPUT120), .A3(new_n1059), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT120), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1074));
  NOR3_X1   g649(.A1(new_n1073), .A2(new_n1074), .A3(new_n982), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT122), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1066), .A2(KEYINPUT122), .A3(new_n1068), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1075), .A2(new_n1080), .A3(KEYINPUT123), .A4(new_n1054), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1031), .A2(new_n961), .A3(new_n1032), .ZN(new_n1082));
  XNOR2_X1  g657(.A(KEYINPUT112), .B(G1956), .ZN(new_n1083));
  XOR2_X1   g658(.A(KEYINPUT56), .B(G2072), .Z(new_n1084));
  OAI22_X1  g659(.A1(new_n1082), .A2(new_n1083), .B1(new_n1028), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT57), .B1(new_n543), .B2(KEYINPUT113), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n762), .B(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n993), .A2(new_n946), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n972), .A2(new_n961), .ZN(new_n1090));
  OAI22_X1  g665(.A1(new_n1089), .A2(G1348), .B1(G2067), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n586), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1088), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT114), .ZN(new_n1095));
  OR2_X1    g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n535), .A2(KEYINPUT116), .ZN(new_n1098));
  XOR2_X1   g673(.A(KEYINPUT115), .B(G1996), .Z(new_n1099));
  NAND2_X1  g674(.A1(new_n1003), .A2(new_n1099), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT58), .B(G1341), .Z(new_n1101));
  NAND2_X1  g676(.A1(new_n1090), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1098), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  XOR2_X1   g678(.A(new_n1103), .B(KEYINPUT59), .Z(new_n1104));
  INV_X1    g679(.A(KEYINPUT61), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1093), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1105), .B1(new_n1106), .B2(new_n1088), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1088), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1108), .A2(KEYINPUT61), .A3(new_n1093), .ZN(new_n1109));
  OR3_X1    g684(.A1(new_n1091), .A2(KEYINPUT60), .A3(new_n597), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1104), .A2(new_n1107), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT60), .ZN(new_n1112));
  OR2_X1    g687(.A1(new_n1091), .A2(new_n586), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1112), .B1(new_n1113), .B2(new_n1092), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1096), .B(new_n1097), .C1(new_n1111), .C2(new_n1114), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1072), .A2(new_n1081), .A3(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(G288), .A2(G1976), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1027), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1022), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1013), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1120), .B1(new_n1059), .B2(new_n1055), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n976), .A2(G286), .A3(new_n957), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1058), .A2(new_n1122), .A3(new_n1059), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT63), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n991), .B1(new_n1004), .B2(G8), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n1055), .A2(new_n1126), .A3(new_n1124), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1127), .A2(new_n1059), .A3(new_n1122), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1121), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n983), .A2(KEYINPUT62), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n982), .A2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1132), .A2(new_n1048), .A3(new_n1036), .A4(new_n1060), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT124), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1130), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n1073), .A2(new_n1074), .A3(new_n1047), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT124), .B1(new_n1136), .B2(new_n1132), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1129), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n955), .B1(new_n1116), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n948), .A2(new_n951), .ZN(new_n1140));
  OAI22_X1  g715(.A1(new_n1140), .A2(new_n952), .B1(G2067), .B2(new_n801), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n947), .ZN(new_n1142));
  INV_X1    g717(.A(new_n948), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n947), .B1(new_n1143), .B2(new_n755), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1144), .B(KEYINPUT125), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n947), .A2(new_n950), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(KEYINPUT46), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT47), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n953), .A2(new_n947), .ZN(new_n1150));
  XOR2_X1   g725(.A(new_n1150), .B(KEYINPUT126), .Z(new_n1151));
  NOR2_X1   g726(.A1(G290), .A2(G1986), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n947), .A2(new_n1152), .ZN(new_n1153));
  XOR2_X1   g728(.A(new_n1153), .B(KEYINPUT48), .Z(new_n1154));
  OAI221_X1 g729(.A(new_n1142), .B1(new_n1148), .B2(new_n1149), .C1(new_n1151), .C2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1155), .B1(new_n1149), .B2(new_n1148), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1139), .A2(new_n1156), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g732(.A1(new_n914), .A2(new_n923), .ZN(new_n1159));
  NAND3_X1  g733(.A1(new_n631), .A2(G319), .A3(new_n647), .ZN(new_n1160));
  XNOR2_X1  g734(.A(new_n1160), .B(KEYINPUT127), .ZN(new_n1161));
  OAI21_X1  g735(.A(new_n1161), .B1(new_n670), .B2(new_n671), .ZN(new_n1162));
  INV_X1    g736(.A(new_n1162), .ZN(new_n1163));
  AND3_X1   g737(.A1(new_n1159), .A2(new_n863), .A3(new_n1163), .ZN(G308));
  NAND3_X1  g738(.A1(new_n1159), .A2(new_n1163), .A3(new_n863), .ZN(G225));
endmodule


