//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 1 1 1 1 1 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 0 0 0 0 1 0 1 0 1 1 1 1 0 0 1 1 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n549, new_n550, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n600, new_n603, new_n605,
    new_n606, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1122, new_n1123, new_n1124;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT64), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT66), .Z(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(G101), .A3(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT67), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n469), .A2(new_n466), .A3(G101), .A4(G2104), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n465), .A2(G137), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n472), .B1(new_n463), .B2(new_n464), .ZN(new_n473));
  AND2_X1   g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  OAI21_X1  g049(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G112), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n465), .A2(G136), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT68), .Z(new_n482));
  AOI21_X1  g057(.A(new_n466), .B1(new_n463), .B2(new_n464), .ZN(new_n483));
  AOI211_X1 g058(.A(new_n480), .B(new_n482), .C1(G124), .C2(new_n483), .ZN(G162));
  OAI21_X1  g059(.A(KEYINPUT69), .B1(new_n466), .B2(G114), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n486));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n486), .A2(new_n487), .A3(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(KEYINPUT70), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n493));
  AOI211_X1 g068(.A(new_n493), .B(new_n490), .C1(new_n485), .C2(new_n488), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n483), .A2(G126), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NOR2_X1   g074(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n500));
  AND2_X1   g075(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n498), .B(new_n499), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT3), .B(G2104), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n499), .B1(new_n504), .B2(new_n498), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n496), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n495), .A2(new_n506), .ZN(G164));
  XNOR2_X1  g082(.A(KEYINPUT5), .B(G543), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT71), .ZN(new_n518));
  OR3_X1    g093(.A1(new_n514), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n514), .B2(new_n517), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(G166));
  NAND2_X1  g096(.A1(new_n508), .A2(G651), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n509), .A2(G543), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n523), .A2(G63), .B1(new_n524), .B2(G51), .ZN(new_n525));
  XOR2_X1   g100(.A(new_n525), .B(KEYINPUT72), .Z(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  INV_X1    g103(.A(G89), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n528), .B1(new_n510), .B2(new_n529), .ZN(new_n530));
  XOR2_X1   g105(.A(new_n530), .B(KEYINPUT73), .Z(new_n531));
  NAND2_X1  g106(.A1(new_n526), .A2(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n510), .A2(new_n534), .B1(new_n512), .B2(new_n535), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n516), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n536), .A2(new_n538), .ZN(G301));
  INV_X1    g114(.A(G301), .ZN(G171));
  AND2_X1   g115(.A1(new_n508), .A2(new_n509), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G81), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n524), .A2(G43), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  OAI211_X1 g119(.A(new_n542), .B(new_n543), .C1(new_n516), .C2(new_n544), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT74), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND4_X1  g125(.A1(G319), .A2(G483), .A3(G661), .A4(new_n550), .ZN(G188));
  NAND2_X1  g126(.A1(new_n524), .A2(G53), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT9), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n508), .A2(G65), .ZN(new_n555));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n557), .A2(G651), .B1(new_n541), .B2(G91), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(G299));
  INV_X1    g136(.A(G166), .ZN(G303));
  NAND3_X1  g137(.A1(new_n509), .A2(G49), .A3(G543), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT75), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n509), .A2(new_n565), .A3(G49), .A4(G543), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT76), .ZN(new_n568));
  NAND2_X1  g143(.A1(G74), .A2(G651), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n522), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  OAI211_X1 g145(.A(KEYINPUT76), .B(G651), .C1(new_n508), .C2(G74), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n541), .A2(G87), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n567), .A2(new_n572), .A3(new_n573), .ZN(G288));
  INV_X1    g149(.A(G86), .ZN(new_n575));
  INV_X1    g150(.A(G48), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n510), .A2(new_n575), .B1(new_n512), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n508), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n578), .A2(new_n516), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G305));
  AOI22_X1  g156(.A1(G85), .A2(new_n541), .B1(new_n524), .B2(G47), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n516), .B2(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  AND3_X1   g160(.A1(new_n508), .A2(new_n509), .A3(G92), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT10), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n508), .A2(G66), .ZN(new_n588));
  INV_X1    g163(.A(G79), .ZN(new_n589));
  INV_X1    g164(.A(G543), .ZN(new_n590));
  OAI21_X1  g165(.A(KEYINPUT77), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OR3_X1    g166(.A1(new_n589), .A2(new_n590), .A3(KEYINPUT77), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n588), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n593), .A2(G651), .B1(G54), .B2(new_n524), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n587), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n585), .B1(new_n596), .B2(G868), .ZN(G284));
  OAI21_X1  g172(.A(new_n585), .B1(new_n596), .B2(G868), .ZN(G321));
  INV_X1    g173(.A(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(G299), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(G168), .B2(new_n599), .ZN(G280));
  XNOR2_X1  g176(.A(G280), .B(KEYINPUT78), .ZN(G297));
  INV_X1    g177(.A(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n596), .B1(new_n603), .B2(G860), .ZN(G148));
  NAND2_X1  g179(.A1(new_n596), .A2(new_n603), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G868), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g182(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g183(.A1(new_n465), .A2(G135), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n483), .A2(G123), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n466), .A2(G111), .ZN(new_n611));
  OAI21_X1  g186(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n612));
  OAI211_X1 g187(.A(new_n609), .B(new_n610), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(G2096), .Z(new_n614));
  NAND3_X1  g189(.A1(new_n466), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT13), .ZN(new_n617));
  XOR2_X1   g192(.A(KEYINPUT79), .B(G2100), .Z(new_n618));
  OR2_X1    g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n617), .A2(new_n618), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n614), .A2(new_n619), .A3(new_n620), .ZN(G156));
  XNOR2_X1  g196(.A(G2427), .B(G2438), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2430), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2435), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n625), .A2(KEYINPUT14), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(G1341), .B(G1348), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n627), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2451), .B(G2454), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT81), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n631), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(G14), .A3(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(G401));
  INV_X1    g214(.A(KEYINPUT18), .ZN(new_n640));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(KEYINPUT17), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n641), .A2(new_n642), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n640), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2096), .B(G2100), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2072), .B(G2078), .Z(new_n649));
  AOI21_X1  g224(.A(new_n649), .B1(new_n643), .B2(KEYINPUT18), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT82), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n648), .B(new_n651), .ZN(G227));
  XNOR2_X1  g227(.A(G1956), .B(G2474), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT84), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1961), .B(G1966), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1971), .B(G1976), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n656), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n656), .A2(new_n660), .ZN(new_n662));
  AND2_X1   g237(.A1(new_n662), .A2(KEYINPUT20), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(KEYINPUT20), .ZN(new_n664));
  OAI221_X1 g239(.A(new_n661), .B1(new_n660), .B2(new_n657), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1981), .B(G1986), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT85), .B(KEYINPUT86), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n670));
  XNOR2_X1  g245(.A(G1991), .B(G1996), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n669), .B(new_n672), .ZN(G229));
  INV_X1    g248(.A(KEYINPUT92), .ZN(new_n674));
  NAND2_X1  g249(.A1(G288), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g250(.A1(new_n567), .A2(new_n572), .A3(KEYINPUT92), .A4(new_n573), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(G16), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n678), .B2(G23), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT33), .B(G1976), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n678), .A2(G22), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT93), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(G166), .B2(new_n678), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n686), .A2(G1971), .ZN(new_n687));
  NOR2_X1   g262(.A1(G6), .A2(G16), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(new_n580), .B2(G16), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT32), .B(G1981), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT90), .B(KEYINPUT91), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n689), .B(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(G1971), .B2(new_n686), .ZN(new_n694));
  NAND4_X1  g269(.A1(new_n682), .A2(new_n683), .A3(new_n687), .A4(new_n694), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n695), .A2(KEYINPUT34), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(KEYINPUT34), .ZN(new_n697));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G25), .ZN(new_n699));
  OR2_X1    g274(.A1(G95), .A2(G2105), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n700), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT87), .ZN(new_n702));
  AOI22_X1  g277(.A1(G119), .A2(new_n483), .B1(new_n465), .B2(G131), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n699), .B1(new_n705), .B2(new_n698), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT35), .B(G1991), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT88), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n706), .B(new_n708), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n709), .A2(KEYINPUT89), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n709), .A2(KEYINPUT89), .ZN(new_n711));
  MUX2_X1   g286(.A(G24), .B(G290), .S(G16), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G1986), .ZN(new_n713));
  NOR3_X1   g288(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n696), .A2(new_n697), .A3(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT36), .Z(new_n716));
  NOR2_X1   g291(.A1(G29), .A2(G35), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G162), .B2(G29), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT100), .B(KEYINPUT29), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(G2090), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n698), .A2(G27), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT98), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G164), .B2(new_n698), .ZN(new_n724));
  INV_X1    g299(.A(G2078), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  AOI22_X1  g301(.A1(new_n720), .A2(new_n721), .B1(KEYINPUT99), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n721), .B2(new_n720), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n698), .A2(G26), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT28), .Z(new_n730));
  OAI21_X1  g305(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n731));
  INV_X1    g306(.A(G116), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(G2105), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT94), .Z(new_n734));
  NAND2_X1  g309(.A1(new_n465), .A2(G140), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n483), .A2(G128), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n730), .B1(new_n738), .B2(G29), .ZN(new_n739));
  INV_X1    g314(.A(G2067), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G1348), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n596), .A2(G16), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G4), .B2(G16), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n741), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT30), .B(G28), .ZN(new_n746));
  OR2_X1    g321(.A1(KEYINPUT31), .A2(G11), .ZN(new_n747));
  NAND2_X1  g322(.A1(KEYINPUT31), .A2(G11), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n746), .A2(new_n698), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n613), .B2(new_n698), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n678), .A2(G5), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G171), .B2(new_n678), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n750), .B1(new_n752), .B2(G1961), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n745), .B(new_n753), .C1(G1961), .C2(new_n752), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n744), .A2(new_n742), .ZN(new_n755));
  INV_X1    g330(.A(G34), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n756), .A2(KEYINPUT24), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n756), .A2(KEYINPUT24), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n698), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G160), .B2(new_n698), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G2084), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n698), .A2(G32), .ZN(new_n762));
  NAND3_X1  g337(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT96), .Z(new_n764));
  AND2_X1   g339(.A1(new_n764), .A2(KEYINPUT26), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n764), .A2(KEYINPUT26), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n465), .A2(G141), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n483), .A2(G129), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n466), .A2(G105), .A3(G2104), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NOR3_X1   g345(.A1(new_n765), .A2(new_n766), .A3(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n762), .B1(new_n771), .B2(new_n698), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT27), .B(G1996), .Z(new_n773));
  AND2_X1   g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR4_X1   g349(.A1(new_n754), .A2(new_n755), .A3(new_n761), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n698), .A2(G33), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT25), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n777), .A2(new_n778), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n779), .A2(new_n780), .B1(new_n465), .B2(G139), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n504), .A2(G127), .ZN(new_n783));
  NAND2_X1  g358(.A1(G115), .A2(G2104), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n466), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT95), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n776), .B1(new_n787), .B2(new_n698), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(G2072), .Z(new_n789));
  OAI211_X1 g364(.A(new_n775), .B(new_n789), .C1(KEYINPUT99), .C2(new_n726), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n678), .A2(G21), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G168), .B2(new_n678), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT97), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n772), .A2(new_n773), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n792), .A2(G1966), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G1966), .B2(new_n792), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n678), .A2(G19), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n546), .B2(new_n678), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(G1341), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n678), .A2(G20), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT23), .Z(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G299), .B2(G16), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1956), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n799), .B(new_n803), .C1(new_n793), .C2(new_n794), .ZN(new_n804));
  OR4_X1    g379(.A1(new_n728), .A2(new_n790), .A3(new_n796), .A4(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n716), .A2(new_n805), .ZN(G311));
  OR2_X1    g381(.A1(new_n716), .A2(new_n805), .ZN(G150));
  NAND2_X1  g382(.A1(new_n596), .A2(G559), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT103), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT38), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n541), .A2(G93), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT101), .B(G55), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n524), .A2(new_n812), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n811), .B(new_n813), .C1(new_n516), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n546), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(KEYINPUT102), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(new_n545), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n810), .B(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT39), .ZN(new_n821));
  AOI21_X1  g396(.A(G860), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n821), .B2(new_n820), .ZN(new_n823));
  INV_X1    g398(.A(new_n817), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(G860), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT37), .Z(new_n826));
  NAND2_X1  g401(.A1(new_n823), .A2(new_n826), .ZN(G145));
  INV_X1    g402(.A(new_n786), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n738), .B(G164), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(new_n771), .ZN(new_n830));
  MUX2_X1   g405(.A(new_n787), .B(new_n828), .S(new_n830), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n704), .B(new_n616), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n483), .A2(G130), .ZN(new_n833));
  OR2_X1    g408(.A1(G106), .A2(G2105), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n834), .B(G2104), .C1(G118), .C2(new_n466), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(G142), .B2(new_n465), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n832), .B(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n831), .B(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n613), .B(new_n476), .ZN(new_n840));
  XOR2_X1   g415(.A(G162), .B(new_n840), .Z(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(G37), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n839), .A2(new_n842), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g422(.A1(new_n560), .A2(new_n595), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT104), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(G299), .A2(new_n596), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT41), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(G299), .B2(new_n596), .ZN(new_n854));
  AOI22_X1  g429(.A1(new_n852), .A2(new_n853), .B1(new_n848), .B2(new_n854), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n819), .B(new_n605), .Z(new_n856));
  OR3_X1    g431(.A1(new_n855), .A2(new_n856), .A3(KEYINPUT105), .ZN(new_n857));
  OAI21_X1  g432(.A(KEYINPUT105), .B1(new_n855), .B2(new_n856), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n851), .A2(new_n848), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n857), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT42), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n677), .B(G305), .ZN(new_n863));
  XNOR2_X1  g438(.A(G166), .B(G290), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT42), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n857), .A2(new_n858), .A3(new_n866), .A4(new_n860), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n862), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n865), .B1(new_n862), .B2(new_n867), .ZN(new_n869));
  OAI21_X1  g444(.A(G868), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n824), .A2(new_n599), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(G295));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n871), .ZN(G331));
  AOI21_X1  g448(.A(G301), .B1(new_n816), .B2(new_n818), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n816), .A2(new_n818), .A3(G301), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(G168), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n876), .ZN(new_n878));
  OAI21_X1  g453(.A(G286), .B1(new_n878), .B2(new_n874), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n877), .A2(new_n879), .A3(new_n859), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n877), .A2(new_n879), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n865), .B(new_n880), .C1(new_n881), .C2(new_n855), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n844), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT107), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT43), .ZN(new_n886));
  INV_X1    g461(.A(new_n865), .ZN(new_n887));
  INV_X1    g462(.A(new_n880), .ZN(new_n888));
  AOI21_X1  g463(.A(KEYINPUT41), .B1(new_n851), .B2(new_n848), .ZN(new_n889));
  AOI22_X1  g464(.A1(new_n850), .A2(new_n854), .B1(new_n889), .B2(KEYINPUT106), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n889), .A2(KEYINPUT106), .ZN(new_n891));
  AOI22_X1  g466(.A1(new_n877), .A2(new_n879), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n887), .B1(new_n888), .B2(new_n892), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n884), .A2(new_n885), .A3(new_n886), .A4(new_n893), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n893), .A2(new_n882), .A3(new_n886), .A4(new_n844), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(KEYINPUT107), .ZN(new_n896));
  INV_X1    g471(.A(new_n855), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n877), .A2(new_n879), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n865), .B1(new_n899), .B2(new_n880), .ZN(new_n900));
  OAI21_X1  g475(.A(KEYINPUT43), .B1(new_n883), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n894), .A2(new_n896), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n884), .A2(KEYINPUT43), .A3(new_n893), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n886), .B1(new_n883), .B2(new_n900), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT44), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n904), .A2(new_n908), .ZN(G397));
  INV_X1    g484(.A(KEYINPUT113), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n675), .A2(G1976), .A3(new_n676), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT112), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n675), .A2(KEYINPUT112), .A3(G1976), .A4(new_n676), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n490), .B1(new_n485), .B2(new_n488), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(KEYINPUT70), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n498), .B1(new_n501), .B2(new_n500), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT4), .ZN(new_n918));
  AOI22_X1  g493(.A1(new_n918), .A2(new_n502), .B1(new_n483), .B2(G126), .ZN(new_n919));
  AOI21_X1  g494(.A(G1384), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n471), .A2(new_n475), .A3(G40), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT108), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT108), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n471), .A2(new_n475), .A3(new_n923), .A4(G40), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n920), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n914), .A2(G8), .A3(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n910), .B1(new_n913), .B2(new_n926), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n925), .A2(G8), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n911), .A2(new_n912), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n928), .A2(new_n929), .A3(KEYINPUT113), .A4(new_n914), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n927), .A2(KEYINPUT52), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT45), .ZN(new_n932));
  AOI211_X1 g507(.A(new_n932), .B(G1384), .C1(new_n916), .C2(new_n919), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n918), .A2(new_n502), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n934), .B(new_n496), .C1(new_n492), .C2(new_n494), .ZN(new_n935));
  INV_X1    g510(.A(G1384), .ZN(new_n936));
  AOI21_X1  g511(.A(KEYINPUT45), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n922), .A2(new_n924), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n933), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  XNOR2_X1  g514(.A(KEYINPUT110), .B(G1971), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT50), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n920), .A2(new_n941), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n922), .A2(new_n924), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n936), .B1(new_n495), .B2(new_n506), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT50), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n942), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  OAI22_X1  g521(.A1(new_n939), .A2(new_n940), .B1(new_n946), .B2(G2090), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(G8), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n519), .A2(G8), .A3(new_n520), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n949), .B(KEYINPUT55), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(G305), .A2(G1981), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT49), .ZN(new_n953));
  INV_X1    g528(.A(G1981), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n580), .A2(new_n954), .ZN(new_n955));
  OR3_X1    g530(.A1(new_n952), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n953), .B1(new_n952), .B2(new_n955), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n956), .A2(new_n928), .A3(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(G1976), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT52), .B1(G288), .B2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n928), .A2(new_n929), .A3(new_n914), .A4(new_n960), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n931), .A2(new_n951), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT111), .B1(new_n948), .B2(new_n950), .ZN(new_n964));
  INV_X1    g539(.A(new_n950), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT111), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n965), .A2(new_n966), .A3(G8), .A4(new_n947), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n963), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(G168), .A2(G8), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n939), .A2(G1966), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT115), .ZN(new_n971));
  INV_X1    g546(.A(G2084), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n922), .B(new_n924), .C1(new_n920), .C2(new_n941), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n944), .A2(KEYINPUT50), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n970), .A2(new_n971), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT115), .B1(new_n939), .B2(G1966), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n969), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT116), .B1(new_n968), .B2(new_n978), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n931), .A2(new_n951), .A3(new_n962), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n964), .A2(new_n967), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n980), .A2(new_n978), .A3(KEYINPUT116), .A4(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT63), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n981), .A2(KEYINPUT63), .A3(new_n978), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n963), .A2(KEYINPUT117), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n963), .A2(KEYINPUT117), .ZN(new_n988));
  OAI22_X1  g563(.A1(new_n979), .A2(new_n984), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(G288), .A2(G1976), .ZN(new_n990));
  XOR2_X1   g565(.A(new_n990), .B(KEYINPUT114), .Z(new_n991));
  AND2_X1   g566(.A1(new_n958), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n928), .B1(new_n992), .B2(new_n952), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n931), .A2(new_n962), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n993), .B1(new_n981), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT62), .ZN(new_n996));
  AOI21_X1  g571(.A(G168), .B1(new_n976), .B2(new_n977), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n975), .A2(new_n972), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n944), .A2(new_n932), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n935), .A2(KEYINPUT45), .A3(new_n936), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n943), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G1966), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1001), .A2(new_n971), .A3(new_n1002), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n977), .A2(new_n998), .A3(G168), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(G8), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT51), .B1(new_n997), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1004), .A2(new_n1007), .A3(G8), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n996), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT118), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n946), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G1961), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n941), .B1(new_n935), .B2(new_n936), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1013), .A2(new_n938), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1014), .A2(KEYINPUT118), .A3(new_n942), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1011), .A2(new_n1012), .A3(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n939), .A2(KEYINPUT53), .A3(new_n725), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT123), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1020), .B1(new_n1001), .B2(G2078), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT123), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1016), .A2(new_n1022), .A3(new_n1017), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1019), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n980), .A2(new_n1024), .A3(new_n981), .A4(G171), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1009), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1006), .A2(new_n996), .A3(new_n1008), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n995), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G1956), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1029), .B1(new_n973), .B2(new_n974), .ZN(new_n1030));
  NOR3_X1   g605(.A1(new_n554), .A2(KEYINPUT57), .A3(new_n559), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n552), .B(KEYINPUT9), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1032), .B1(new_n1033), .B2(new_n558), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT56), .B(G2072), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n943), .A2(new_n999), .A3(new_n1000), .A4(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1030), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1011), .A2(new_n742), .A3(new_n1015), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n943), .A2(new_n740), .A3(new_n920), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OR2_X1    g617(.A1(new_n1042), .A2(new_n595), .ZN(new_n1043));
  OR2_X1    g618(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1044));
  AOI21_X1  g619(.A(G1956), .B1(new_n1014), .B2(new_n942), .ZN(new_n1045));
  AND4_X1   g620(.A1(new_n943), .A2(new_n999), .A3(new_n1000), .A4(new_n1036), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1044), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1039), .B1(new_n1043), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1047), .A2(KEYINPUT61), .A3(new_n1038), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT119), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT119), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1047), .A2(new_n1051), .A3(new_n1038), .A4(KEYINPUT61), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT120), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT61), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1047), .A2(new_n1038), .ZN(new_n1056));
  XOR2_X1   g631(.A(KEYINPUT58), .B(G1341), .Z(new_n1057));
  NAND2_X1  g632(.A1(new_n925), .A2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(new_n1001), .B2(G1996), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n546), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT59), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT59), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(new_n1062), .A3(new_n546), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1055), .A2(new_n1056), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1053), .A2(new_n1054), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1054), .B1(new_n1053), .B2(new_n1064), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1040), .A2(KEYINPUT60), .A3(new_n1041), .ZN(new_n1068));
  OR3_X1    g643(.A1(new_n1068), .A2(KEYINPUT121), .A3(new_n596), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n596), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT122), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT121), .B1(new_n1068), .B2(new_n596), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT122), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1068), .A2(new_n1073), .A3(new_n596), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1069), .A2(new_n1071), .A3(new_n1072), .A4(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1075), .B1(KEYINPUT60), .B2(new_n1042), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1048), .B1(new_n1067), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1023), .A2(new_n1021), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1022), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1079));
  OAI21_X1  g654(.A(G171), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT124), .B(G2078), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n921), .A2(new_n1020), .A3(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n999), .A2(new_n1000), .A3(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1016), .A2(new_n1021), .A3(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1080), .B1(G171), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1019), .A2(G301), .A3(new_n1023), .A4(new_n1021), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT125), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1084), .A2(new_n1090), .A3(G171), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1090), .B1(new_n1084), .B2(G171), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1089), .B(KEYINPUT54), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1087), .A2(new_n968), .A3(new_n1088), .A4(new_n1093), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n989), .B(new_n1028), .C1(new_n1077), .C2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n999), .A2(new_n938), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n738), .B(G2067), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n1097), .B(KEYINPUT109), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n771), .B(G1996), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n705), .A2(new_n707), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n705), .A2(new_n707), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(G290), .B(G1986), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1096), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1095), .A2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(G290), .A2(G1986), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1096), .A2(new_n1106), .ZN(new_n1107));
  XOR2_X1   g682(.A(new_n1107), .B(KEYINPUT48), .Z(new_n1108));
  AOI21_X1  g683(.A(new_n1108), .B1(new_n1102), .B2(new_n1096), .ZN(new_n1109));
  INV_X1    g684(.A(G1996), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT46), .B1(new_n1096), .B2(new_n1110), .ZN(new_n1111));
  XOR2_X1   g686(.A(new_n1111), .B(KEYINPUT126), .Z(new_n1112));
  NAND2_X1  g687(.A1(new_n1110), .A2(KEYINPUT46), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1098), .A2(new_n771), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1112), .B1(new_n1096), .B2(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n1115), .B(KEYINPUT47), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1117));
  OAI22_X1  g692(.A1(new_n1117), .A2(new_n1100), .B1(G2067), .B2(new_n738), .ZN(new_n1118));
  AOI211_X1 g693(.A(new_n1109), .B(new_n1116), .C1(new_n1096), .C2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1105), .A2(new_n1119), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g695(.A(G319), .ZN(new_n1122));
  OR2_X1    g696(.A1(G227), .A2(new_n1122), .ZN(new_n1123));
  NOR3_X1   g697(.A1(G229), .A2(G401), .A3(new_n1123), .ZN(new_n1124));
  AND3_X1   g698(.A1(new_n902), .A2(new_n1124), .A3(new_n846), .ZN(G308));
  NAND3_X1  g699(.A1(new_n902), .A2(new_n1124), .A3(new_n846), .ZN(G225));
endmodule


