

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782;

  INV_X1 U377 ( .A(n370), .ZN(n357) );
  XNOR2_X1 U378 ( .A(n544), .B(KEYINPUT38), .ZN(n710) );
  XNOR2_X1 U379 ( .A(n467), .B(n466), .ZN(n587) );
  XNOR2_X1 U380 ( .A(n450), .B(n449), .ZN(n399) );
  XNOR2_X1 U381 ( .A(KEYINPUT70), .B(G131), .ZN(n483) );
  BUF_X1 U382 ( .A(G128), .Z(n356) );
  NAND2_X1 U383 ( .A1(n671), .A2(n584), .ZN(n382) );
  XNOR2_X2 U384 ( .A(n376), .B(KEYINPUT35), .ZN(n671) );
  XNOR2_X2 U385 ( .A(n770), .B(G146), .ZN(n385) );
  AND2_X2 U386 ( .A1(n394), .A2(n393), .ZN(n392) );
  INV_X2 U387 ( .A(KEYINPUT79), .ZN(n443) );
  NOR2_X1 U388 ( .A1(n643), .A2(n357), .ZN(n371) );
  OR2_X1 U389 ( .A1(n652), .A2(G902), .ZN(n430) );
  XNOR2_X1 U390 ( .A(n399), .B(n385), .ZN(n682) );
  AND2_X2 U391 ( .A1(n372), .A2(n418), .ZN(n374) );
  XNOR2_X2 U392 ( .A(n563), .B(KEYINPUT0), .ZN(n582) );
  AND2_X2 U393 ( .A1(n692), .A2(n693), .ZN(n701) );
  XNOR2_X2 U394 ( .A(G116), .B(G113), .ZN(n432) );
  XNOR2_X1 U395 ( .A(n405), .B(KEYINPUT104), .ZN(n669) );
  XNOR2_X1 U396 ( .A(n572), .B(KEYINPUT32), .ZN(n577) );
  XNOR2_X1 U397 ( .A(n591), .B(KEYINPUT31), .ZN(n751) );
  NOR2_X1 U398 ( .A1(n583), .A2(n590), .ZN(n591) );
  OR2_X1 U399 ( .A1(n507), .A2(n452), .ZN(n458) );
  XNOR2_X1 U400 ( .A(n504), .B(n424), .ZN(n770) );
  XNOR2_X1 U401 ( .A(n483), .B(n425), .ZN(n424) );
  XNOR2_X1 U402 ( .A(n525), .B(G134), .ZN(n504) );
  XNOR2_X1 U403 ( .A(KEYINPUT4), .B(G137), .ZN(n425) );
  NAND2_X1 U404 ( .A1(n390), .A2(n392), .ZN(n358) );
  NAND2_X1 U405 ( .A1(n390), .A2(n392), .ZN(n718) );
  OR2_X1 U406 ( .A1(n581), .A2(n391), .ZN(n390) );
  XNOR2_X2 U407 ( .A(n762), .B(n446), .ZN(n519) );
  XNOR2_X2 U408 ( .A(n445), .B(n444), .ZN(n762) );
  INV_X1 U409 ( .A(G237), .ZN(n441) );
  NAND2_X1 U410 ( .A1(n383), .A2(n364), .ZN(n380) );
  NOR2_X1 U411 ( .A1(n669), .A2(KEYINPUT105), .ZN(n403) );
  XNOR2_X1 U412 ( .A(n589), .B(n387), .ZN(n602) );
  INV_X1 U413 ( .A(KEYINPUT106), .ZN(n387) );
  NOR2_X1 U414 ( .A1(n359), .A2(n362), .ZN(n377) );
  XNOR2_X1 U415 ( .A(KEYINPUT18), .B(KEYINPUT81), .ZN(n520) );
  XOR2_X1 U416 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n436) );
  NAND2_X1 U417 ( .A1(n640), .A2(n420), .ZN(n419) );
  NAND2_X1 U418 ( .A1(KEYINPUT2), .A2(KEYINPUT66), .ZN(n420) );
  XNOR2_X1 U419 ( .A(KEYINPUT68), .B(G101), .ZN(n446) );
  INV_X1 U420 ( .A(KEYINPUT33), .ZN(n375) );
  XNOR2_X1 U421 ( .A(n512), .B(n511), .ZN(n564) );
  INV_X1 U422 ( .A(G902), .ZN(n510) );
  NOR2_X1 U423 ( .A1(n380), .A2(n403), .ZN(n379) );
  XNOR2_X1 U424 ( .A(G107), .B(G104), .ZN(n444) );
  XNOR2_X1 U425 ( .A(n443), .B(G110), .ZN(n445) );
  AND2_X1 U426 ( .A1(n595), .A2(n365), .ZN(n428) );
  NAND2_X1 U427 ( .A1(n555), .A2(n709), .ZN(n557) );
  NAND2_X1 U428 ( .A1(n413), .A2(n363), .ZN(n412) );
  INV_X1 U429 ( .A(G469), .ZN(n400) );
  INV_X1 U430 ( .A(KEYINPUT64), .ZN(n447) );
  AND2_X1 U431 ( .A1(n597), .A2(KEYINPUT105), .ZN(n402) );
  OR2_X1 U432 ( .A1(n597), .A2(KEYINPUT105), .ZN(n384) );
  NOR2_X1 U433 ( .A1(G953), .A2(G237), .ZN(n488) );
  XNOR2_X1 U434 ( .A(G104), .B(G113), .ZN(n482) );
  XNOR2_X1 U435 ( .A(G143), .B(G122), .ZN(n484) );
  XOR2_X1 U436 ( .A(KEYINPUT95), .B(KEYINPUT11), .Z(n490) );
  XNOR2_X1 U437 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n521) );
  XNOR2_X1 U438 ( .A(n406), .B(KEYINPUT110), .ZN(n714) );
  XNOR2_X1 U439 ( .A(n385), .B(n440), .ZN(n652) );
  BUF_X1 U440 ( .A(n643), .Z(n772) );
  XOR2_X1 U441 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n459) );
  XNOR2_X1 U442 ( .A(n356), .B(G110), .ZN(n453) );
  XOR2_X1 U443 ( .A(G137), .B(G119), .Z(n454) );
  NAND2_X1 U444 ( .A1(n421), .A2(n419), .ZN(n418) );
  NAND2_X1 U445 ( .A1(n530), .A2(KEYINPUT66), .ZN(n421) );
  NAND2_X1 U446 ( .A1(n417), .A2(n409), .ZN(n422) );
  NOR2_X1 U447 ( .A1(n772), .A2(n638), .ZN(n417) );
  NAND2_X1 U448 ( .A1(G234), .A2(G237), .ZN(n472) );
  AND2_X1 U449 ( .A1(n396), .A2(n360), .ZN(n395) );
  NAND2_X1 U450 ( .A1(n583), .A2(n427), .ZN(n396) );
  XNOR2_X1 U451 ( .A(n386), .B(n442), .ZN(n547) );
  OR2_X1 U452 ( .A1(n602), .A2(n554), .ZN(n386) );
  XNOR2_X1 U453 ( .A(n498), .B(n497), .ZN(n565) );
  XOR2_X1 U454 ( .A(KEYINPUT62), .B(n652), .Z(n653) );
  XNOR2_X1 U455 ( .A(n509), .B(n508), .ZN(n665) );
  XNOR2_X1 U456 ( .A(n659), .B(n660), .ZN(n661) );
  NAND2_X1 U457 ( .A1(n648), .A2(n647), .ZN(n676) );
  INV_X1 U458 ( .A(n422), .ZN(n688) );
  XNOR2_X1 U459 ( .A(n388), .B(KEYINPUT40), .ZN(n407) );
  NAND2_X1 U460 ( .A1(n389), .A2(n744), .ZN(n388) );
  NOR2_X2 U461 ( .A1(n612), .A2(n611), .ZN(n745) );
  NOR2_X1 U462 ( .A1(n575), .A2(n693), .ZN(n433) );
  NAND2_X1 U463 ( .A1(n588), .A2(n587), .ZN(n405) );
  XNOR2_X1 U464 ( .A(n411), .B(n410), .ZN(n588) );
  INV_X1 U465 ( .A(KEYINPUT86), .ZN(n410) );
  AND2_X1 U466 ( .A1(n745), .A2(n613), .ZN(n359) );
  INV_X1 U467 ( .A(KEYINPUT66), .ZN(n423) );
  XNOR2_X1 U468 ( .A(n557), .B(n556), .ZN(n610) );
  XOR2_X1 U469 ( .A(n514), .B(KEYINPUT108), .Z(n360) );
  INV_X1 U470 ( .A(n583), .ZN(n595) );
  AND2_X1 U471 ( .A1(n639), .A2(n638), .ZN(n361) );
  XNOR2_X1 U472 ( .A(n589), .B(n366), .ZN(n586) );
  NAND2_X1 U473 ( .A1(n619), .A2(n618), .ZN(n362) );
  NOR2_X1 U474 ( .A1(n713), .A2(n690), .ZN(n363) );
  AND2_X1 U475 ( .A1(n384), .A2(n599), .ZN(n364) );
  XOR2_X1 U476 ( .A(KEYINPUT74), .B(KEYINPUT34), .Z(n365) );
  XOR2_X1 U477 ( .A(KEYINPUT102), .B(KEYINPUT6), .Z(n366) );
  XOR2_X1 U478 ( .A(KEYINPUT84), .B(KEYINPUT45), .Z(n367) );
  INV_X1 U479 ( .A(n530), .ZN(n640) );
  AND2_X1 U480 ( .A1(n638), .A2(n423), .ZN(n368) );
  AND2_X1 U481 ( .A1(n585), .A2(KEYINPUT72), .ZN(n369) );
  AND2_X1 U482 ( .A1(n640), .A2(KEYINPUT66), .ZN(n370) );
  NAND2_X1 U483 ( .A1(n371), .A2(n409), .ZN(n372) );
  NAND2_X1 U484 ( .A1(n409), .A2(n637), .ZN(n639) );
  NAND2_X1 U485 ( .A1(n374), .A2(n373), .ZN(n416) );
  NAND2_X1 U486 ( .A1(n639), .A2(n368), .ZN(n373) );
  XNOR2_X1 U487 ( .A(n378), .B(n367), .ZN(n641) );
  NAND2_X1 U488 ( .A1(n586), .A2(n375), .ZN(n391) );
  NAND2_X1 U489 ( .A1(n381), .A2(n379), .ZN(n378) );
  NOR2_X2 U490 ( .A1(n426), .A2(n429), .ZN(n376) );
  XNOR2_X1 U491 ( .A(n382), .B(n369), .ZN(n381) );
  NOR2_X1 U492 ( .A1(n587), .A2(n538), .ZN(n539) );
  NAND2_X1 U493 ( .A1(n620), .A2(n377), .ZN(n622) );
  NAND2_X1 U494 ( .A1(n669), .A2(n402), .ZN(n383) );
  INV_X1 U495 ( .A(n589), .ZN(n698) );
  INV_X1 U496 ( .A(n407), .ZN(n670) );
  INV_X1 U497 ( .A(n600), .ZN(n389) );
  NAND2_X1 U498 ( .A1(n358), .A2(n428), .ZN(n397) );
  NAND2_X1 U499 ( .A1(n580), .A2(KEYINPUT33), .ZN(n393) );
  NAND2_X1 U500 ( .A1(n581), .A2(KEYINPUT33), .ZN(n394) );
  NAND2_X1 U501 ( .A1(n397), .A2(n395), .ZN(n426) );
  XNOR2_X2 U502 ( .A(n398), .B(n400), .ZN(n605) );
  NOR2_X2 U503 ( .A1(n682), .A2(G902), .ZN(n398) );
  NAND2_X1 U504 ( .A1(n401), .A2(n577), .ZN(n578) );
  XNOR2_X1 U505 ( .A(n401), .B(G110), .ZN(G12) );
  NAND2_X1 U506 ( .A1(n576), .A2(n689), .ZN(n401) );
  XNOR2_X1 U507 ( .A(n404), .B(n664), .ZN(G51) );
  NAND2_X1 U508 ( .A1(n663), .A2(n676), .ZN(n404) );
  NOR2_X1 U509 ( .A1(n586), .A2(n693), .ZN(n434) );
  NAND2_X1 U510 ( .A1(n710), .A2(n709), .ZN(n406) );
  XNOR2_X1 U511 ( .A(n601), .B(KEYINPUT41), .ZN(n727) );
  NAND2_X1 U512 ( .A1(n408), .A2(n407), .ZN(n609) );
  INV_X1 U513 ( .A(n782), .ZN(n408) );
  XNOR2_X1 U514 ( .A(n607), .B(KEYINPUT42), .ZN(n782) );
  INV_X1 U515 ( .A(n641), .ZN(n409) );
  NAND2_X1 U516 ( .A1(n574), .A2(n434), .ZN(n411) );
  XNOR2_X2 U517 ( .A(n412), .B(n568), .ZN(n574) );
  INV_X1 U518 ( .A(n582), .ZN(n413) );
  XNOR2_X2 U519 ( .A(n414), .B(KEYINPUT65), .ZN(n678) );
  NAND2_X1 U520 ( .A1(n416), .A2(n422), .ZN(n414) );
  XNOR2_X1 U521 ( .A(n415), .B(KEYINPUT67), .ZN(n576) );
  NAND2_X1 U522 ( .A1(n574), .A2(n433), .ZN(n415) );
  XNOR2_X2 U523 ( .A(G143), .B(G128), .ZN(n525) );
  INV_X1 U524 ( .A(n365), .ZN(n427) );
  NOR2_X1 U525 ( .A1(n718), .A2(n365), .ZN(n429) );
  XNOR2_X2 U526 ( .A(n430), .B(G472), .ZN(n589) );
  XNOR2_X2 U527 ( .A(n432), .B(n431), .ZN(n518) );
  XNOR2_X2 U528 ( .A(KEYINPUT3), .B(G119), .ZN(n431) );
  NAND2_X1 U529 ( .A1(n488), .A2(G210), .ZN(n435) );
  XNOR2_X1 U530 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U531 ( .A(n437), .B(n518), .ZN(n439) );
  XNOR2_X1 U532 ( .A(n446), .B(KEYINPUT5), .ZN(n438) );
  XNOR2_X1 U533 ( .A(n439), .B(n438), .ZN(n440) );
  NAND2_X1 U534 ( .A1(n441), .A2(n510), .ZN(n531) );
  NAND2_X1 U535 ( .A1(n531), .A2(G214), .ZN(n709) );
  INV_X1 U536 ( .A(n709), .ZN(n554) );
  XNOR2_X1 U537 ( .A(KEYINPUT109), .B(KEYINPUT30), .ZN(n442) );
  INV_X1 U538 ( .A(n519), .ZN(n450) );
  XNOR2_X2 U539 ( .A(n447), .B(G953), .ZN(n773) );
  NAND2_X1 U540 ( .A1(n773), .A2(G227), .ZN(n448) );
  XNOR2_X1 U541 ( .A(n448), .B(G140), .ZN(n449) );
  NAND2_X1 U542 ( .A1(n773), .A2(G234), .ZN(n451) );
  XNOR2_X1 U543 ( .A(n451), .B(KEYINPUT8), .ZN(n507) );
  INV_X1 U544 ( .A(G221), .ZN(n452) );
  XNOR2_X1 U545 ( .A(n454), .B(n453), .ZN(n456) );
  XNOR2_X1 U546 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n455) );
  XNOR2_X1 U547 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U548 ( .A(n458), .B(n457), .ZN(n461) );
  XNOR2_X1 U549 ( .A(G146), .B(G125), .ZN(n524) );
  XNOR2_X1 U550 ( .A(n524), .B(G140), .ZN(n460) );
  XNOR2_X1 U551 ( .A(n460), .B(n459), .ZN(n493) );
  XNOR2_X1 U552 ( .A(n461), .B(n493), .ZN(n673) );
  NAND2_X1 U553 ( .A1(n673), .A2(n510), .ZN(n467) );
  XNOR2_X1 U554 ( .A(G902), .B(KEYINPUT15), .ZN(n530) );
  NAND2_X1 U555 ( .A1(n530), .A2(G234), .ZN(n463) );
  XNOR2_X1 U556 ( .A(KEYINPUT20), .B(KEYINPUT90), .ZN(n462) );
  XNOR2_X1 U557 ( .A(n463), .B(n462), .ZN(n468) );
  NAND2_X1 U558 ( .A1(G217), .A2(n468), .ZN(n465) );
  XNOR2_X1 U559 ( .A(KEYINPUT91), .B(KEYINPUT25), .ZN(n464) );
  XNOR2_X1 U560 ( .A(n465), .B(n464), .ZN(n466) );
  NAND2_X1 U561 ( .A1(n468), .A2(G221), .ZN(n470) );
  XNOR2_X1 U562 ( .A(KEYINPUT92), .B(KEYINPUT21), .ZN(n469) );
  XNOR2_X1 U563 ( .A(n470), .B(n469), .ZN(n690) );
  INV_X1 U564 ( .A(KEYINPUT14), .ZN(n471) );
  XNOR2_X1 U565 ( .A(n472), .B(n471), .ZN(n724) );
  INV_X1 U566 ( .A(n724), .ZN(n478) );
  INV_X1 U567 ( .A(G900), .ZN(n473) );
  NAND2_X1 U568 ( .A1(n473), .A2(G902), .ZN(n474) );
  OR2_X1 U569 ( .A1(n773), .A2(n474), .ZN(n476) );
  INV_X1 U570 ( .A(G953), .ZN(n475) );
  NAND2_X1 U571 ( .A1(n475), .A2(G952), .ZN(n559) );
  NAND2_X1 U572 ( .A1(n476), .A2(n559), .ZN(n477) );
  NAND2_X1 U573 ( .A1(n478), .A2(n477), .ZN(n479) );
  OR2_X1 U574 ( .A1(n690), .A2(n479), .ZN(n538) );
  INV_X1 U575 ( .A(n538), .ZN(n480) );
  AND2_X1 U576 ( .A1(n587), .A2(n480), .ZN(n481) );
  AND2_X1 U577 ( .A1(n605), .A2(n481), .ZN(n545) );
  AND2_X1 U578 ( .A1(n547), .A2(n545), .ZN(n537) );
  XNOR2_X1 U579 ( .A(n483), .B(n482), .ZN(n487) );
  XOR2_X1 U580 ( .A(KEYINPUT96), .B(KEYINPUT12), .Z(n485) );
  XNOR2_X1 U581 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U582 ( .A(n487), .B(n486), .ZN(n492) );
  NAND2_X1 U583 ( .A1(G214), .A2(n488), .ZN(n489) );
  XNOR2_X1 U584 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U585 ( .A(n492), .B(n491), .ZN(n494) );
  INV_X1 U586 ( .A(n493), .ZN(n771) );
  XNOR2_X1 U587 ( .A(n494), .B(n771), .ZN(n644) );
  NAND2_X1 U588 ( .A1(n644), .A2(n510), .ZN(n498) );
  XOR2_X1 U589 ( .A(KEYINPUT98), .B(KEYINPUT13), .Z(n496) );
  XNOR2_X1 U590 ( .A(KEYINPUT97), .B(G475), .ZN(n495) );
  XNOR2_X1 U591 ( .A(n496), .B(n495), .ZN(n497) );
  INV_X1 U592 ( .A(n565), .ZN(n513) );
  XNOR2_X1 U593 ( .A(G107), .B(G116), .ZN(n499) );
  XNOR2_X1 U594 ( .A(n499), .B(KEYINPUT100), .ZN(n503) );
  XOR2_X1 U595 ( .A(KEYINPUT9), .B(KEYINPUT99), .Z(n501) );
  XNOR2_X1 U596 ( .A(G122), .B(KEYINPUT7), .ZN(n500) );
  XNOR2_X1 U597 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U598 ( .A(n503), .B(n502), .Z(n505) );
  XNOR2_X1 U599 ( .A(n504), .B(n505), .ZN(n509) );
  INV_X1 U600 ( .A(G217), .ZN(n506) );
  OR2_X1 U601 ( .A1(n507), .A2(n506), .ZN(n508) );
  NAND2_X1 U602 ( .A1(n665), .A2(n510), .ZN(n512) );
  XNOR2_X1 U603 ( .A(G478), .B(KEYINPUT101), .ZN(n511) );
  INV_X1 U604 ( .A(n564), .ZN(n552) );
  NAND2_X1 U605 ( .A1(n513), .A2(n552), .ZN(n514) );
  XNOR2_X1 U606 ( .A(KEYINPUT77), .B(KEYINPUT16), .ZN(n516) );
  XNOR2_X1 U607 ( .A(G122), .B(KEYINPUT76), .ZN(n515) );
  XNOR2_X1 U608 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U609 ( .A(n518), .B(n517), .ZN(n764) );
  XNOR2_X1 U610 ( .A(n519), .B(n764), .ZN(n529) );
  NAND2_X1 U611 ( .A1(n773), .A2(G224), .ZN(n523) );
  XNOR2_X1 U612 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U613 ( .A(n523), .B(n522), .ZN(n527) );
  XNOR2_X1 U614 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U615 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U616 ( .A(n529), .B(n528), .ZN(n658) );
  NOR2_X1 U617 ( .A1(n658), .A2(n640), .ZN(n535) );
  NAND2_X1 U618 ( .A1(n531), .A2(G210), .ZN(n533) );
  INV_X1 U619 ( .A(KEYINPUT89), .ZN(n532) );
  XOR2_X1 U620 ( .A(n533), .B(n532), .Z(n534) );
  XNOR2_X1 U621 ( .A(n535), .B(n534), .ZN(n553) );
  BUF_X1 U622 ( .A(n553), .Z(n544) );
  INV_X1 U623 ( .A(n544), .ZN(n623) );
  AND2_X1 U624 ( .A1(n360), .A2(n623), .ZN(n536) );
  NAND2_X1 U625 ( .A1(n537), .A2(n536), .ZN(n619) );
  XNOR2_X1 U626 ( .A(n619), .B(G143), .ZN(G45) );
  XNOR2_X1 U627 ( .A(n539), .B(KEYINPUT71), .ZN(n603) );
  OR2_X1 U628 ( .A1(n552), .A2(n565), .ZN(n748) );
  INV_X1 U629 ( .A(n748), .ZN(n744) );
  NAND2_X1 U630 ( .A1(n744), .A2(n709), .ZN(n540) );
  NOR2_X1 U631 ( .A1(n603), .A2(n540), .ZN(n541) );
  AND2_X1 U632 ( .A1(n541), .A2(n586), .ZN(n624) );
  XNOR2_X2 U633 ( .A(n605), .B(KEYINPUT1), .ZN(n693) );
  INV_X1 U634 ( .A(n693), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n624), .A2(n573), .ZN(n542) );
  XNOR2_X1 U636 ( .A(n542), .B(KEYINPUT43), .ZN(n543) );
  NAND2_X1 U637 ( .A1(n543), .A2(n544), .ZN(n633) );
  XNOR2_X1 U638 ( .A(n633), .B(G140), .ZN(G42) );
  AND2_X1 U639 ( .A1(n545), .A2(n710), .ZN(n546) );
  NAND2_X1 U640 ( .A1(n547), .A2(n546), .ZN(n551) );
  XNOR2_X1 U641 ( .A(KEYINPUT85), .B(KEYINPUT39), .ZN(n549) );
  INV_X1 U642 ( .A(KEYINPUT73), .ZN(n548) );
  XNOR2_X1 U643 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U644 ( .A(n551), .B(n550), .ZN(n600) );
  NAND2_X1 U645 ( .A1(n552), .A2(n565), .ZN(n752) );
  OR2_X1 U646 ( .A1(n600), .A2(n752), .ZN(n634) );
  XNOR2_X1 U647 ( .A(n634), .B(G134), .ZN(G36) );
  INV_X1 U648 ( .A(n553), .ZN(n555) );
  XNOR2_X1 U649 ( .A(KEYINPUT80), .B(KEYINPUT19), .ZN(n556) );
  INV_X1 U650 ( .A(G898), .ZN(n765) );
  AND2_X1 U651 ( .A1(n765), .A2(G902), .ZN(n558) );
  NAND2_X1 U652 ( .A1(n558), .A2(G953), .ZN(n560) );
  AND2_X1 U653 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U654 ( .A1(n724), .A2(n561), .ZN(n562) );
  NAND2_X1 U655 ( .A1(n610), .A2(n562), .ZN(n563) );
  NAND2_X1 U656 ( .A1(n565), .A2(n564), .ZN(n567) );
  INV_X1 U657 ( .A(KEYINPUT103), .ZN(n566) );
  XNOR2_X1 U658 ( .A(n567), .B(n566), .ZN(n713) );
  XNOR2_X1 U659 ( .A(KEYINPUT75), .B(KEYINPUT22), .ZN(n568) );
  INV_X1 U660 ( .A(n586), .ZN(n580) );
  INV_X1 U661 ( .A(n587), .ZN(n689) );
  NAND2_X1 U662 ( .A1(n580), .A2(n689), .ZN(n569) );
  NOR2_X1 U663 ( .A1(n569), .A2(n573), .ZN(n570) );
  XNOR2_X1 U664 ( .A(n570), .B(KEYINPUT82), .ZN(n571) );
  NAND2_X1 U665 ( .A1(n574), .A2(n571), .ZN(n572) );
  XNOR2_X1 U666 ( .A(n577), .B(G119), .ZN(G21) );
  INV_X1 U667 ( .A(n602), .ZN(n575) );
  XNOR2_X1 U668 ( .A(n578), .B(KEYINPUT87), .ZN(n584) );
  INV_X1 U669 ( .A(n690), .ZN(n579) );
  AND2_X1 U670 ( .A1(n587), .A2(n579), .ZN(n692) );
  XNOR2_X1 U671 ( .A(n701), .B(KEYINPUT107), .ZN(n581) );
  BUF_X1 U672 ( .A(n582), .Z(n583) );
  INV_X1 U673 ( .A(KEYINPUT44), .ZN(n585) );
  NAND2_X1 U674 ( .A1(n701), .A2(n589), .ZN(n590) );
  NAND2_X1 U675 ( .A1(n698), .A2(n692), .ZN(n593) );
  INV_X1 U676 ( .A(n605), .ZN(n592) );
  NOR2_X1 U677 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U678 ( .A1(n595), .A2(n594), .ZN(n738) );
  NAND2_X1 U679 ( .A1(n751), .A2(n738), .ZN(n596) );
  AND2_X1 U680 ( .A1(n748), .A2(n752), .ZN(n715) );
  INV_X1 U681 ( .A(n715), .ZN(n614) );
  NAND2_X1 U682 ( .A1(n596), .A2(n614), .ZN(n597) );
  INV_X1 U683 ( .A(KEYINPUT72), .ZN(n598) );
  NAND2_X1 U684 ( .A1(n598), .A2(KEYINPUT44), .ZN(n599) );
  NOR2_X1 U685 ( .A1(n714), .A2(n713), .ZN(n601) );
  NOR2_X1 U686 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U687 ( .A(n604), .B(KEYINPUT28), .ZN(n606) );
  NAND2_X1 U688 ( .A1(n606), .A2(n605), .ZN(n612) );
  NOR2_X1 U689 ( .A1(n727), .A2(n612), .ZN(n607) );
  INV_X1 U690 ( .A(KEYINPUT46), .ZN(n608) );
  XNOR2_X1 U691 ( .A(n609), .B(n608), .ZN(n630) );
  INV_X1 U692 ( .A(n610), .ZN(n611) );
  NOR2_X1 U693 ( .A1(n715), .A2(KEYINPUT47), .ZN(n613) );
  OR2_X1 U694 ( .A1(KEYINPUT83), .A2(n614), .ZN(n615) );
  NAND2_X1 U695 ( .A1(n745), .A2(n615), .ZN(n616) );
  NAND2_X1 U696 ( .A1(n616), .A2(KEYINPUT47), .ZN(n620) );
  NAND2_X1 U697 ( .A1(n715), .A2(KEYINPUT47), .ZN(n617) );
  NAND2_X1 U698 ( .A1(n617), .A2(KEYINPUT83), .ZN(n618) );
  INV_X1 U699 ( .A(KEYINPUT78), .ZN(n621) );
  XNOR2_X1 U700 ( .A(n622), .B(n621), .ZN(n628) );
  NAND2_X1 U701 ( .A1(n624), .A2(n623), .ZN(n626) );
  INV_X1 U702 ( .A(KEYINPUT36), .ZN(n625) );
  XNOR2_X1 U703 ( .A(n626), .B(n625), .ZN(n627) );
  NAND2_X1 U704 ( .A1(n627), .A2(n693), .ZN(n754) );
  AND2_X1 U705 ( .A1(n628), .A2(n754), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n630), .A2(n629), .ZN(n632) );
  INV_X1 U707 ( .A(KEYINPUT48), .ZN(n631) );
  XNOR2_X1 U708 ( .A(n632), .B(n631), .ZN(n636) );
  AND2_X1 U709 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U710 ( .A1(n636), .A2(n635), .ZN(n643) );
  INV_X1 U711 ( .A(n643), .ZN(n637) );
  INV_X1 U712 ( .A(KEYINPUT2), .ZN(n638) );
  BUF_X1 U713 ( .A(n641), .Z(n642) );
  NAND2_X1 U714 ( .A1(n678), .A2(G475), .ZN(n646) );
  XOR2_X1 U715 ( .A(n644), .B(KEYINPUT59), .Z(n645) );
  XNOR2_X1 U716 ( .A(n646), .B(n645), .ZN(n649) );
  INV_X1 U717 ( .A(n773), .ZN(n648) );
  INV_X1 U718 ( .A(G952), .ZN(n647) );
  NAND2_X1 U719 ( .A1(n649), .A2(n676), .ZN(n651) );
  XOR2_X1 U720 ( .A(KEYINPUT120), .B(KEYINPUT60), .Z(n650) );
  XNOR2_X1 U721 ( .A(n651), .B(n650), .ZN(G60) );
  NAND2_X1 U722 ( .A1(n678), .A2(G472), .ZN(n654) );
  XNOR2_X1 U723 ( .A(n654), .B(n653), .ZN(n655) );
  NAND2_X1 U724 ( .A1(n655), .A2(n676), .ZN(n657) );
  XNOR2_X1 U725 ( .A(KEYINPUT88), .B(KEYINPUT63), .ZN(n656) );
  XNOR2_X1 U726 ( .A(n657), .B(n656), .ZN(G57) );
  INV_X1 U727 ( .A(KEYINPUT56), .ZN(n664) );
  NAND2_X1 U728 ( .A1(n678), .A2(G210), .ZN(n662) );
  BUF_X1 U729 ( .A(n658), .Z(n659) );
  XNOR2_X1 U730 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n660) );
  XNOR2_X1 U731 ( .A(n662), .B(n661), .ZN(n663) );
  NAND2_X1 U732 ( .A1(n678), .A2(G478), .ZN(n666) );
  XNOR2_X1 U733 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U734 ( .A1(n667), .A2(n676), .ZN(n668) );
  XNOR2_X1 U735 ( .A(n668), .B(KEYINPUT121), .ZN(G63) );
  XNOR2_X1 U736 ( .A(n669), .B(G101), .ZN(G3) );
  XOR2_X1 U737 ( .A(n670), .B(G131), .Z(G33) );
  XNOR2_X1 U738 ( .A(n671), .B(G122), .ZN(G24) );
  NAND2_X1 U739 ( .A1(n679), .A2(G217), .ZN(n675) );
  XNOR2_X1 U740 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n672) );
  XNOR2_X1 U741 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U742 ( .A(n675), .B(n674), .ZN(n677) );
  INV_X1 U743 ( .A(n676), .ZN(n686) );
  NOR2_X1 U744 ( .A1(n677), .A2(n686), .ZN(G66) );
  BUF_X1 U745 ( .A(n678), .Z(n679) );
  NAND2_X1 U746 ( .A1(n679), .A2(G469), .ZN(n685) );
  XOR2_X1 U747 ( .A(KEYINPUT119), .B(KEYINPUT118), .Z(n681) );
  XNOR2_X1 U748 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n680) );
  XNOR2_X1 U749 ( .A(n681), .B(n680), .ZN(n683) );
  XOR2_X1 U750 ( .A(n683), .B(n682), .Z(n684) );
  XNOR2_X1 U751 ( .A(n685), .B(n684), .ZN(n687) );
  NOR2_X1 U752 ( .A1(n687), .A2(n686), .ZN(G54) );
  NOR2_X1 U753 ( .A1(n361), .A2(n688), .ZN(n732) );
  AND2_X1 U754 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U755 ( .A(KEYINPUT49), .B(n691), .Z(n697) );
  NOR2_X1 U756 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U757 ( .A(KEYINPUT50), .B(n694), .Z(n695) );
  XNOR2_X1 U758 ( .A(KEYINPUT115), .B(n695), .ZN(n696) );
  NOR2_X1 U759 ( .A1(n697), .A2(n696), .ZN(n704) );
  NAND2_X1 U760 ( .A1(n704), .A2(KEYINPUT116), .ZN(n699) );
  NAND2_X1 U761 ( .A1(n699), .A2(n698), .ZN(n703) );
  NAND2_X1 U762 ( .A1(n589), .A2(KEYINPUT116), .ZN(n700) );
  OR2_X1 U763 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U764 ( .A1(n703), .A2(n702), .ZN(n706) );
  OR2_X1 U765 ( .A1(n704), .A2(KEYINPUT116), .ZN(n705) );
  NAND2_X1 U766 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U767 ( .A(KEYINPUT51), .B(n707), .ZN(n708) );
  NOR2_X1 U768 ( .A1(n708), .A2(n727), .ZN(n721) );
  NOR2_X1 U769 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U770 ( .A(KEYINPUT117), .B(n711), .Z(n712) );
  NOR2_X1 U771 ( .A1(n713), .A2(n712), .ZN(n717) );
  NOR2_X1 U772 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U773 ( .A1(n717), .A2(n716), .ZN(n719) );
  INV_X1 U774 ( .A(n358), .ZN(n726) );
  NOR2_X1 U775 ( .A1(n719), .A2(n726), .ZN(n720) );
  NOR2_X1 U776 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U777 ( .A(n722), .B(KEYINPUT52), .ZN(n723) );
  NOR2_X1 U778 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U779 ( .A1(n725), .A2(G952), .ZN(n730) );
  NOR2_X1 U780 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U781 ( .A1(n728), .A2(G953), .ZN(n729) );
  NAND2_X1 U782 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U783 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U784 ( .A(n733), .B(KEYINPUT53), .ZN(G75) );
  NOR2_X1 U785 ( .A1(n738), .A2(n748), .ZN(n735) );
  XNOR2_X1 U786 ( .A(G104), .B(KEYINPUT111), .ZN(n734) );
  XNOR2_X1 U787 ( .A(n735), .B(n734), .ZN(G6) );
  XOR2_X1 U788 ( .A(KEYINPUT112), .B(KEYINPUT26), .Z(n737) );
  XNOR2_X1 U789 ( .A(G107), .B(KEYINPUT27), .ZN(n736) );
  XNOR2_X1 U790 ( .A(n737), .B(n736), .ZN(n740) );
  NOR2_X1 U791 ( .A1(n738), .A2(n752), .ZN(n739) );
  XOR2_X1 U792 ( .A(n740), .B(n739), .Z(G9) );
  XOR2_X1 U793 ( .A(n356), .B(KEYINPUT29), .Z(n743) );
  INV_X1 U794 ( .A(n752), .ZN(n741) );
  NAND2_X1 U795 ( .A1(n745), .A2(n741), .ZN(n742) );
  XNOR2_X1 U796 ( .A(n743), .B(n742), .ZN(G30) );
  XOR2_X1 U797 ( .A(G146), .B(KEYINPUT113), .Z(n747) );
  NAND2_X1 U798 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U799 ( .A(n747), .B(n746), .ZN(G48) );
  NOR2_X1 U800 ( .A1(n748), .A2(n751), .ZN(n749) );
  XOR2_X1 U801 ( .A(KEYINPUT114), .B(n749), .Z(n750) );
  XNOR2_X1 U802 ( .A(G113), .B(n750), .ZN(G15) );
  NOR2_X1 U803 ( .A1(n752), .A2(n751), .ZN(n753) );
  XOR2_X1 U804 ( .A(G116), .B(n753), .Z(G18) );
  XOR2_X1 U805 ( .A(G125), .B(n754), .Z(n755) );
  XNOR2_X1 U806 ( .A(n755), .B(KEYINPUT37), .ZN(G27) );
  NOR2_X1 U807 ( .A1(n642), .A2(G953), .ZN(n760) );
  NAND2_X1 U808 ( .A1(G224), .A2(G953), .ZN(n756) );
  XNOR2_X1 U809 ( .A(n756), .B(KEYINPUT124), .ZN(n757) );
  XNOR2_X1 U810 ( .A(KEYINPUT61), .B(n757), .ZN(n758) );
  AND2_X1 U811 ( .A1(n758), .A2(G898), .ZN(n759) );
  NOR2_X1 U812 ( .A1(n760), .A2(n759), .ZN(n769) );
  XOR2_X1 U813 ( .A(G101), .B(KEYINPUT125), .Z(n761) );
  XNOR2_X1 U814 ( .A(n762), .B(n761), .ZN(n763) );
  XNOR2_X1 U815 ( .A(n764), .B(n763), .ZN(n767) );
  NAND2_X1 U816 ( .A1(n765), .A2(G953), .ZN(n766) );
  AND2_X1 U817 ( .A1(n767), .A2(n766), .ZN(n768) );
  XOR2_X1 U818 ( .A(n769), .B(n768), .Z(G69) );
  XNOR2_X1 U819 ( .A(n770), .B(n771), .ZN(n775) );
  XNOR2_X1 U820 ( .A(n772), .B(n775), .ZN(n774) );
  NAND2_X1 U821 ( .A1(n774), .A2(n773), .ZN(n780) );
  XNOR2_X1 U822 ( .A(n775), .B(G227), .ZN(n776) );
  XNOR2_X1 U823 ( .A(n776), .B(KEYINPUT126), .ZN(n777) );
  NAND2_X1 U824 ( .A1(n777), .A2(G900), .ZN(n778) );
  NAND2_X1 U825 ( .A1(G953), .A2(n778), .ZN(n779) );
  NAND2_X1 U826 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U827 ( .A(KEYINPUT127), .B(n781), .Z(G72) );
  XOR2_X1 U828 ( .A(n782), .B(G137), .Z(G39) );
endmodule

