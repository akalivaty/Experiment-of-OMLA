//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 0 1 0 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n872, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977, new_n978;
  INV_X1    g000(.A(G8gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n203), .A2(G1gat), .ZN(new_n204));
  AOI21_X1  g003(.A(new_n202), .B1(new_n204), .B2(KEYINPUT95), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n203), .B1(new_n206), .B2(G1gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(new_n205), .B(new_n208), .Z(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT21), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT100), .B1(G71gat), .B2(G78gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(G57gat), .B(G64gat), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G71gat), .B(G78gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n215), .B(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT101), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n217), .B(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n210), .A2(new_n211), .A3(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n217), .B(KEYINPUT101), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n209), .B1(new_n221), .B2(KEYINPUT21), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n219), .A2(new_n211), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n220), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(G127gat), .B(G155gat), .Z(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G231gat), .A2(G233gat), .ZN(new_n227));
  INV_X1    g026(.A(new_n225), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n220), .B(new_n228), .C1(new_n222), .C2(new_n223), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n226), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n227), .B1(new_n226), .B2(new_n229), .ZN(new_n232));
  XNOR2_X1  g031(.A(G183gat), .B(G211gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n233), .B(KEYINPUT20), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT102), .B(KEYINPUT19), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n234), .B(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  OR3_X1    g036(.A1(new_n231), .A2(new_n232), .A3(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n237), .B1(new_n231), .B2(new_n232), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT92), .B(G29gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G36gat), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NOR3_X1   g044(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT15), .ZN(new_n248));
  XOR2_X1   g047(.A(G43gat), .B(G50gat), .Z(new_n249));
  AOI22_X1  g048(.A1(new_n245), .A2(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n249), .A2(new_n248), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT93), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AND2_X1   g054(.A1(new_n246), .A2(KEYINPUT91), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n243), .B1(new_n246), .B2(KEYINPUT91), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n242), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(new_n251), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n250), .A2(KEYINPUT93), .A3(new_n252), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n255), .A2(KEYINPUT17), .A3(new_n259), .A4(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(KEYINPUT97), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n255), .A2(new_n259), .A3(new_n260), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT94), .B(KEYINPUT17), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G85gat), .A2(G92gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(KEYINPUT7), .ZN(new_n267));
  NAND2_X1  g066(.A1(G99gat), .A2(G106gat), .ZN(new_n268));
  INV_X1    g067(.A(G85gat), .ZN(new_n269));
  INV_X1    g068(.A(G92gat), .ZN(new_n270));
  AOI22_X1  g069(.A1(KEYINPUT8), .A2(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G99gat), .B(G106gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  XOR2_X1   g073(.A(new_n274), .B(KEYINPUT104), .Z(new_n275));
  NAND3_X1  g074(.A1(new_n262), .A2(new_n265), .A3(new_n275), .ZN(new_n276));
  AND2_X1   g075(.A1(G232gat), .A2(G233gat), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n263), .A2(new_n274), .B1(KEYINPUT41), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  XOR2_X1   g078(.A(G190gat), .B(G218gat), .Z(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n276), .A2(new_n280), .A3(new_n278), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(KEYINPUT105), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT105), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n276), .A2(new_n285), .A3(new_n280), .A4(new_n278), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n277), .A2(KEYINPUT41), .ZN(new_n287));
  XNOR2_X1  g086(.A(G134gat), .B(G162gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT103), .ZN(new_n290));
  AND2_X1   g089(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n284), .A2(new_n291), .A3(KEYINPUT103), .ZN(new_n292));
  AOI22_X1  g091(.A1(new_n284), .A2(new_n291), .B1(new_n282), .B2(new_n283), .ZN(new_n293));
  INV_X1    g092(.A(new_n289), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n240), .B(new_n292), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(G230gat), .A2(G233gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n217), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(new_n274), .ZN(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT106), .B(KEYINPUT10), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n298), .B(new_n299), .C1(new_n221), .C2(new_n274), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT107), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n221), .A2(KEYINPUT10), .A3(new_n274), .ZN(new_n302));
  AND3_X1   g101(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n301), .B1(new_n300), .B2(new_n302), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n296), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G120gat), .B(G148gat), .ZN(new_n306));
  INV_X1    g105(.A(G176gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G204gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n298), .B1(new_n221), .B2(new_n274), .ZN(new_n312));
  INV_X1    g111(.A(new_n296), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n305), .A2(new_n311), .A3(new_n315), .ZN(new_n316));
  XOR2_X1   g115(.A(new_n310), .B(KEYINPUT108), .Z(new_n317));
  AOI21_X1  g116(.A(new_n313), .B1(new_n300), .B2(new_n302), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n317), .B1(new_n318), .B2(new_n314), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n295), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G169gat), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n323), .A2(new_n307), .A3(KEYINPUT66), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT66), .B1(new_n323), .B2(new_n307), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT23), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(G169gat), .A2(G176gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT23), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n323), .A2(new_n307), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT67), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n336));
  INV_X1    g135(.A(G183gat), .ZN(new_n337));
  INV_X1    g136(.A(G190gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(new_n336), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n335), .A2(new_n336), .B1(new_n334), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT25), .B1(new_n331), .B2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT65), .B(G176gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT64), .B(G169gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT25), .B1(new_n345), .B2(KEYINPUT23), .ZN(new_n346));
  INV_X1    g145(.A(new_n340), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n347), .A2(new_n333), .B1(new_n329), .B2(new_n328), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT70), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n337), .A2(KEYINPUT27), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT27), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n352), .A2(G183gat), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n350), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(G183gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n337), .A2(KEYINPUT27), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT70), .ZN(new_n357));
  AOI21_X1  g156(.A(G190gat), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT68), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT27), .B(G183gat), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n338), .B(new_n361), .C1(new_n362), .C2(new_n360), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n358), .A2(KEYINPUT28), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT26), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n365), .B1(new_n324), .B2(new_n325), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n329), .A2(KEYINPUT26), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(new_n327), .A3(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n337), .A2(new_n338), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n342), .B(new_n349), .C1(new_n364), .C2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(G120gat), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT72), .B1(new_n373), .B2(G113gat), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT72), .ZN(new_n375));
  INV_X1    g174(.A(G113gat), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n376), .A3(G120gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT71), .B(G120gat), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n374), .B(new_n377), .C1(new_n378), .C2(new_n376), .ZN(new_n379));
  NOR2_X1   g178(.A1(G127gat), .A2(G134gat), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G127gat), .A2(G134gat), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT1), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT1), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n373), .A2(G113gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n376), .A2(G120gat), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n382), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n388), .A2(new_n380), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n379), .A2(new_n383), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n372), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT73), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n336), .B1(new_n332), .B2(KEYINPUT67), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n395), .B1(new_n347), .B2(KEYINPUT67), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n396), .A2(new_n330), .A3(new_n326), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n397), .A2(KEYINPUT25), .B1(new_n346), .B2(new_n348), .ZN(new_n398));
  INV_X1    g197(.A(new_n357), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT70), .B1(new_n355), .B2(new_n356), .ZN(new_n400));
  OAI211_X1 g199(.A(KEYINPUT28), .B(new_n338), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n363), .A2(new_n359), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n403), .A2(new_n370), .A3(new_n368), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n398), .A2(new_n404), .A3(new_n390), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n372), .A2(KEYINPUT73), .A3(new_n391), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n394), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(G227gat), .A2(G233gat), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT33), .ZN(new_n411));
  XNOR2_X1  g210(.A(G15gat), .B(G43gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(G71gat), .ZN(new_n413));
  INV_X1    g212(.A(G99gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n410), .B(KEYINPUT32), .C1(new_n411), .C2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n416), .B1(new_n410), .B2(new_n411), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n410), .A2(KEYINPUT32), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n418), .A2(KEYINPUT74), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT74), .B1(new_n418), .B2(new_n419), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n417), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n407), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT34), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n424), .A2(KEYINPUT76), .A3(new_n425), .A4(new_n408), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT76), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n394), .A2(new_n405), .A3(new_n425), .A4(new_n406), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n427), .B1(new_n428), .B2(new_n409), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  OR2_X1    g229(.A1(new_n407), .A2(KEYINPUT75), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n407), .A2(KEYINPUT75), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(new_n408), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n430), .B1(KEYINPUT34), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n423), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n418), .A2(new_n419), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT74), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n420), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n440), .A2(new_n417), .A3(new_n434), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT6), .ZN(new_n442));
  AND2_X1   g241(.A1(new_n442), .A2(KEYINPUT83), .ZN(new_n443));
  XNOR2_X1  g242(.A(G155gat), .B(G162gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(G141gat), .B(G148gat), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT2), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n444), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  XNOR2_X1  g248(.A(KEYINPUT78), .B(G155gat), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n447), .B1(new_n450), .B2(G162gat), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n446), .B1(new_n451), .B2(KEYINPUT79), .ZN(new_n452));
  INV_X1    g251(.A(G155gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT78), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT78), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(G155gat), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n456), .A3(G162gat), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n457), .A2(KEYINPUT79), .A3(KEYINPUT2), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n444), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n449), .B1(new_n452), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT4), .B1(new_n460), .B2(new_n391), .ZN(new_n461));
  INV_X1    g260(.A(new_n444), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n462), .B1(new_n451), .B2(KEYINPUT79), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n457), .A2(KEYINPUT2), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT79), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n445), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n448), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT4), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(new_n468), .A3(new_n390), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n461), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n373), .A2(KEYINPUT71), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT71), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(G120gat), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n376), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n374), .A2(new_n377), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n383), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT80), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n387), .A2(new_n389), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n478), .B1(new_n477), .B2(new_n479), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT3), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n483), .B(new_n449), .C1(new_n452), .C2(new_n459), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n471), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(G225gat), .A2(G233gat), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n487), .A2(KEYINPUT5), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n470), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n384), .B1(new_n388), .B2(new_n380), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n374), .A2(new_n377), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n473), .A2(G120gat), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n373), .A2(KEYINPUT71), .ZN(new_n493));
  OAI21_X1  g292(.A(G113gat), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n490), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n381), .A2(new_n382), .ZN(new_n496));
  XOR2_X1   g295(.A(G113gat), .B(G120gat), .Z(new_n497));
  AOI21_X1  g296(.A(new_n496), .B1(new_n497), .B2(new_n384), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT80), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n460), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n390), .B(new_n449), .C1(new_n452), .C2(new_n459), .ZN(new_n502));
  AOI211_X1 g301(.A(KEYINPUT82), .B(new_n486), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT82), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n499), .A2(new_n500), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n502), .B1(new_n505), .B2(new_n467), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n504), .B1(new_n506), .B2(new_n487), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT5), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT81), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n461), .A2(new_n469), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n502), .A2(KEYINPUT81), .A3(KEYINPUT4), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n510), .A2(new_n511), .A3(new_n485), .A4(new_n486), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n489), .B1(new_n508), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G1gat), .B(G29gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(KEYINPUT0), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(G57gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n517), .B(new_n269), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n443), .B1(new_n514), .B2(new_n519), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n512), .B(KEYINPUT5), .C1(new_n507), .C2(new_n503), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n521), .A2(new_n518), .A3(new_n489), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(new_n442), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n518), .B1(new_n521), .B2(new_n489), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n442), .B(new_n522), .C1(new_n525), .C2(KEYINPUT83), .ZN(new_n526));
  XNOR2_X1  g325(.A(G8gat), .B(G36gat), .ZN(new_n527));
  INV_X1    g326(.A(G64gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(new_n270), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(G211gat), .A2(G218gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(G211gat), .A2(G218gat), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(G197gat), .B(G204gat), .ZN(new_n535));
  AOI211_X1 g334(.A(new_n532), .B(new_n534), .C1(new_n535), .C2(KEYINPUT22), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n532), .A2(KEYINPUT22), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(new_n533), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n538), .A2(new_n535), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT29), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n372), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(G226gat), .A2(G233gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n543), .B(KEYINPUT77), .Z(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n372), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n540), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n546), .B1(new_n372), .B2(new_n541), .ZN(new_n549));
  INV_X1    g348(.A(new_n540), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n543), .B1(new_n398), .B2(new_n404), .ZN(new_n551));
  NOR3_X1   g350(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n531), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n543), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n372), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT29), .B1(new_n398), .B2(new_n404), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n555), .B(new_n540), .C1(new_n556), .C2(new_n546), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n542), .A2(new_n543), .B1(new_n372), .B2(new_n546), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n557), .B(new_n530), .C1(new_n558), .C2(new_n540), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n553), .A2(KEYINPUT30), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n557), .B1(new_n558), .B2(new_n540), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT30), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n561), .A2(new_n562), .A3(new_n531), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  AND3_X1   g363(.A1(new_n524), .A2(new_n526), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(G22gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(G228gat), .A2(G233gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n539), .B(KEYINPUT85), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n541), .B1(new_n568), .B2(new_n536), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n467), .B1(new_n569), .B2(new_n483), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n550), .B1(new_n484), .B2(new_n541), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n567), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n483), .B1(new_n540), .B2(KEYINPUT29), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n571), .B1(new_n460), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n574), .A2(G228gat), .A3(G233gat), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n566), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(G78gat), .B(G106gat), .Z(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT84), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT31), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(G50gat), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT86), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n572), .A2(new_n575), .A3(new_n566), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n577), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n572), .A2(new_n575), .A3(new_n566), .A4(new_n581), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n583), .B1(new_n577), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n436), .A2(new_n441), .A3(new_n565), .A4(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT35), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n565), .A2(new_n589), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT37), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n561), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n558), .A2(new_n540), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n550), .B1(new_n549), .B2(new_n551), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n596), .A2(KEYINPUT37), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT38), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n595), .A2(new_n598), .A3(new_n599), .A4(new_n530), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(new_n553), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n601), .B1(new_n524), .B2(new_n526), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT89), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n531), .B1(new_n561), .B2(new_n594), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n557), .B(KEYINPUT37), .C1(new_n558), .C2(new_n540), .ZN(new_n605));
  AOI211_X1 g404(.A(new_n603), .B(new_n599), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n595), .A2(new_n530), .A3(new_n605), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT89), .B1(new_n607), .B2(KEYINPUT38), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n602), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(new_n589), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n506), .A2(new_n487), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT87), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT87), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n470), .A2(new_n485), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n614), .B1(new_n615), .B2(new_n487), .ZN(new_n616));
  OAI211_X1 g415(.A(KEYINPUT39), .B(new_n613), .C1(new_n616), .C2(new_n612), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n486), .B1(new_n470), .B2(new_n485), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT39), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n519), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(KEYINPUT40), .B1(new_n617), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n564), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n617), .A2(new_n620), .A3(KEYINPUT40), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n514), .A2(new_n519), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT88), .B1(new_n622), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT88), .ZN(new_n628));
  NOR4_X1   g427(.A1(new_n625), .A2(new_n564), .A3(new_n621), .A4(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g429(.A(KEYINPUT90), .B1(new_n611), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n617), .A2(new_n620), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT40), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n634), .A2(new_n563), .A3(new_n560), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n628), .B1(new_n635), .B2(new_n625), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n622), .A2(new_n626), .A3(KEYINPUT88), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n588), .B1(new_n602), .B2(new_n609), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT90), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n593), .B1(new_n631), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT36), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n423), .A2(new_n435), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n434), .B1(new_n440), .B2(new_n417), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n436), .A2(KEYINPUT36), .A3(new_n441), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n592), .B1(new_n642), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n210), .A2(KEYINPUT96), .ZN(new_n650));
  OR2_X1    g449(.A1(new_n210), .A2(KEYINPUT96), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n262), .A2(new_n265), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(G229gat), .A2(G233gat), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n210), .A2(new_n263), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT18), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n210), .A2(new_n263), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n658), .A2(KEYINPUT98), .A3(new_n654), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n653), .B(KEYINPUT13), .Z(new_n660));
  INV_X1    g459(.A(KEYINPUT98), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n210), .A2(new_n661), .A3(new_n263), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n659), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n652), .A2(KEYINPUT18), .A3(new_n653), .A4(new_n654), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n657), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(G113gat), .B(G141gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G197gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT11), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(new_n323), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT12), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n665), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n657), .A2(new_n663), .A3(new_n670), .A4(new_n664), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  OR3_X1    g474(.A1(new_n649), .A2(KEYINPUT99), .A3(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n593), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n638), .A2(new_n640), .A3(new_n639), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n640), .B1(new_n638), .B2(new_n639), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n677), .B(new_n648), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n590), .B(KEYINPUT35), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n674), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(KEYINPUT99), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n322), .B1(new_n676), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n524), .A2(new_n526), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(G1gat), .ZN(G1324gat));
  INV_X1    g487(.A(new_n564), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n206), .A2(new_n202), .ZN(new_n690));
  NAND2_X1  g489(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n685), .A2(new_n689), .A3(new_n690), .A4(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n202), .B1(new_n685), .B2(new_n689), .ZN(new_n694));
  OAI21_X1  g493(.A(KEYINPUT42), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT42), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(G1325gat));
  NOR2_X1   g497(.A1(new_n644), .A2(new_n645), .ZN(new_n699));
  AOI21_X1  g498(.A(G15gat), .B1(new_n685), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT109), .ZN(new_n701));
  INV_X1    g500(.A(new_n647), .ZN(new_n702));
  AOI21_X1  g501(.A(KEYINPUT36), .B1(new_n436), .B2(new_n441), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n646), .A2(KEYINPUT109), .A3(new_n647), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AND2_X1   g505(.A1(new_n706), .A2(G15gat), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n700), .B1(new_n685), .B2(new_n707), .ZN(G1326gat));
  NAND2_X1  g507(.A1(new_n685), .A2(new_n588), .ZN(new_n709));
  XNOR2_X1  g508(.A(KEYINPUT43), .B(G22gat), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1327gat));
  INV_X1    g510(.A(KEYINPUT111), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n712), .B(KEYINPUT44), .C1(new_n649), .C2(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n714), .B1(new_n680), .B2(new_n681), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT111), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n681), .B1(new_n706), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n720), .A2(new_n717), .A3(new_n713), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n715), .A2(new_n718), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n320), .B(KEYINPUT110), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n675), .A2(new_n240), .A3(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n722), .A2(new_n686), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n241), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT45), .ZN(new_n727));
  INV_X1    g526(.A(new_n240), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n714), .A2(new_n320), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n683), .A2(KEYINPUT99), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n683), .A2(KEYINPUT99), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n728), .B(new_n729), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n732), .A2(new_n241), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n727), .B1(new_n733), .B2(new_n686), .ZN(new_n734));
  INV_X1    g533(.A(new_n686), .ZN(new_n735));
  NOR4_X1   g534(.A1(new_n732), .A2(KEYINPUT45), .A3(new_n735), .A4(new_n241), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n726), .B1(new_n734), .B2(new_n736), .ZN(G1328gat));
  AOI21_X1  g536(.A(new_n240), .B1(new_n676), .B2(new_n684), .ZN(new_n738));
  INV_X1    g537(.A(G36gat), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n738), .A2(new_n739), .A3(new_n689), .A4(new_n729), .ZN(new_n740));
  OR2_X1    g539(.A1(new_n740), .A2(KEYINPUT46), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(KEYINPUT46), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n722), .A2(new_n689), .A3(new_n724), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(G36gat), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n741), .A2(new_n742), .A3(new_n744), .ZN(G1329gat));
  NAND3_X1  g544(.A1(new_n722), .A2(new_n706), .A3(new_n724), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(G43gat), .ZN(new_n747));
  INV_X1    g546(.A(new_n699), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(G43gat), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n738), .A2(new_n729), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT47), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n747), .A2(KEYINPUT47), .A3(new_n750), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(G1330gat));
  NAND3_X1  g554(.A1(new_n722), .A2(new_n588), .A3(new_n724), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(G50gat), .ZN(new_n757));
  INV_X1    g556(.A(G50gat), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n738), .A2(new_n758), .A3(new_n588), .A4(new_n729), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT48), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n757), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n760), .B1(new_n757), .B2(new_n759), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n761), .A2(new_n762), .ZN(G1331gat));
  NAND2_X1  g562(.A1(new_n631), .A2(new_n641), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n764), .A2(new_n677), .A3(new_n704), .A4(new_n705), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n674), .B1(new_n765), .B2(new_n681), .ZN(new_n766));
  INV_X1    g565(.A(new_n723), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n295), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n686), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(G57gat), .ZN(G1332gat));
  INV_X1    g571(.A(KEYINPUT49), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n773), .A2(new_n528), .ZN(new_n774));
  OR4_X1    g573(.A1(KEYINPUT112), .A2(new_n769), .A3(new_n564), .A4(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n774), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n770), .A2(new_n689), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT112), .ZN(new_n778));
  AND4_X1   g577(.A1(new_n773), .A2(new_n775), .A3(new_n778), .A4(new_n528), .ZN(new_n779));
  AOI22_X1  g578(.A1(new_n775), .A2(new_n778), .B1(new_n773), .B2(new_n528), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n779), .A2(new_n780), .ZN(G1333gat));
  INV_X1    g580(.A(G71gat), .ZN(new_n782));
  XOR2_X1   g581(.A(new_n699), .B(KEYINPUT114), .Z(new_n783));
  OAI21_X1  g582(.A(new_n782), .B1(new_n769), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n766), .A2(G71gat), .A3(new_n768), .ZN(new_n785));
  INV_X1    g584(.A(new_n706), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n785), .A2(KEYINPUT113), .A3(new_n786), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n784), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT50), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n793), .B(new_n784), .C1(new_n789), .C2(new_n790), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(G1334gat));
  NAND2_X1  g594(.A1(new_n770), .A2(new_n588), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(G78gat), .ZN(G1335gat));
  INV_X1    g596(.A(new_n320), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n674), .A2(new_n240), .A3(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n722), .A2(new_n686), .A3(new_n799), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n800), .A2(KEYINPUT115), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(KEYINPUT115), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(G85gat), .A3(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n674), .A2(new_n240), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n720), .A2(new_n713), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT51), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n714), .B1(new_n765), .B2(new_n681), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n808), .A2(KEYINPUT51), .A3(new_n804), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n807), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  AND4_X1   g610(.A1(KEYINPUT51), .A2(new_n720), .A3(new_n713), .A4(new_n804), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(KEYINPUT116), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n735), .A2(G85gat), .A3(new_n798), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n811), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n803), .A2(new_n815), .ZN(G1336gat));
  NAND3_X1  g615(.A1(new_n722), .A2(new_n689), .A3(new_n799), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n817), .A2(G92gat), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n767), .A2(G92gat), .A3(new_n564), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n811), .A2(new_n813), .A3(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n809), .ZN(new_n823));
  AOI22_X1  g622(.A1(new_n817), .A2(G92gat), .B1(new_n823), .B2(new_n819), .ZN(new_n824));
  OAI22_X1  g623(.A1(new_n818), .A2(new_n822), .B1(new_n824), .B2(new_n821), .ZN(G1337gat));
  AND3_X1   g624(.A1(new_n722), .A2(new_n706), .A3(new_n799), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n813), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n699), .A2(new_n414), .A3(new_n320), .ZN(new_n828));
  OAI22_X1  g627(.A1(new_n826), .A2(new_n414), .B1(new_n827), .B2(new_n828), .ZN(G1338gat));
  NAND3_X1  g628(.A1(new_n722), .A2(new_n588), .A3(new_n799), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(G106gat), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n767), .A2(G106gat), .A3(new_n589), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT51), .B1(new_n808), .B2(new_n804), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(new_n833), .B2(new_n812), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n823), .A2(KEYINPUT117), .A3(new_n832), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n831), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT53), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n811), .A2(new_n813), .A3(new_n832), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n831), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n839), .A2(new_n842), .ZN(G1339gat));
  NOR3_X1   g642(.A1(new_n295), .A2(new_n674), .A3(new_n320), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n653), .B1(new_n652), .B2(new_n654), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n660), .B1(new_n659), .B2(new_n662), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n669), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n673), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n300), .A2(new_n313), .A3(new_n302), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n305), .A2(KEYINPUT54), .A3(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT54), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n311), .B1(new_n318), .B2(new_n851), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n850), .A2(KEYINPUT55), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT55), .B1(new_n850), .B2(new_n852), .ZN(new_n854));
  INV_X1    g653(.A(new_n316), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n713), .A2(new_n848), .A3(new_n856), .ZN(new_n857));
  AOI22_X1  g656(.A1(new_n674), .A2(new_n856), .B1(new_n848), .B2(new_n320), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n857), .B1(new_n858), .B2(new_n713), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n844), .B1(new_n859), .B2(new_n728), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n860), .A2(new_n735), .A3(new_n689), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n748), .A2(new_n588), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n675), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n376), .A2(KEYINPUT118), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n376), .A2(KEYINPUT118), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n867), .B1(new_n864), .B2(new_n865), .ZN(G1340gat));
  OAI21_X1  g667(.A(G120gat), .B1(new_n863), .B2(new_n767), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n320), .B1(new_n492), .B2(new_n493), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n869), .B1(new_n863), .B2(new_n870), .ZN(G1341gat));
  NOR2_X1   g670(.A1(new_n863), .A2(new_n728), .ZN(new_n872));
  XOR2_X1   g671(.A(new_n872), .B(G127gat), .Z(G1342gat));
  NOR2_X1   g672(.A1(new_n863), .A2(new_n714), .ZN(new_n874));
  NOR2_X1   g673(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n875));
  AND2_X1   g674(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n877), .B1(new_n874), .B2(new_n875), .ZN(G1343gat));
  INV_X1    g677(.A(KEYINPUT57), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n879), .B1(new_n860), .B2(new_n589), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n674), .A2(new_n856), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n848), .A2(new_n320), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n714), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n240), .B1(new_n884), .B2(new_n857), .ZN(new_n885));
  OAI211_X1 g684(.A(KEYINPUT57), .B(new_n588), .C1(new_n885), .C2(new_n844), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n706), .B1(new_n880), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n735), .A2(new_n689), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(G141gat), .B1(new_n889), .B2(new_n675), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n706), .A2(new_n589), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n861), .A2(new_n891), .ZN(new_n892));
  OR3_X1    g691(.A1(new_n892), .A2(G141gat), .A3(new_n675), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(KEYINPUT58), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT58), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n890), .A2(new_n896), .A3(new_n893), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(new_n897), .ZN(G1344gat));
  OR3_X1    g697(.A1(new_n892), .A2(G148gat), .A3(new_n798), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n887), .A2(new_n320), .A3(new_n888), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n900), .A2(new_n901), .A3(G148gat), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n901), .B1(new_n900), .B2(G148gat), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n899), .B1(new_n902), .B2(new_n903), .ZN(G1345gat));
  OAI21_X1  g703(.A(new_n450), .B1(new_n889), .B2(new_n728), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n728), .A2(new_n450), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n905), .B1(new_n892), .B2(new_n906), .ZN(G1346gat));
  OAI21_X1  g706(.A(G162gat), .B1(new_n889), .B2(new_n714), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n714), .A2(G162gat), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n892), .B2(new_n909), .ZN(G1347gat));
  NOR2_X1   g709(.A1(new_n686), .A2(new_n564), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n860), .A2(new_n912), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n913), .A2(new_n862), .ZN(new_n914));
  XOR2_X1   g713(.A(new_n914), .B(KEYINPUT119), .Z(new_n915));
  NOR2_X1   g714(.A1(new_n675), .A2(new_n344), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n860), .A2(new_n783), .A3(new_n912), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n589), .ZN(new_n919));
  OAI21_X1  g718(.A(G169gat), .B1(new_n919), .B2(new_n675), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n917), .A2(new_n920), .ZN(G1348gat));
  INV_X1    g720(.A(new_n919), .ZN(new_n922));
  AND3_X1   g721(.A1(new_n922), .A2(new_n343), .A3(new_n723), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n915), .A2(new_n320), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(new_n924), .B2(new_n307), .ZN(G1349gat));
  OAI21_X1  g724(.A(KEYINPUT120), .B1(new_n919), .B2(new_n728), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT120), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n918), .A2(new_n927), .A3(new_n589), .A4(new_n240), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n926), .A2(G183gat), .A3(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT121), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n728), .B1(new_n354), .B2(new_n357), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n914), .B2(new_n931), .ZN(new_n932));
  XNOR2_X1  g731(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n929), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n933), .B1(new_n929), .B2(new_n932), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n934), .A2(new_n935), .ZN(G1350gat));
  NAND3_X1  g735(.A1(new_n915), .A2(new_n338), .A3(new_n713), .ZN(new_n937));
  OAI21_X1  g736(.A(G190gat), .B1(new_n919), .B2(new_n714), .ZN(new_n938));
  XOR2_X1   g737(.A(KEYINPUT123), .B(KEYINPUT61), .Z(new_n939));
  NOR2_X1   g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n938), .A2(new_n939), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n937), .B1(new_n940), .B2(new_n941), .ZN(G1351gat));
  AOI21_X1  g741(.A(new_n713), .B1(new_n881), .B2(new_n882), .ZN(new_n943));
  AND3_X1   g742(.A1(new_n713), .A2(new_n848), .A3(new_n856), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n728), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(new_n844), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(KEYINPUT57), .B1(new_n947), .B2(new_n588), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n860), .A2(new_n879), .A3(new_n589), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OR2_X1    g749(.A1(new_n950), .A2(KEYINPUT124), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n706), .B1(new_n950), .B2(KEYINPUT124), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n951), .A2(new_n911), .A3(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(G197gat), .B1(new_n953), .B2(new_n675), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n913), .A2(new_n891), .ZN(new_n955));
  OR3_X1    g754(.A1(new_n955), .A2(G197gat), .A3(new_n675), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(G1352gat));
  OAI21_X1  g756(.A(G204gat), .B1(new_n953), .B2(new_n767), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n955), .A2(G204gat), .A3(new_n798), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT62), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(G1353gat));
  INV_X1    g760(.A(G211gat), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n913), .A2(new_n962), .A3(new_n240), .A4(new_n891), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT63), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n912), .A2(new_n728), .ZN(new_n965));
  AOI211_X1 g764(.A(new_n964), .B(new_n962), .C1(new_n887), .C2(new_n965), .ZN(new_n966));
  OAI211_X1 g765(.A(new_n786), .B(new_n965), .C1(new_n948), .C2(new_n949), .ZN(new_n967));
  AOI21_X1  g766(.A(KEYINPUT63), .B1(new_n967), .B2(G211gat), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n963), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT125), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI211_X1 g770(.A(KEYINPUT125), .B(new_n963), .C1(new_n966), .C2(new_n968), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(G1354gat));
  INV_X1    g772(.A(G218gat), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n974), .B1(new_n955), .B2(new_n714), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n975), .B(KEYINPUT126), .ZN(new_n976));
  INV_X1    g775(.A(new_n953), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n714), .A2(new_n974), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(G1355gat));
endmodule


