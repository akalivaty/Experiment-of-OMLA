//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 0 0 0 1 0 0 1 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1255,
    new_n1256, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT64), .Z(G353));
  INV_X1    g0006(.A(G97), .ZN(new_n207));
  INV_X1    g0007(.A(G107), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G87), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n202), .A2(new_n203), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n221), .A2(new_n212), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  INV_X1    g0024(.A(G238), .ZN(new_n225));
  INV_X1    g0025(.A(G87), .ZN(new_n226));
  INV_X1    g0026(.A(G250), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n224), .B1(new_n203), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n214), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n217), .B(new_n223), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n201), .A2(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n203), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n246), .B(new_n251), .Z(G351));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  AND2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  OAI211_X1 g0055(.A(G223), .B(new_n253), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  OAI211_X1 g0056(.A(G226), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G33), .A2(G87), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G1), .A3(G13), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  INV_X1    g0064(.A(G45), .ZN(new_n265));
  AOI21_X1  g0065(.A(G1), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(new_n261), .A3(G274), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n261), .A2(G232), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n263), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G169), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n270), .B1(new_n262), .B2(new_n259), .ZN(new_n275));
  INV_X1    g0075(.A(G179), .ZN(new_n276));
  AND3_X1   g0076(.A1(new_n275), .A2(KEYINPUT76), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(KEYINPUT76), .B1(new_n275), .B2(new_n276), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n274), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT8), .B(G58), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT67), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT67), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(new_n202), .A3(KEYINPUT8), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n221), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n286), .B1(new_n211), .B2(G20), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n288), .B1(new_n289), .B2(new_n284), .ZN(new_n290));
  INV_X1    g0090(.A(new_n286), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n254), .A2(new_n255), .ZN(new_n292));
  AOI21_X1  g0092(.A(KEYINPUT7), .B1(new_n292), .B2(new_n212), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT7), .ZN(new_n294));
  NOR4_X1   g0094(.A1(new_n254), .A2(new_n255), .A3(new_n294), .A4(G20), .ZN(new_n295));
  OAI21_X1  g0095(.A(G68), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(KEYINPUT75), .B1(new_n202), .B2(new_n203), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT75), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n298), .A2(G58), .A3(G68), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n297), .A2(new_n299), .A3(new_n218), .ZN(new_n300));
  NOR2_X1   g0100(.A1(G20), .A2(G33), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n300), .A2(G20), .B1(G159), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT16), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n291), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n296), .A2(KEYINPUT16), .A3(new_n302), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n290), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT18), .B1(new_n279), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT17), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT77), .ZN(new_n310));
  INV_X1    g0110(.A(G190), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n263), .A2(new_n271), .A3(new_n310), .A4(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(G200), .B2(new_n275), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n310), .B1(new_n275), .B2(new_n311), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT3), .B(G33), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n294), .B1(new_n316), .B2(G20), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n292), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n203), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n300), .A2(G20), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n301), .A2(G159), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n304), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n323), .A2(new_n286), .A3(new_n306), .ZN(new_n324));
  INV_X1    g0124(.A(new_n290), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n309), .B1(new_n315), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT76), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(new_n272), .B2(G179), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n275), .A2(KEYINPUT76), .A3(new_n276), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n329), .A2(new_n330), .B1(new_n273), .B2(new_n272), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT18), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n331), .A2(new_n332), .A3(new_n326), .ZN(new_n333));
  OAI21_X1  g0133(.A(KEYINPUT77), .B1(new_n272), .B2(G190), .ZN(new_n334));
  INV_X1    g0134(.A(G200), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n272), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n336), .A3(new_n312), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n307), .A2(KEYINPUT17), .A3(new_n337), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n308), .A2(new_n327), .A3(new_n333), .A4(new_n338), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n339), .B(KEYINPUT78), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT66), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n316), .A2(G222), .A3(new_n253), .ZN(new_n342));
  INV_X1    g0142(.A(G77), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n342), .B1(new_n343), .B2(new_n316), .ZN(new_n344));
  OAI21_X1  g0144(.A(G1698), .B1(new_n254), .B2(new_n255), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT65), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT65), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n347), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n344), .B1(G223), .B2(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n350), .A2(new_n261), .ZN(new_n351));
  INV_X1    g0151(.A(G226), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n261), .A2(new_n268), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n267), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n341), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n354), .ZN(new_n356));
  OAI211_X1 g0156(.A(KEYINPUT66), .B(new_n356), .C1(new_n350), .C2(new_n261), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n276), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n212), .A2(G33), .ZN(new_n360));
  OR2_X1    g0160(.A1(new_n284), .A2(new_n360), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n301), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n291), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n201), .B1(new_n211), .B2(G20), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n364), .B(KEYINPUT68), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n365), .A2(new_n291), .A3(new_n289), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(G50), .B2(new_n289), .ZN(new_n367));
  OR2_X1    g0167(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n355), .A2(new_n273), .A3(new_n357), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n359), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n355), .A2(G200), .A3(new_n357), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT9), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  OR3_X1    g0174(.A1(new_n363), .A2(new_n367), .A3(new_n373), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n372), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n311), .B1(new_n355), .B2(new_n357), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT10), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n374), .A2(new_n375), .ZN(new_n379));
  INV_X1    g0179(.A(new_n377), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT10), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n379), .A2(new_n380), .A3(new_n381), .A4(new_n372), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n371), .B1(new_n378), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n301), .ZN(new_n384));
  OAI22_X1  g0184(.A1(new_n280), .A2(new_n384), .B1(new_n212), .B2(new_n343), .ZN(new_n385));
  XNOR2_X1  g0185(.A(KEYINPUT15), .B(G87), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n386), .A2(new_n360), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n286), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n289), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n343), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n287), .A2(G77), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n388), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(G244), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n267), .B1(new_n393), .B2(new_n353), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n347), .B1(new_n316), .B2(G1698), .ZN(new_n395));
  INV_X1    g0195(.A(new_n348), .ZN(new_n396));
  OAI21_X1  g0196(.A(G238), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n316), .A2(G232), .A3(new_n253), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n292), .A2(G107), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n394), .B1(new_n402), .B2(new_n262), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n392), .B1(new_n403), .B2(G169), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n225), .B1(new_n346), .B2(new_n348), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n262), .B1(new_n405), .B2(new_n400), .ZN(new_n406));
  INV_X1    g0206(.A(new_n394), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n408), .A2(G179), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT69), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n335), .B1(new_n406), .B2(new_n407), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n411), .B1(new_n412), .B2(new_n392), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n408), .A2(new_n311), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n392), .B1(new_n408), .B2(G200), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n414), .B1(new_n415), .B2(KEYINPUT69), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n410), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n340), .A2(new_n383), .A3(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n384), .A2(new_n201), .ZN(new_n419));
  OAI22_X1  g0219(.A1(new_n360), .A2(new_n343), .B1(new_n212), .B2(G68), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n286), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n421), .B(KEYINPUT11), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT12), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT71), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n203), .B1(new_n423), .B2(KEYINPUT71), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n424), .B1(new_n425), .B2(new_n289), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n389), .A2(KEYINPUT71), .A3(new_n423), .A4(new_n203), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n426), .A2(new_n427), .B1(new_n287), .B2(G68), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n422), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT74), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT73), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n236), .A2(G1698), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(G226), .B2(G1698), .ZN(new_n433));
  INV_X1    g0233(.A(G33), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n433), .A2(new_n292), .B1(new_n434), .B2(new_n207), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n262), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n261), .A2(G238), .A3(new_n268), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT70), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n267), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n438), .B1(new_n267), .B2(new_n437), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n436), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT13), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT13), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n436), .B(new_n443), .C1(new_n439), .C2(new_n440), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n273), .B1(new_n442), .B2(new_n444), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT14), .ZN(new_n447));
  AOI22_X1  g0247(.A1(G179), .A2(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT14), .B1(new_n445), .B2(new_n273), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n431), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n442), .A2(new_n444), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n451), .A2(new_n447), .A3(G169), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n442), .A2(G179), .A3(new_n444), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n446), .A2(new_n447), .ZN(new_n455));
  NOR3_X1   g0255(.A1(new_n454), .A2(KEYINPUT73), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n430), .B1(new_n450), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n442), .A2(G190), .A3(new_n444), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n429), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n335), .B1(new_n442), .B2(new_n444), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT72), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n460), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT72), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n462), .A2(new_n463), .A3(new_n458), .A4(new_n429), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n457), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n418), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT81), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(new_n264), .A3(KEYINPUT5), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT5), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n470), .B1(KEYINPUT81), .B2(G41), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n265), .A2(G1), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n469), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(G257), .A3(new_n261), .ZN(new_n474));
  INV_X1    g0274(.A(G274), .ZN(new_n475));
  AND2_X1   g0275(.A1(G1), .A2(G13), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n475), .B1(new_n476), .B2(new_n260), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n477), .A2(new_n469), .A3(new_n471), .A4(new_n472), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(G244), .B(new_n253), .C1(new_n254), .C2(new_n255), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT4), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT80), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT80), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n480), .A2(new_n484), .A3(new_n481), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n316), .A2(KEYINPUT4), .A3(G244), .A4(new_n253), .ZN(new_n486));
  OAI211_X1 g0286(.A(G250), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n483), .A2(new_n485), .A3(new_n486), .A4(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n479), .B1(new_n490), .B2(new_n262), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(G190), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT6), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G97), .A2(G107), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(G97), .A2(G107), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AND2_X1   g0297(.A1(KEYINPUT79), .A2(G97), .ZN(new_n498));
  NOR2_X1   g0298(.A1(KEYINPUT79), .A2(G97), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n208), .A2(KEYINPUT6), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n497), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n502), .A2(G20), .B1(G77), .B2(new_n301), .ZN(new_n503));
  OAI21_X1  g0303(.A(G107), .B1(new_n293), .B2(new_n295), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n291), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n211), .A2(G33), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n289), .A2(new_n506), .A3(new_n221), .A4(new_n285), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G97), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n389), .A2(new_n207), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n492), .B(new_n512), .C1(new_n335), .C2(new_n491), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT82), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n490), .A2(new_n262), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n479), .A2(G179), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OR2_X1    g0317(.A1(KEYINPUT79), .A2(G97), .ZN(new_n518));
  NAND2_X1  g0318(.A1(KEYINPUT79), .A2(G97), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n501), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(KEYINPUT6), .B1(new_n209), .B2(new_n494), .ZN(new_n521));
  OAI21_X1  g0321(.A(G20), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n301), .A2(G77), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n208), .B1(new_n317), .B2(new_n318), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n286), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n526), .A2(new_n509), .A3(new_n510), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n517), .B(new_n527), .C1(G169), .C2(new_n491), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n513), .A2(new_n514), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n513), .A2(new_n528), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(KEYINPUT82), .ZN(new_n531));
  INV_X1    g0331(.A(new_n386), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n532), .A2(new_n289), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n507), .A2(new_n226), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT19), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n500), .B2(new_n360), .ZN(new_n536));
  NOR2_X1   g0336(.A1(G87), .A2(G107), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n518), .A2(new_n519), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n212), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n212), .B(G68), .C1(new_n254), .C2(new_n255), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n536), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI211_X1 g0343(.A(new_n533), .B(new_n534), .C1(new_n543), .C2(new_n286), .ZN(new_n544));
  OAI211_X1 g0344(.A(G244), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n545));
  OAI211_X1 g0345(.A(G238), .B(new_n253), .C1(new_n254), .C2(new_n255), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G116), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n262), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n472), .A2(new_n227), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n261), .A2(new_n550), .B1(new_n477), .B2(new_n472), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G200), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n549), .A2(G190), .A3(new_n551), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n544), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n552), .A2(new_n273), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n360), .B1(new_n518), .B2(new_n519), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n542), .B1(new_n557), .B2(KEYINPUT19), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n538), .A2(new_n540), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n286), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n533), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n532), .A2(KEYINPUT83), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT83), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n386), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n508), .A3(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n560), .A2(new_n561), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n549), .A2(new_n276), .A3(new_n551), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n556), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n555), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n316), .A2(G257), .A3(G1698), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n316), .A2(G250), .A3(new_n253), .ZN(new_n571));
  NAND2_X1  g0371(.A1(G33), .A2(G294), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n473), .A2(new_n261), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n573), .A2(new_n262), .B1(new_n574), .B2(G264), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n478), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n273), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n276), .A3(new_n478), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n212), .B(G87), .C1(new_n254), .C2(new_n255), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT22), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT22), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n316), .A2(new_n581), .A3(new_n212), .A4(G87), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n547), .A2(G20), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT23), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n212), .B2(G107), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n208), .A2(KEYINPUT23), .A3(G20), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n584), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n583), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT24), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT24), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n583), .A2(new_n591), .A3(new_n588), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n291), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT25), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n289), .B2(G107), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  NOR3_X1   g0396(.A1(new_n289), .A2(new_n594), .A3(G107), .ZN(new_n597));
  OAI22_X1  g0397(.A1(new_n596), .A2(new_n597), .B1(new_n208), .B2(new_n507), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n577), .B(new_n578), .C1(new_n593), .C2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n592), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n591), .B1(new_n583), .B2(new_n588), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n286), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n598), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n575), .A2(new_n311), .A3(new_n478), .ZN(new_n604));
  AOI21_X1  g0404(.A(G200), .B1(new_n575), .B2(new_n478), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n602), .B(new_n603), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n569), .A2(new_n599), .A3(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT21), .ZN(new_n608));
  OAI211_X1 g0408(.A(G264), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n609));
  OAI211_X1 g0409(.A(G257), .B(new_n253), .C1(new_n254), .C2(new_n255), .ZN(new_n610));
  INV_X1    g0410(.A(G303), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n609), .B(new_n610), .C1(new_n611), .C2(new_n316), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n262), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n473), .A2(G270), .A3(new_n261), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(new_n478), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G169), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n289), .A2(G116), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n508), .B2(G116), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n212), .B(new_n488), .C1(new_n500), .C2(G33), .ZN(new_n620));
  INV_X1    g0420(.A(G116), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n285), .A2(new_n221), .B1(G20), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT20), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n620), .A2(KEYINPUT20), .A3(new_n622), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n619), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n608), .B1(new_n616), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n615), .A2(G200), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n628), .B(new_n626), .C1(new_n311), .C2(new_n615), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n615), .A2(new_n276), .ZN(new_n630));
  INV_X1    g0430(.A(new_n625), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n618), .B1(new_n631), .B2(new_n623), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n632), .A2(KEYINPUT21), .A3(G169), .A4(new_n615), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n627), .A2(new_n629), .A3(new_n633), .A4(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n607), .A2(new_n635), .ZN(new_n636));
  AND4_X1   g0436(.A1(new_n467), .A2(new_n529), .A3(new_n531), .A4(new_n636), .ZN(G372));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n488), .B(new_n487), .C1(new_n480), .C2(new_n481), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n484), .B1(new_n480), .B2(new_n481), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n261), .B1(new_n641), .B2(new_n485), .ZN(new_n642));
  INV_X1    g0442(.A(new_n516), .ZN(new_n643));
  OAI22_X1  g0443(.A1(new_n642), .A2(new_n643), .B1(new_n505), .B2(new_n511), .ZN(new_n644));
  INV_X1    g0444(.A(new_n479), .ZN(new_n645));
  AOI21_X1  g0445(.A(G169), .B1(new_n515), .B2(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n638), .B1(new_n647), .B2(new_n569), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n555), .A2(new_n568), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n528), .A2(new_n649), .A3(KEYINPUT26), .ZN(new_n650));
  OAI21_X1  g0450(.A(KEYINPUT84), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n568), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n647), .A2(new_n569), .ZN(new_n653));
  NOR2_X1   g0453(.A1(KEYINPUT84), .A2(KEYINPUT26), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n651), .A2(KEYINPUT85), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT85), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT84), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n647), .A2(new_n569), .A3(new_n638), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT26), .B1(new_n528), .B2(new_n649), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n528), .A2(new_n649), .ZN(new_n662));
  INV_X1    g0462(.A(new_n654), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n568), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n657), .B1(new_n661), .B2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n599), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n627), .A2(new_n633), .A3(new_n634), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n513), .A2(new_n569), .A3(new_n528), .A4(new_n606), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n656), .A2(new_n665), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n467), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n308), .A2(new_n333), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n430), .ZN(new_n676));
  OAI21_X1  g0476(.A(KEYINPUT73), .B1(new_n454), .B2(new_n455), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n449), .A2(new_n431), .A3(new_n453), .A4(new_n452), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n679), .B1(new_n465), .B2(new_n410), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n327), .A2(new_n338), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n675), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n378), .A2(new_n382), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n371), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n673), .A2(new_n684), .ZN(G369));
  NAND3_X1  g0485(.A1(new_n211), .A2(new_n212), .A3(G13), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G213), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G343), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n626), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT86), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n693), .B1(new_n635), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n694), .B2(new_n635), .ZN(new_n696));
  INV_X1    g0496(.A(new_n667), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n693), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n696), .A2(G330), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n599), .A2(new_n606), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n692), .B1(new_n602), .B2(new_n603), .ZN(new_n702));
  OAI22_X1  g0502(.A1(new_n701), .A2(new_n702), .B1(new_n599), .B2(new_n692), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n666), .A2(new_n692), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n667), .A2(new_n692), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n706), .A2(new_n701), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(new_n705), .A3(new_n707), .ZN(G399));
  INV_X1    g0508(.A(new_n215), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G41), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(G1), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n500), .A2(new_n621), .A3(new_n537), .ZN(new_n713));
  OAI22_X1  g0513(.A1(new_n712), .A2(new_n713), .B1(new_n219), .B2(new_n711), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT28), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT29), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n672), .A2(new_n716), .A3(new_n692), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n659), .A2(new_n660), .A3(new_n568), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n692), .B1(new_n670), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(KEYINPUT29), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(G330), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT30), .ZN(new_n724));
  INV_X1    g0524(.A(new_n552), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n614), .A2(new_n478), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n726), .B1(new_n262), .B2(new_n612), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n725), .A2(new_n727), .A3(G179), .A4(new_n575), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n515), .A2(new_n645), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n724), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n727), .A2(G179), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n729), .A2(new_n731), .A3(new_n576), .A4(new_n552), .ZN(new_n732));
  AND3_X1   g0532(.A1(new_n575), .A2(new_n549), .A3(new_n551), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n733), .A2(new_n630), .A3(KEYINPUT30), .A4(new_n491), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n730), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n691), .ZN(new_n736));
  AOI21_X1  g0536(.A(KEYINPUT31), .B1(new_n735), .B2(new_n691), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n636), .A2(new_n529), .A3(new_n531), .A4(new_n692), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n723), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n722), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n715), .B1(new_n743), .B2(G1), .ZN(G364));
  AND2_X1   g0544(.A1(new_n212), .A2(G13), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n211), .B1(new_n745), .B2(G45), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n710), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n221), .B1(G20), .B2(new_n273), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n212), .A2(new_n276), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n752), .A2(new_n311), .A3(G200), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(G317), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(KEYINPUT33), .ZN(new_n756));
  OR2_X1    g0556(.A1(new_n755), .A2(KEYINPUT33), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n754), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n212), .A2(G179), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n759), .A2(G190), .A3(G200), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n758), .B1(new_n611), .B2(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n752), .A2(G190), .A3(new_n335), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G190), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n763), .A2(G322), .B1(new_n766), .B2(G329), .ZN(new_n767));
  INV_X1    g0567(.A(G311), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n752), .A2(new_n764), .ZN(new_n769));
  OAI211_X1 g0569(.A(new_n767), .B(new_n292), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n752), .A2(G200), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n311), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n761), .B(new_n770), .C1(G326), .C2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(G283), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n759), .A2(new_n311), .A3(G200), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT87), .ZN(new_n776));
  INV_X1    g0576(.A(G294), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n335), .A2(G190), .ZN(new_n778));
  OAI21_X1  g0578(.A(G20), .B1(new_n778), .B2(G179), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT88), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n779), .A2(new_n780), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n773), .B1(new_n774), .B2(new_n776), .C1(new_n777), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n766), .A2(G159), .ZN(new_n785));
  INV_X1    g0585(.A(new_n760), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n785), .A2(KEYINPUT32), .B1(G87), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(new_n203), .B2(new_n753), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n316), .B1(new_n769), .B2(new_n343), .C1(new_n202), .C2(new_n762), .ZN(new_n789));
  INV_X1    g0589(.A(new_n772), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n790), .A2(new_n201), .B1(new_n785), .B2(KEYINPUT32), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n783), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G97), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n792), .B(new_n794), .C1(new_n208), .C2(new_n776), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n751), .B1(new_n784), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(G13), .A2(G33), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(G20), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n750), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n709), .A2(new_n292), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n801), .A2(G355), .B1(new_n621), .B2(new_n709), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n709), .A2(new_n316), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(G45), .B2(new_n219), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n251), .A2(new_n265), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n749), .B(new_n796), .C1(new_n800), .C2(new_n806), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT89), .Z(new_n808));
  NAND2_X1  g0608(.A1(new_n696), .A2(new_n698), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n799), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n809), .A2(new_n723), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n812), .A2(new_n699), .A3(new_n749), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(G396));
  NAND2_X1  g0615(.A1(new_n672), .A2(new_n692), .ZN(new_n816));
  INV_X1    g0616(.A(new_n392), .ZN(new_n817));
  OAI211_X1 g0617(.A(KEYINPUT69), .B(new_n817), .C1(new_n403), .C2(new_n335), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n403), .A2(G190), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n818), .A2(new_n413), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n817), .A2(new_n692), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n410), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  NOR3_X1   g0623(.A1(new_n404), .A2(new_n409), .A3(new_n691), .ZN(new_n824));
  OAI21_X1  g0624(.A(KEYINPUT94), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT94), .ZN(new_n826));
  INV_X1    g0626(.A(new_n824), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n821), .B1(new_n416), .B2(new_n413), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n826), .B(new_n827), .C1(new_n828), .C2(new_n410), .ZN(new_n829));
  AND3_X1   g0629(.A1(new_n825), .A2(new_n829), .A3(KEYINPUT95), .ZN(new_n830));
  AOI21_X1  g0630(.A(KEYINPUT95), .B1(new_n825), .B2(new_n829), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n816), .A2(new_n832), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT96), .Z(new_n834));
  AND3_X1   g0634(.A1(new_n825), .A2(new_n829), .A3(new_n692), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n672), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n748), .B1(new_n837), .B2(new_n741), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n834), .A2(new_n740), .A3(new_n836), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n825), .A2(new_n829), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n797), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n750), .A2(new_n797), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n748), .B1(G77), .B2(new_n844), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n790), .A2(new_n611), .B1(new_n769), .B2(new_n621), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n753), .A2(KEYINPUT90), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n753), .A2(KEYINPUT90), .ZN(new_n848));
  OR2_X1    g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n846), .B1(new_n849), .B2(G283), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(KEYINPUT91), .Z(new_n851));
  INV_X1    g0651(.A(new_n776), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(G87), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n292), .B1(new_n760), .B2(new_n208), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT92), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n763), .A2(G294), .B1(new_n766), .B2(G311), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n794), .A2(new_n853), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  XNOR2_X1  g0657(.A(KEYINPUT93), .B(G143), .ZN(new_n858));
  INV_X1    g0658(.A(new_n769), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n763), .A2(new_n858), .B1(new_n859), .B2(G159), .ZN(new_n860));
  INV_X1    g0660(.A(G150), .ZN(new_n861));
  INV_X1    g0661(.A(G137), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n860), .B1(new_n861), .B2(new_n753), .C1(new_n862), .C2(new_n790), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n863), .B(KEYINPUT34), .Z(new_n864));
  NAND2_X1  g0664(.A1(new_n852), .A2(G68), .ZN(new_n865));
  INV_X1    g0665(.A(G132), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n316), .B1(new_n765), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(G50), .B2(new_n786), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n865), .B(new_n868), .C1(new_n202), .C2(new_n783), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n851), .A2(new_n857), .B1(new_n864), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n845), .B1(new_n870), .B2(new_n750), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n842), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n840), .A2(new_n872), .ZN(G384));
  OR2_X1    g0673(.A1(new_n502), .A2(KEYINPUT35), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n502), .A2(KEYINPUT35), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n874), .A2(G116), .A3(new_n222), .A4(new_n875), .ZN(new_n876));
  XOR2_X1   g0676(.A(new_n876), .B(KEYINPUT36), .Z(new_n877));
  NAND4_X1  g0677(.A1(new_n220), .A2(G77), .A3(new_n299), .A4(new_n297), .ZN(new_n878));
  AOI211_X1 g0678(.A(new_n211), .B(G13), .C1(new_n878), .C2(new_n247), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT39), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n307), .A2(new_n689), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n339), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n307), .B1(new_n279), .B2(new_n689), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n315), .A2(new_n326), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT37), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n689), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n326), .B1(new_n331), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT37), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n307), .A2(new_n337), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n886), .A2(new_n891), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n883), .A2(new_n892), .A3(KEYINPUT38), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT38), .B1(new_n883), .B2(new_n892), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n881), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n883), .A2(new_n892), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT38), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n883), .A2(new_n892), .A3(KEYINPUT38), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n898), .A2(KEYINPUT39), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n895), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n679), .A2(new_n692), .ZN(new_n902));
  OAI22_X1  g0702(.A1(new_n901), .A2(new_n902), .B1(new_n675), .B2(new_n887), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n824), .B1(new_n672), .B2(new_n835), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n898), .A2(new_n899), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n430), .A2(new_n691), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n457), .B2(new_n465), .ZN(new_n908));
  INV_X1    g0708(.A(new_n465), .ZN(new_n909));
  INV_X1    g0709(.A(new_n907), .ZN(new_n910));
  NOR3_X1   g0710(.A1(new_n679), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NOR3_X1   g0712(.A1(new_n904), .A2(new_n906), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n903), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n721), .A2(new_n467), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n684), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n914), .B(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT40), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n825), .A2(new_n829), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n738), .A2(new_n739), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n919), .B(new_n920), .C1(new_n893), .C2(new_n894), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n918), .B1(new_n921), .B2(new_n912), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n841), .B1(new_n739), .B2(new_n738), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n457), .A2(new_n465), .A3(new_n907), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n910), .B1(new_n679), .B2(new_n909), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n923), .A2(new_n905), .A3(new_n926), .A4(KEYINPUT40), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n922), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n467), .A2(new_n920), .ZN(new_n929));
  OAI21_X1  g0729(.A(G330), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n928), .B2(new_n929), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n917), .A2(new_n931), .B1(new_n211), .B2(new_n745), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n917), .A2(new_n931), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n880), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT97), .ZN(G367));
  NAND2_X1  g0735(.A1(new_n707), .A2(new_n705), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n513), .B(new_n528), .C1(new_n512), .C2(new_n692), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n647), .A2(new_n691), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n936), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT44), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n936), .A2(KEYINPUT44), .A3(new_n940), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT45), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n936), .B2(new_n940), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n707), .A2(new_n939), .A3(KEYINPUT45), .A4(new_n705), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n945), .A2(new_n704), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(KEYINPUT101), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n945), .A2(new_n949), .ZN(new_n952));
  INV_X1    g0752(.A(new_n704), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n706), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n707), .B(KEYINPUT102), .C1(new_n703), .C2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(KEYINPUT102), .B2(new_n707), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(new_n699), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n952), .A2(KEYINPUT101), .A3(new_n953), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n743), .A2(new_n955), .A3(new_n959), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n743), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n710), .B(KEYINPUT41), .Z(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n747), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n706), .A2(new_n701), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT42), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n939), .B(new_n966), .C1(KEYINPUT100), .C2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(KEYINPUT100), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n968), .B(new_n969), .Z(new_n970));
  XOR2_X1   g0770(.A(new_n939), .B(KEYINPUT99), .Z(new_n971));
  AOI21_X1  g0771(.A(new_n647), .B1(new_n971), .B2(new_n666), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n970), .B1(new_n972), .B2(new_n691), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n544), .A2(new_n692), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n569), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n568), .B2(new_n974), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(KEYINPUT43), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT43), .B1(new_n976), .B2(KEYINPUT98), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(KEYINPUT98), .B2(new_n976), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n973), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n973), .B2(new_n979), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n953), .A2(new_n971), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n981), .B(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n793), .A2(G68), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n861), .B2(new_n762), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT104), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n316), .B1(new_n765), .B2(new_n862), .C1(new_n201), .C2(new_n769), .ZN(new_n987));
  INV_X1    g0787(.A(new_n775), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n772), .A2(new_n858), .B1(new_n988), .B2(G77), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n202), .B2(new_n760), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n987), .B(new_n990), .C1(G159), .C2(new_n849), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n986), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT105), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n786), .A2(G116), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT46), .Z(new_n995));
  OAI22_X1  g0795(.A1(new_n790), .A2(new_n768), .B1(new_n775), .B2(new_n500), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n292), .B1(new_n769), .B2(new_n774), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n762), .A2(new_n611), .B1(new_n765), .B2(new_n755), .ZN(new_n998));
  NOR4_X1   g0798(.A1(new_n995), .A2(new_n996), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n849), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n999), .B1(new_n208), .B2(new_n783), .C1(new_n777), .C2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n993), .A2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT47), .Z(new_n1003));
  NOR2_X1   g0803(.A1(new_n1003), .A2(new_n751), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n803), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n800), .B1(new_n215), .B2(new_n386), .C1(new_n1005), .C2(new_n242), .ZN(new_n1006));
  AND2_X1   g0806(.A1(new_n1006), .A2(KEYINPUT103), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1007), .A2(new_n749), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n799), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1008), .B1(KEYINPUT103), .B2(new_n1006), .C1(new_n976), .C2(new_n1009), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n965), .A2(new_n983), .B1(new_n1004), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT106), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1011), .B(new_n1012), .ZN(G387));
  INV_X1    g0813(.A(new_n959), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n742), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n959), .A2(new_n722), .A3(new_n741), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1015), .A2(new_n710), .A3(new_n1016), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n239), .A2(new_n265), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n1018), .A2(new_n803), .B1(new_n713), .B2(new_n801), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n280), .A2(G50), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT50), .Z(new_n1021));
  OAI21_X1  g0821(.A(new_n265), .B1(new_n203), .B2(new_n343), .ZN(new_n1022));
  NOR3_X1   g0822(.A1(new_n1021), .A2(new_n713), .A3(new_n1022), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n1019), .A2(new_n1023), .B1(G107), .B2(new_n215), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n749), .B1(new_n1024), .B2(new_n800), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n703), .B2(new_n1009), .ZN(new_n1026));
  INV_X1    g0826(.A(G159), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n790), .A2(new_n1027), .B1(new_n760), .B2(new_n343), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n316), .B1(new_n769), .B2(new_n203), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n762), .A2(new_n201), .B1(new_n765), .B2(new_n861), .ZN(new_n1030));
  NOR3_X1   g0830(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n284), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n754), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n852), .A2(G97), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n562), .A2(new_n564), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n793), .A2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .A4(new_n1036), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n783), .A2(new_n774), .B1(new_n777), .B2(new_n760), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n763), .A2(G317), .B1(new_n859), .B2(G303), .ZN(new_n1039));
  INV_X1    g0839(.A(G322), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1039), .B1(new_n1040), .B2(new_n790), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G311), .B2(new_n849), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1038), .B1(new_n1042), .B2(KEYINPUT48), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT107), .Z(new_n1044));
  OR2_X1    g0844(.A1(new_n1042), .A2(KEYINPUT48), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1044), .A2(KEYINPUT49), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n316), .B1(new_n766), .B2(G326), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1046), .B(new_n1047), .C1(new_n621), .C2(new_n775), .ZN(new_n1048));
  AOI21_X1  g0848(.A(KEYINPUT49), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1037), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1026), .B1(new_n1050), .B2(new_n750), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n747), .B2(new_n959), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1017), .A2(new_n1052), .ZN(G393));
  NAND2_X1  g0853(.A1(new_n803), .A2(new_n246), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n500), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n799), .B(new_n750), .C1(new_n709), .C2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n749), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n292), .B1(new_n765), .B2(new_n1040), .C1(new_n774), .C2(new_n760), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n852), .B2(G107), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT109), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n790), .A2(new_n755), .B1(new_n768), .B2(new_n762), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT52), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n849), .A2(G303), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n793), .A2(G116), .B1(G294), .B2(new_n859), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1060), .A2(new_n1062), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT110), .Z(new_n1066));
  AOI22_X1  g0866(.A1(G150), .A2(new_n772), .B1(new_n763), .B2(G159), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  XOR2_X1   g0868(.A(KEYINPUT108), .B(KEYINPUT51), .Z(new_n1069));
  AOI22_X1  g0869(.A1(new_n1068), .A2(new_n1069), .B1(new_n793), .B2(G77), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n760), .A2(new_n203), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n316), .B1(new_n769), .B2(new_n280), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(new_n766), .C2(new_n858), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1069), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n849), .A2(G50), .B1(new_n1067), .B2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1070), .A2(new_n853), .A3(new_n1073), .A4(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1066), .A2(new_n1076), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT111), .Z(new_n1078));
  OAI221_X1 g0878(.A(new_n1057), .B1(new_n1009), .B2(new_n971), .C1(new_n1078), .C2(new_n751), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n954), .A2(new_n747), .A3(new_n950), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n954), .A2(new_n950), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n1082), .A2(new_n1016), .A3(KEYINPUT112), .ZN(new_n1083));
  AOI21_X1  g0883(.A(KEYINPUT112), .B1(new_n1082), .B2(new_n1016), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n961), .A2(new_n710), .ZN(new_n1086));
  OAI21_X1  g0886(.A(KEYINPUT113), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1082), .A2(new_n1016), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT112), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1082), .A2(new_n1016), .A3(KEYINPUT112), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT113), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1092), .A2(new_n961), .A3(new_n1093), .A4(new_n710), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1081), .B1(new_n1087), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(G390));
  NAND2_X1  g0896(.A1(new_n467), .A2(new_n740), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n915), .A2(new_n684), .A3(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n740), .B1(new_n830), .B2(new_n831), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n912), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT116), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n926), .A2(new_n740), .A3(new_n919), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n827), .B1(new_n841), .B2(new_n719), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT114), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g0906(.A(KEYINPUT114), .B(new_n827), .C1(new_n841), .C2(new_n719), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1099), .A2(KEYINPUT116), .A3(new_n912), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1102), .A2(new_n1103), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n836), .A2(new_n827), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1103), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n926), .B1(new_n740), .B2(new_n919), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1098), .B1(new_n1110), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n905), .B(new_n902), .C1(new_n1108), .C2(new_n912), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1111), .A2(new_n926), .ZN(new_n1118));
  AOI21_X1  g0918(.A(KEYINPUT115), .B1(new_n1118), .B2(new_n902), .ZN(new_n1119));
  OAI211_X1 g0919(.A(KEYINPUT115), .B(new_n902), .C1(new_n904), .C2(new_n912), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n901), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1103), .B(new_n1117), .C1(new_n1119), .C2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n902), .B1(new_n904), .B2(new_n912), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT115), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1126), .A2(new_n901), .A3(new_n1120), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1103), .B1(new_n1127), .B2(new_n1117), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1116), .B1(new_n1123), .B2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1117), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n1112), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1131), .A2(new_n1115), .A3(new_n1122), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1129), .A2(new_n710), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1131), .A2(new_n747), .A3(new_n1122), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n901), .A2(new_n797), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n748), .B1(new_n1032), .B2(new_n844), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT117), .Z(new_n1137));
  INV_X1    g0937(.A(G125), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n762), .A2(new_n866), .B1(new_n765), .B2(new_n1138), .ZN(new_n1139));
  XOR2_X1   g0939(.A(KEYINPUT54), .B(G143), .Z(new_n1140));
  AOI211_X1 g0940(.A(new_n292), .B(new_n1139), .C1(new_n859), .C2(new_n1140), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n772), .A2(G128), .B1(new_n988), .B2(G50), .ZN(new_n1142));
  OAI21_X1  g0942(.A(KEYINPUT53), .B1(new_n760), .B2(new_n861), .ZN(new_n1143));
  OR3_X1    g0943(.A1(new_n760), .A2(KEYINPUT53), .A3(new_n861), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n1000), .A2(new_n862), .B1(new_n1027), .B2(new_n783), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n1000), .A2(new_n208), .B1(new_n343), .B2(new_n783), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n316), .B1(new_n763), .B2(G116), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n1055), .A2(new_n859), .B1(new_n766), .B2(G294), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n772), .A2(G283), .B1(new_n786), .B2(G87), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n865), .A2(new_n1148), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n1145), .A2(new_n1146), .B1(new_n1147), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1137), .B1(new_n1152), .B2(new_n750), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1135), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1133), .A2(new_n1134), .A3(new_n1154), .ZN(G378));
  XOR2_X1   g0955(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n683), .A2(new_n370), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n368), .A2(new_n887), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT55), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n383), .A2(new_n1160), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1157), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n383), .A2(new_n1160), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1165), .A2(new_n1156), .A3(new_n1166), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n797), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n748), .B1(G50), .B2(new_n844), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n316), .A2(G41), .ZN(new_n1171));
  AOI211_X1 g0971(.A(G50), .B(new_n1171), .C1(new_n434), .C2(new_n264), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1171), .B1(new_n774), .B2(new_n765), .C1(new_n208), .C2(new_n762), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n1035), .B2(new_n859), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n786), .A2(G77), .B1(new_n988), .B2(G58), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(G116), .A2(new_n772), .B1(new_n754), .B2(G97), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1174), .A2(new_n984), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT58), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1172), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  XOR2_X1   g0979(.A(KEYINPUT118), .B(G124), .Z(new_n1180));
  AOI211_X1 g0980(.A(G33), .B(G41), .C1(new_n766), .C2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n1027), .B2(new_n775), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT119), .ZN(new_n1183));
  INV_X1    g0983(.A(G128), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n762), .A2(new_n1184), .B1(new_n769), .B2(new_n862), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G132), .B2(new_n754), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n772), .A2(G125), .B1(new_n786), .B2(new_n1140), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(new_n861), .C2(new_n783), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1183), .A2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1179), .B1(new_n1178), .B2(new_n1177), .C1(new_n1190), .C2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1170), .B1(new_n1192), .B2(new_n750), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1169), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n922), .A2(G330), .A3(new_n927), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(new_n1168), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1198), .A2(new_n922), .A3(G330), .A4(new_n927), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n914), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT121), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  AND3_X1   g1003(.A1(new_n1197), .A2(new_n914), .A3(new_n1199), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n914), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1203), .B1(new_n1206), .B2(KEYINPUT121), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1195), .B1(new_n1207), .B2(new_n747), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1098), .B(KEYINPUT122), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1123), .A2(new_n1128), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1210), .B1(new_n1211), .B2(new_n1115), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1197), .A2(new_n914), .A3(new_n1199), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(KEYINPUT57), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n710), .B1(new_n1212), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1132), .A2(new_n1209), .ZN(new_n1218));
  AOI21_X1  g1018(.A(KEYINPUT57), .B1(new_n1207), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1208), .B1(new_n1217), .B2(new_n1219), .ZN(G375));
  NAND2_X1  g1020(.A1(new_n1110), .A2(new_n1114), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n747), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT123), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n912), .A2(new_n797), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n748), .B1(G68), .B2(new_n844), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n790), .A2(new_n866), .B1(new_n202), .B2(new_n775), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G159), .B2(new_n786), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n762), .A2(new_n862), .B1(new_n765), .B2(new_n1184), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n292), .B(new_n1228), .C1(G150), .C2(new_n859), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n849), .A2(new_n1140), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n793), .A2(G50), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1227), .A2(new_n1229), .A3(new_n1230), .A4(new_n1231), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n769), .A2(new_n208), .B1(new_n765), .B2(new_n611), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n316), .B(new_n1233), .C1(G283), .C2(new_n763), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n772), .A2(G294), .B1(new_n786), .B2(G97), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1234), .A2(new_n1036), .A3(new_n1235), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n1000), .A2(new_n621), .B1(new_n343), .B2(new_n776), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1232), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1225), .B1(new_n1238), .B2(new_n750), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1224), .A2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1222), .A2(new_n1223), .A3(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n746), .B1(new_n1110), .B2(new_n1114), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1240), .ZN(new_n1243));
  OAI21_X1  g1043(.A(KEYINPUT123), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1241), .A2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1110), .A2(new_n1114), .A3(new_n1098), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1116), .A2(new_n964), .A3(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1245), .A2(new_n1247), .ZN(G381));
  XNOR2_X1  g1048(.A(G375), .B(KEYINPUT124), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n838), .A2(new_n839), .B1(new_n842), .B2(new_n871), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(G393), .A2(G396), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1095), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  OR2_X1    g1052(.A1(new_n1252), .A2(G381), .ZN(new_n1253));
  OR4_X1    g1053(.A1(G387), .A2(new_n1249), .A3(G378), .A4(new_n1253), .ZN(G407));
  NAND2_X1  g1054(.A1(new_n690), .A2(G213), .ZN(new_n1255));
  OR3_X1    g1055(.A1(new_n1249), .A2(G378), .A3(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(G407), .A2(G213), .A3(new_n1256), .ZN(G409));
  INV_X1    g1057(.A(new_n1011), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1087), .A2(new_n1094), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n814), .B1(new_n1052), .B2(new_n1017), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1012), .B1(new_n1251), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1081), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1259), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1251), .A2(new_n1260), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(new_n1259), .B2(new_n1262), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1258), .B1(new_n1263), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1095), .A2(new_n1261), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1267), .B(new_n1011), .C1(new_n1095), .C2(new_n1264), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G378), .B(new_n1208), .C1(new_n1217), .C2(new_n1219), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1194), .B1(new_n1206), .B2(new_n746), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1213), .A2(KEYINPUT121), .A3(new_n1214), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1205), .A2(new_n1202), .ZN(new_n1273));
  AND3_X1   g1073(.A1(new_n1272), .A2(new_n964), .A3(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1271), .B1(new_n1274), .B2(new_n1218), .ZN(new_n1275));
  OAI21_X1  g1075(.A(KEYINPUT125), .B1(new_n1275), .B2(G378), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1195), .B1(new_n1215), .B2(new_n747), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1272), .A2(new_n964), .A3(new_n1273), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1277), .B1(new_n1212), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT125), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1134), .A2(new_n1154), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1131), .A2(new_n1122), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n711), .B1(new_n1282), .B2(new_n1116), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1281), .B1(new_n1283), .B2(new_n1132), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1279), .A2(new_n1280), .A3(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1270), .A2(new_n1276), .A3(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT62), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT60), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1246), .B1(new_n1115), .B2(new_n1288), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1110), .A2(new_n1098), .A3(KEYINPUT60), .A4(new_n1114), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1289), .A2(new_n710), .A3(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n1245), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n1250), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(G384), .A2(new_n1291), .A3(new_n1245), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1286), .A2(new_n1287), .A3(new_n1255), .A4(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT61), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1255), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1279), .A2(new_n1280), .A3(new_n1284), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1280), .B1(new_n1279), .B2(new_n1284), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1299), .B1(new_n1302), .B2(new_n1270), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1296), .A2(KEYINPUT126), .ZN(new_n1304));
  INV_X1    g1104(.A(G2897), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1255), .A2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT126), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1307), .B1(new_n1295), .B2(new_n1308), .ZN(new_n1309));
  AOI211_X1 g1109(.A(KEYINPUT126), .B(new_n1306), .C1(new_n1293), .C2(new_n1294), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1304), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1297), .B(new_n1298), .C1(new_n1303), .C2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1286), .A2(new_n1255), .A3(new_n1296), .ZN(new_n1313));
  AND2_X1   g1113(.A1(new_n1313), .A2(KEYINPUT62), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1269), .B1(new_n1312), .B2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1266), .A2(new_n1268), .A3(new_n1298), .ZN(new_n1316));
  XNOR2_X1  g1116(.A(new_n1316), .B(KEYINPUT127), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1286), .A2(new_n1255), .ZN(new_n1318));
  OAI211_X1 g1118(.A(new_n1318), .B(new_n1304), .C1(new_n1310), .C2(new_n1309), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1303), .A2(KEYINPUT63), .A3(new_n1296), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT63), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1313), .A2(new_n1321), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1317), .A2(new_n1319), .A3(new_n1320), .A4(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1315), .A2(new_n1323), .ZN(G405));
  XNOR2_X1  g1124(.A(G375), .B(G378), .ZN(new_n1325));
  XNOR2_X1  g1125(.A(new_n1325), .B(new_n1296), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1269), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  AND2_X1   g1128(.A1(new_n1325), .A2(new_n1295), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1325), .A2(new_n1295), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1269), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1328), .A2(new_n1331), .ZN(G402));
endmodule


