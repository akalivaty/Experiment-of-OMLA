

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733;

  NAND2_X1 U365 ( .A1(n541), .A2(n661), .ZN(n539) );
  XNOR2_X1 U366 ( .A(n611), .B(n610), .ZN(n612) );
  XNOR2_X2 U367 ( .A(n539), .B(n530), .ZN(n564) );
  XNOR2_X2 U368 ( .A(n550), .B(n437), .ZN(n647) );
  NOR2_X1 U369 ( .A1(n699), .A2(G902), .ZN(n502) );
  NOR2_X1 U370 ( .A1(n580), .A2(n344), .ZN(n401) );
  XNOR2_X1 U371 ( .A(n502), .B(n501), .ZN(n644) );
  XNOR2_X1 U372 ( .A(n445), .B(n444), .ZN(n484) );
  INV_X1 U373 ( .A(KEYINPUT64), .ZN(n386) );
  INV_X1 U374 ( .A(n612), .ZN(n343) );
  NOR2_X1 U375 ( .A1(n731), .A2(n349), .ZN(n593) );
  XNOR2_X1 U376 ( .A(n401), .B(KEYINPUT32), .ZN(n731) );
  XNOR2_X1 U377 ( .A(n387), .B(KEYINPUT67), .ZN(n648) );
  NOR2_X1 U378 ( .A1(n644), .A2(n643), .ZN(n387) );
  INV_X1 U379 ( .A(KEYINPUT72), .ZN(n391) );
  NOR2_X1 U380 ( .A1(n604), .A2(n603), .ZN(n607) );
  NOR2_X1 U381 ( .A1(n543), .A2(n425), .ZN(n424) );
  NOR2_X1 U382 ( .A1(n647), .A2(n648), .ZN(n589) );
  XNOR2_X1 U383 ( .A(n398), .B(KEYINPUT0), .ZN(n570) );
  XOR2_X1 U384 ( .A(KEYINPUT101), .B(n548), .Z(n632) );
  NOR2_X1 U385 ( .A1(n554), .A2(n517), .ZN(n548) );
  XNOR2_X1 U386 ( .A(n481), .B(G478), .ZN(n554) );
  OR2_X1 U387 ( .A1(n689), .A2(G902), .ZN(n438) );
  XNOR2_X1 U388 ( .A(n452), .B(n484), .ZN(n407) );
  XNOR2_X1 U389 ( .A(n605), .B(KEYINPUT45), .ZN(n606) );
  XNOR2_X1 U390 ( .A(n391), .B(G119), .ZN(n445) );
  XNOR2_X1 U391 ( .A(n373), .B(G134), .ZN(n478) );
  XNOR2_X1 U392 ( .A(G107), .B(KEYINPUT91), .ZN(n443) );
  XNOR2_X2 U393 ( .A(n446), .B(G113), .ZN(n465) );
  XNOR2_X2 U394 ( .A(G122), .B(G104), .ZN(n446) );
  XNOR2_X2 U395 ( .A(n441), .B(n439), .ZN(n541) );
  NOR2_X1 U396 ( .A1(n510), .A2(n416), .ZN(n415) );
  INV_X1 U397 ( .A(n544), .ZN(n416) );
  XNOR2_X1 U398 ( .A(n468), .B(n467), .ZN(n553) );
  BUF_X1 U399 ( .A(n644), .Z(n394) );
  AND2_X1 U400 ( .A1(n565), .A2(n678), .ZN(n399) );
  INV_X1 U401 ( .A(n609), .ZN(n610) );
  INV_X1 U402 ( .A(G902), .ZN(n479) );
  INV_X1 U403 ( .A(KEYINPUT75), .ZN(n372) );
  OR2_X1 U404 ( .A1(n733), .A2(n732), .ZN(n370) );
  XNOR2_X1 U405 ( .A(G113), .B(G101), .ZN(n483) );
  INV_X1 U406 ( .A(KEYINPUT76), .ZN(n427) );
  XNOR2_X1 U407 ( .A(n430), .B(n429), .ZN(n428) );
  XNOR2_X1 U408 ( .A(G137), .B(KEYINPUT5), .ZN(n429) );
  AND2_X1 U409 ( .A1(n482), .A2(G210), .ZN(n430) );
  XNOR2_X1 U410 ( .A(n478), .B(n454), .ZN(n719) );
  XNOR2_X1 U411 ( .A(KEYINPUT4), .B(G131), .ZN(n453) );
  XNOR2_X1 U412 ( .A(G140), .B(KEYINPUT68), .ZN(n450) );
  XOR2_X1 U413 ( .A(KEYINPUT78), .B(G104), .Z(n448) );
  XNOR2_X1 U414 ( .A(n719), .B(G146), .ZN(n486) );
  OR2_X1 U415 ( .A1(G902), .A2(G237), .ZN(n456) );
  XNOR2_X1 U416 ( .A(KEYINPUT15), .B(G902), .ZN(n609) );
  NOR2_X1 U417 ( .A1(n641), .A2(n421), .ZN(n420) );
  INV_X1 U418 ( .A(n639), .ZN(n421) );
  XNOR2_X1 U419 ( .A(n442), .B(n403), .ZN(n402) );
  XNOR2_X1 U420 ( .A(n463), .B(n345), .ZN(n442) );
  XNOR2_X1 U421 ( .A(n406), .B(n404), .ZN(n403) );
  XNOR2_X1 U422 ( .A(n436), .B(n590), .ZN(n671) );
  NAND2_X1 U423 ( .A1(n589), .A2(n588), .ZN(n436) );
  AND2_X1 U424 ( .A1(n632), .A2(n512), .ZN(n513) );
  NOR2_X1 U425 ( .A1(n511), .A2(n529), .ZN(n512) );
  NOR2_X1 U426 ( .A1(n671), .A2(n570), .ZN(n435) );
  INV_X1 U427 ( .A(KEYINPUT1), .ZN(n437) );
  XNOR2_X1 U428 ( .A(KEYINPUT66), .B(KEYINPUT22), .ZN(n568) );
  NOR2_X1 U429 ( .A1(n570), .A2(n643), .ZN(n567) );
  NAND2_X1 U430 ( .A1(n343), .A2(n363), .ZN(n434) );
  INV_X1 U431 ( .A(G478), .ZN(n364) );
  XNOR2_X1 U432 ( .A(n478), .B(n477), .ZN(n381) );
  NAND2_X1 U433 ( .A1(n343), .A2(n361), .ZN(n616) );
  INV_X1 U434 ( .A(G210), .ZN(n362) );
  NAND2_X1 U435 ( .A1(n383), .A2(n581), .ZN(n368) );
  XNOR2_X1 U436 ( .A(n540), .B(KEYINPUT36), .ZN(n383) );
  AND2_X1 U437 ( .A1(n538), .A2(n397), .ZN(n540) );
  INV_X1 U438 ( .A(n539), .ZN(n397) );
  INV_X1 U439 ( .A(KEYINPUT83), .ZN(n411) );
  XNOR2_X1 U440 ( .A(G125), .B(G146), .ZN(n464) );
  XNOR2_X1 U441 ( .A(n500), .B(n499), .ZN(n501) );
  NAND2_X1 U442 ( .A1(n371), .A2(n369), .ZN(n423) );
  XNOR2_X1 U443 ( .A(n370), .B(n413), .ZN(n369) );
  INV_X1 U444 ( .A(KEYINPUT46), .ZN(n413) );
  XOR2_X1 U445 ( .A(KEYINPUT98), .B(G140), .Z(n460) );
  XOR2_X1 U446 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n458) );
  INV_X1 U447 ( .A(n464), .ZN(n463) );
  NAND2_X1 U448 ( .A1(G237), .A2(G234), .ZN(n505) );
  XNOR2_X1 U449 ( .A(n428), .B(n426), .ZN(n485) );
  XNOR2_X1 U450 ( .A(n483), .B(n427), .ZN(n426) );
  XNOR2_X1 U451 ( .A(G128), .B(G110), .ZN(n489) );
  INV_X1 U452 ( .A(KEYINPUT8), .ZN(n469) );
  XNOR2_X1 U453 ( .A(n486), .B(n455), .ZN(n689) );
  XNOR2_X1 U454 ( .A(n451), .B(n396), .ZN(n455) );
  XNOR2_X1 U455 ( .A(n374), .B(n452), .ZN(n396) );
  XNOR2_X1 U456 ( .A(n547), .B(n385), .ZN(n560) );
  INV_X1 U457 ( .A(KEYINPUT39), .ZN(n385) );
  NOR2_X1 U458 ( .A1(n552), .A2(n546), .ZN(n547) );
  NAND2_X1 U459 ( .A1(n573), .A2(n678), .ZN(n543) );
  XNOR2_X1 U460 ( .A(n447), .B(n440), .ZN(n439) );
  INV_X1 U461 ( .A(KEYINPUT80), .ZN(n440) );
  NOR2_X1 U462 ( .A1(n418), .A2(n529), .ZN(n414) );
  INV_X1 U463 ( .A(KEYINPUT6), .ZN(n417) );
  NAND2_X1 U464 ( .A1(n343), .A2(n360), .ZN(n618) );
  BUF_X1 U465 ( .A(n725), .Z(n384) );
  NAND2_X1 U466 ( .A1(n343), .A2(n358), .ZN(n697) );
  INV_X1 U467 ( .A(G475), .ZN(n359) );
  XNOR2_X1 U468 ( .A(n549), .B(KEYINPUT40), .ZN(n733) );
  AND2_X1 U469 ( .A1(n560), .A2(n548), .ZN(n549) );
  XNOR2_X1 U470 ( .A(n435), .B(n352), .ZN(n395) );
  NAND2_X1 U471 ( .A1(n647), .A2(n418), .ZN(n400) );
  INV_X1 U472 ( .A(KEYINPUT120), .ZN(n431) );
  INV_X1 U473 ( .A(KEYINPUT56), .ZN(n379) );
  XNOR2_X1 U474 ( .A(n688), .B(n375), .ZN(G75) );
  XNOR2_X1 U475 ( .A(n376), .B(KEYINPUT115), .ZN(n375) );
  INV_X1 U476 ( .A(KEYINPUT53), .ZN(n376) );
  INV_X1 U477 ( .A(n368), .ZN(n637) );
  OR2_X1 U478 ( .A1(n350), .A2(n583), .ZN(n344) );
  INV_X1 U479 ( .A(G953), .ZN(n684) );
  XOR2_X1 U480 ( .A(KEYINPUT4), .B(KEYINPUT17), .Z(n345) );
  XOR2_X1 U481 ( .A(KEYINPUT16), .B(n465), .Z(n346) );
  XOR2_X1 U482 ( .A(G101), .B(G110), .Z(n347) );
  XNOR2_X1 U483 ( .A(n654), .B(n417), .ZN(n588) );
  OR2_X1 U484 ( .A1(n400), .A2(n583), .ZN(n348) );
  NOR2_X1 U485 ( .A1(n580), .A2(n348), .ZN(n349) );
  OR2_X1 U486 ( .A1(n588), .A2(n647), .ZN(n350) );
  OR2_X1 U487 ( .A1(n581), .A2(n588), .ZN(n351) );
  XOR2_X1 U488 ( .A(KEYINPUT79), .B(n587), .Z(n352) );
  XNOR2_X1 U489 ( .A(n505), .B(KEYINPUT14), .ZN(n678) );
  INV_X1 U490 ( .A(n703), .ZN(n388) );
  XOR2_X1 U491 ( .A(n617), .B(KEYINPUT62), .Z(n353) );
  XOR2_X1 U492 ( .A(n696), .B(n695), .Z(n354) );
  XNOR2_X1 U493 ( .A(n615), .B(n614), .ZN(n355) );
  XNOR2_X1 U494 ( .A(n381), .B(n476), .ZN(n480) );
  XNOR2_X1 U495 ( .A(KEYINPUT60), .B(KEYINPUT119), .ZN(n356) );
  XOR2_X1 U496 ( .A(KEYINPUT63), .B(KEYINPUT103), .Z(n357) );
  INV_X1 U497 ( .A(G472), .ZN(n419) );
  NOR2_X1 U498 ( .A1(n612), .A2(n642), .ZN(n365) );
  NOR2_X1 U499 ( .A1(n642), .A2(n359), .ZN(n358) );
  NOR2_X1 U500 ( .A1(n642), .A2(n419), .ZN(n360) );
  NOR2_X1 U501 ( .A1(n642), .A2(n362), .ZN(n361) );
  NOR2_X1 U502 ( .A1(n642), .A2(n364), .ZN(n363) );
  NAND2_X1 U503 ( .A1(n365), .A2(G469), .ZN(n692) );
  NAND2_X1 U504 ( .A1(n365), .A2(G217), .ZN(n701) );
  NAND2_X1 U505 ( .A1(n366), .A2(n368), .ZN(n367) );
  XNOR2_X1 U506 ( .A(n537), .B(n372), .ZN(n366) );
  XNOR2_X1 U507 ( .A(n367), .B(KEYINPUT71), .ZN(n371) );
  XNOR2_X1 U508 ( .A(n373), .B(n405), .ZN(n404) );
  XNOR2_X2 U509 ( .A(G143), .B(G128), .ZN(n373) );
  XNOR2_X2 U510 ( .A(n347), .B(n443), .ZN(n452) );
  XNOR2_X2 U511 ( .A(n569), .B(n568), .ZN(n580) );
  NAND2_X1 U512 ( .A1(n531), .A2(KEYINPUT47), .ZN(n412) );
  XNOR2_X1 U513 ( .A(n412), .B(n411), .ZN(n410) );
  XNOR2_X1 U514 ( .A(n414), .B(KEYINPUT28), .ZN(n551) );
  NOR2_X1 U515 ( .A1(n730), .A2(n599), .ZN(n598) );
  XNOR2_X1 U516 ( .A(n592), .B(KEYINPUT35), .ZN(n730) );
  NOR2_X1 U517 ( .A1(n580), .A2(n351), .ZN(n582) );
  XNOR2_X2 U518 ( .A(n608), .B(KEYINPUT2), .ZN(n642) );
  INV_X1 U519 ( .A(n496), .ZN(n374) );
  INV_X1 U520 ( .A(n570), .ZN(n572) );
  XNOR2_X2 U521 ( .A(n576), .B(KEYINPUT96), .ZN(n622) );
  NAND2_X1 U522 ( .A1(n433), .A2(n388), .ZN(n432) );
  XNOR2_X1 U523 ( .A(n434), .B(n480), .ZN(n433) );
  NOR2_X2 U524 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U525 ( .A(n423), .B(n559), .ZN(n422) );
  NAND2_X1 U526 ( .A1(n424), .A2(n522), .ZN(n629) );
  XNOR2_X1 U527 ( .A(n409), .B(KEYINPUT82), .ZN(n536) );
  XNOR2_X1 U528 ( .A(n377), .B(n357), .ZN(G57) );
  NAND2_X1 U529 ( .A1(n393), .A2(n388), .ZN(n377) );
  XNOR2_X1 U530 ( .A(n378), .B(n356), .ZN(G60) );
  NAND2_X1 U531 ( .A1(n392), .A2(n388), .ZN(n378) );
  XNOR2_X1 U532 ( .A(n380), .B(n379), .ZN(G51) );
  NAND2_X1 U533 ( .A1(n389), .A2(n388), .ZN(n380) );
  XNOR2_X1 U534 ( .A(n466), .B(n382), .ZN(n696) );
  XNOR2_X1 U535 ( .A(n495), .B(n465), .ZN(n382) );
  NAND2_X1 U536 ( .A1(n725), .A2(G234), .ZN(n470) );
  XNOR2_X2 U537 ( .A(n386), .B(G953), .ZN(n725) );
  XNOR2_X1 U538 ( .A(n616), .B(n355), .ZN(n389) );
  NOR2_X1 U539 ( .A1(n586), .A2(n390), .ZN(n597) );
  NAND2_X1 U540 ( .A1(n619), .A2(n585), .ZN(n390) );
  NOR2_X2 U541 ( .A1(n648), .A2(n518), .ZN(n573) );
  NAND2_X1 U542 ( .A1(n564), .A2(n399), .ZN(n398) );
  NAND2_X1 U543 ( .A1(n526), .A2(KEYINPUT81), .ZN(n527) );
  NAND2_X1 U544 ( .A1(n629), .A2(n523), .ZN(n526) );
  XNOR2_X1 U545 ( .A(n697), .B(n354), .ZN(n392) );
  XNOR2_X1 U546 ( .A(n618), .B(n353), .ZN(n393) );
  NOR2_X1 U547 ( .A1(n395), .A2(n591), .ZN(n592) );
  NAND2_X1 U548 ( .A1(n480), .A2(n479), .ZN(n481) );
  XNOR2_X2 U549 ( .A(n704), .B(n402), .ZN(n613) );
  XNOR2_X2 U550 ( .A(n346), .B(n407), .ZN(n704) );
  INV_X1 U551 ( .A(KEYINPUT18), .ZN(n405) );
  NAND2_X1 U552 ( .A1(n725), .A2(G224), .ZN(n406) );
  NAND2_X1 U553 ( .A1(n408), .A2(G221), .ZN(n494) );
  NAND2_X1 U554 ( .A1(n408), .A2(G217), .ZN(n477) );
  XNOR2_X2 U555 ( .A(n470), .B(n469), .ZN(n408) );
  NAND2_X1 U556 ( .A1(n532), .A2(n410), .ZN(n409) );
  NAND2_X1 U557 ( .A1(n394), .A2(n415), .ZN(n529) );
  INV_X1 U558 ( .A(n588), .ZN(n511) );
  NAND2_X1 U559 ( .A1(n521), .A2(n541), .ZN(n425) );
  NAND2_X1 U560 ( .A1(n613), .A2(n609), .ZN(n441) );
  NAND2_X1 U561 ( .A1(n572), .A2(n418), .ZN(n575) );
  INV_X1 U562 ( .A(n654), .ZN(n418) );
  XNOR2_X2 U563 ( .A(n488), .B(n419), .ZN(n654) );
  NAND2_X1 U564 ( .A1(n422), .A2(n420), .ZN(n724) );
  XNOR2_X1 U565 ( .A(n432), .B(n431), .ZN(G63) );
  XNOR2_X2 U566 ( .A(n438), .B(G469), .ZN(n550) );
  NOR2_X1 U567 ( .A1(n384), .A2(G952), .ZN(n703) );
  NOR2_X1 U568 ( .A1(n536), .A2(n535), .ZN(n537) );
  INV_X1 U569 ( .A(KEYINPUT48), .ZN(n558) );
  XNOR2_X1 U570 ( .A(n558), .B(KEYINPUT70), .ZN(n559) );
  XNOR2_X1 U571 ( .A(n449), .B(n448), .ZN(n451) );
  XNOR2_X1 U572 ( .A(n485), .B(n484), .ZN(n487) );
  XNOR2_X1 U573 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U574 ( .A(n486), .B(n487), .ZN(n617) );
  INV_X1 U575 ( .A(n542), .ZN(n522) );
  XNOR2_X1 U576 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X1 U577 ( .A(G116), .B(KEYINPUT3), .ZN(n444) );
  NAND2_X1 U578 ( .A1(G210), .A2(n456), .ZN(n447) );
  NAND2_X1 U579 ( .A1(G227), .A2(n725), .ZN(n449) );
  XNOR2_X1 U580 ( .A(n450), .B(G137), .ZN(n496) );
  XNOR2_X1 U581 ( .A(n453), .B(KEYINPUT69), .ZN(n454) );
  INV_X1 U582 ( .A(n647), .ZN(n581) );
  NAND2_X1 U583 ( .A1(G214), .A2(n456), .ZN(n661) );
  XNOR2_X1 U584 ( .A(KEYINPUT13), .B(G475), .ZN(n468) );
  NOR2_X1 U585 ( .A1(G953), .A2(G237), .ZN(n482) );
  NAND2_X1 U586 ( .A1(n482), .A2(G214), .ZN(n457) );
  XNOR2_X1 U587 ( .A(n458), .B(n457), .ZN(n462) );
  XNOR2_X1 U588 ( .A(G143), .B(G131), .ZN(n459) );
  XNOR2_X1 U589 ( .A(n460), .B(n459), .ZN(n461) );
  XOR2_X1 U590 ( .A(n462), .B(n461), .Z(n466) );
  XNOR2_X1 U591 ( .A(KEYINPUT10), .B(n464), .ZN(n495) );
  NOR2_X1 U592 ( .A1(G902), .A2(n696), .ZN(n467) );
  INV_X1 U593 ( .A(n553), .ZN(n517) );
  XNOR2_X1 U594 ( .A(G122), .B(G107), .ZN(n471) );
  XNOR2_X1 U595 ( .A(n471), .B(KEYINPUT99), .ZN(n475) );
  XOR2_X1 U596 ( .A(KEYINPUT9), .B(KEYINPUT100), .Z(n473) );
  XNOR2_X1 U597 ( .A(G116), .B(KEYINPUT7), .ZN(n472) );
  XNOR2_X1 U598 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U599 ( .A(n474), .B(n475), .Z(n476) );
  NOR2_X1 U600 ( .A1(n617), .A2(G902), .ZN(n488) );
  XOR2_X1 U601 ( .A(KEYINPUT23), .B(G119), .Z(n490) );
  XNOR2_X1 U602 ( .A(n490), .B(n489), .ZN(n492) );
  XOR2_X1 U603 ( .A(KEYINPUT24), .B(KEYINPUT94), .Z(n491) );
  XNOR2_X1 U604 ( .A(n494), .B(n493), .ZN(n497) );
  XNOR2_X1 U605 ( .A(n496), .B(n495), .ZN(n718) );
  XNOR2_X1 U606 ( .A(n497), .B(n718), .ZN(n699) );
  NAND2_X1 U607 ( .A1(n609), .A2(G234), .ZN(n498) );
  XNOR2_X1 U608 ( .A(n498), .B(KEYINPUT20), .ZN(n506) );
  NAND2_X1 U609 ( .A1(G217), .A2(n506), .ZN(n500) );
  INV_X1 U610 ( .A(KEYINPUT25), .ZN(n499) );
  NOR2_X1 U611 ( .A1(n384), .A2(G900), .ZN(n503) );
  NAND2_X1 U612 ( .A1(G902), .A2(n503), .ZN(n504) );
  NAND2_X1 U613 ( .A1(G952), .A2(n684), .ZN(n562) );
  NAND2_X1 U614 ( .A1(n504), .A2(n562), .ZN(n544) );
  INV_X1 U615 ( .A(n678), .ZN(n509) );
  XOR2_X1 U616 ( .A(KEYINPUT95), .B(KEYINPUT21), .Z(n508) );
  NAND2_X1 U617 ( .A1(G221), .A2(n506), .ZN(n507) );
  XNOR2_X1 U618 ( .A(n508), .B(n507), .ZN(n643) );
  OR2_X1 U619 ( .A1(n509), .A2(n643), .ZN(n510) );
  XNOR2_X1 U620 ( .A(n513), .B(KEYINPUT102), .ZN(n538) );
  NAND2_X1 U621 ( .A1(n661), .A2(n538), .ZN(n514) );
  NOR2_X1 U622 ( .A1(n581), .A2(n514), .ZN(n515) );
  XNOR2_X1 U623 ( .A(n515), .B(KEYINPUT43), .ZN(n516) );
  NOR2_X1 U624 ( .A1(n541), .A2(n516), .ZN(n641) );
  AND2_X1 U625 ( .A1(n554), .A2(n517), .ZN(n634) );
  NOR2_X1 U626 ( .A1(n548), .A2(n634), .ZN(n667) );
  NAND2_X1 U627 ( .A1(KEYINPUT47), .A2(n667), .ZN(n523) );
  INV_X1 U628 ( .A(n550), .ZN(n518) );
  NAND2_X1 U629 ( .A1(n654), .A2(n661), .ZN(n519) );
  XNOR2_X1 U630 ( .A(KEYINPUT30), .B(n519), .ZN(n542) );
  NAND2_X1 U631 ( .A1(n554), .A2(n553), .ZN(n591) );
  INV_X1 U632 ( .A(n591), .ZN(n520) );
  AND2_X1 U633 ( .A1(n520), .A2(n544), .ZN(n521) );
  INV_X1 U634 ( .A(n526), .ZN(n525) );
  INV_X1 U635 ( .A(KEYINPUT81), .ZN(n524) );
  NAND2_X1 U636 ( .A1(n525), .A2(n524), .ZN(n528) );
  NAND2_X1 U637 ( .A1(n528), .A2(n527), .ZN(n532) );
  XOR2_X1 U638 ( .A(KEYINPUT77), .B(KEYINPUT19), .Z(n530) );
  AND2_X1 U639 ( .A1(n550), .A2(n564), .ZN(n533) );
  NAND2_X1 U640 ( .A1(n551), .A2(n533), .ZN(n531) );
  AND2_X1 U641 ( .A1(n551), .A2(n533), .ZN(n630) );
  XOR2_X1 U642 ( .A(KEYINPUT84), .B(n667), .Z(n578) );
  NAND2_X1 U643 ( .A1(n630), .A2(n578), .ZN(n534) );
  NOR2_X1 U644 ( .A1(n534), .A2(KEYINPUT47), .ZN(n535) );
  XNOR2_X1 U645 ( .A(KEYINPUT38), .B(n541), .ZN(n552) );
  NOR2_X1 U646 ( .A1(n543), .A2(n542), .ZN(n545) );
  NAND2_X1 U647 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U648 ( .A1(n551), .A2(n550), .ZN(n556) );
  INV_X1 U649 ( .A(n552), .ZN(n662) );
  NAND2_X1 U650 ( .A1(n662), .A2(n661), .ZN(n666) );
  NOR2_X1 U651 ( .A1(n554), .A2(n553), .ZN(n566) );
  INV_X1 U652 ( .A(n566), .ZN(n665) );
  NOR2_X1 U653 ( .A1(n666), .A2(n665), .ZN(n555) );
  XNOR2_X1 U654 ( .A(KEYINPUT41), .B(n555), .ZN(n660) );
  NOR2_X1 U655 ( .A1(n556), .A2(n660), .ZN(n557) );
  XNOR2_X1 U656 ( .A(n557), .B(KEYINPUT42), .ZN(n732) );
  NAND2_X1 U657 ( .A1(n560), .A2(n634), .ZN(n639) );
  INV_X1 U658 ( .A(n394), .ZN(n583) );
  XOR2_X1 U659 ( .A(KEYINPUT92), .B(G898), .Z(n711) );
  NAND2_X1 U660 ( .A1(n711), .A2(G953), .ZN(n561) );
  XNOR2_X1 U661 ( .A(n561), .B(KEYINPUT93), .ZN(n706) );
  NAND2_X1 U662 ( .A1(n706), .A2(G902), .ZN(n563) );
  NAND2_X1 U663 ( .A1(n563), .A2(n562), .ZN(n565) );
  NAND2_X1 U664 ( .A1(n567), .A2(n566), .ZN(n569) );
  NOR2_X1 U665 ( .A1(KEYINPUT73), .A2(KEYINPUT44), .ZN(n594) );
  NOR2_X1 U666 ( .A1(n593), .A2(n594), .ZN(n586) );
  AND2_X1 U667 ( .A1(n654), .A2(n589), .ZN(n657) );
  NAND2_X1 U668 ( .A1(n572), .A2(n657), .ZN(n571) );
  XNOR2_X1 U669 ( .A(n571), .B(KEYINPUT31), .ZN(n635) );
  INV_X1 U670 ( .A(n573), .ZN(n574) );
  NOR2_X1 U671 ( .A1(n635), .A2(n622), .ZN(n577) );
  XNOR2_X1 U672 ( .A(n577), .B(KEYINPUT97), .ZN(n579) );
  NAND2_X1 U673 ( .A1(n579), .A2(n578), .ZN(n585) );
  XNOR2_X1 U674 ( .A(n582), .B(KEYINPUT88), .ZN(n584) );
  NAND2_X1 U675 ( .A1(n584), .A2(n583), .ZN(n619) );
  XOR2_X1 U676 ( .A(KEYINPUT74), .B(KEYINPUT34), .Z(n587) );
  XOR2_X1 U677 ( .A(KEYINPUT90), .B(KEYINPUT33), .Z(n590) );
  AND2_X1 U678 ( .A1(n730), .A2(n593), .ZN(n595) );
  NAND2_X1 U679 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U680 ( .A1(n597), .A2(n596), .ZN(n604) );
  INV_X1 U681 ( .A(KEYINPUT44), .ZN(n599) );
  XNOR2_X1 U682 ( .A(n598), .B(KEYINPUT89), .ZN(n602) );
  NAND2_X1 U683 ( .A1(n599), .A2(n730), .ZN(n600) );
  NAND2_X1 U684 ( .A1(n600), .A2(KEYINPUT73), .ZN(n601) );
  NAND2_X1 U685 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U686 ( .A(KEYINPUT65), .B(KEYINPUT87), .ZN(n605) );
  XNOR2_X1 U687 ( .A(n607), .B(n606), .ZN(n707) );
  NOR2_X2 U688 ( .A1(n724), .A2(n707), .ZN(n608) );
  NOR2_X2 U689 ( .A1(n608), .A2(KEYINPUT86), .ZN(n611) );
  XOR2_X1 U690 ( .A(KEYINPUT55), .B(KEYINPUT54), .Z(n615) );
  XNOR2_X1 U691 ( .A(n613), .B(KEYINPUT116), .ZN(n614) );
  XNOR2_X1 U692 ( .A(n619), .B(G101), .ZN(G3) );
  NAND2_X1 U693 ( .A1(n622), .A2(n632), .ZN(n620) );
  XNOR2_X1 U694 ( .A(n620), .B(KEYINPUT104), .ZN(n621) );
  XNOR2_X1 U695 ( .A(G104), .B(n621), .ZN(G6) );
  XOR2_X1 U696 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n624) );
  NAND2_X1 U697 ( .A1(n634), .A2(n622), .ZN(n623) );
  XNOR2_X1 U698 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U699 ( .A(G107), .B(n625), .ZN(G9) );
  XOR2_X1 U700 ( .A(G110), .B(n349), .Z(G12) );
  XOR2_X1 U701 ( .A(KEYINPUT105), .B(KEYINPUT29), .Z(n627) );
  NAND2_X1 U702 ( .A1(n634), .A2(n630), .ZN(n626) );
  XNOR2_X1 U703 ( .A(n627), .B(n626), .ZN(n628) );
  XOR2_X1 U704 ( .A(G128), .B(n628), .Z(G30) );
  XNOR2_X1 U705 ( .A(n629), .B(G143), .ZN(G45) );
  NAND2_X1 U706 ( .A1(n630), .A2(n632), .ZN(n631) );
  XNOR2_X1 U707 ( .A(n631), .B(G146), .ZN(G48) );
  NAND2_X1 U708 ( .A1(n635), .A2(n632), .ZN(n633) );
  XNOR2_X1 U709 ( .A(n633), .B(G113), .ZN(G15) );
  NAND2_X1 U710 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U711 ( .A(n636), .B(G116), .ZN(G18) );
  XNOR2_X1 U712 ( .A(n637), .B(G125), .ZN(n638) );
  XNOR2_X1 U713 ( .A(n638), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U714 ( .A(G134), .B(KEYINPUT106), .ZN(n640) );
  XNOR2_X1 U715 ( .A(n640), .B(n639), .ZN(G36) );
  XOR2_X1 U716 ( .A(G140), .B(n641), .Z(G42) );
  XNOR2_X1 U717 ( .A(n642), .B(KEYINPUT85), .ZN(n687) );
  NOR2_X1 U718 ( .A1(n671), .A2(n660), .ZN(n682) );
  NAND2_X1 U719 ( .A1(n394), .A2(n643), .ZN(n645) );
  XNOR2_X1 U720 ( .A(n645), .B(KEYINPUT107), .ZN(n646) );
  XNOR2_X1 U721 ( .A(KEYINPUT49), .B(n646), .ZN(n652) );
  NAND2_X1 U722 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U723 ( .A(n649), .B(KEYINPUT50), .ZN(n650) );
  XNOR2_X1 U724 ( .A(KEYINPUT108), .B(n650), .ZN(n651) );
  NAND2_X1 U725 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U726 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U727 ( .A(KEYINPUT109), .B(n655), .Z(n656) );
  NOR2_X1 U728 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U729 ( .A(KEYINPUT51), .B(n658), .Z(n659) );
  NOR2_X1 U730 ( .A1(n660), .A2(n659), .ZN(n674) );
  NOR2_X1 U731 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U732 ( .A(n663), .B(KEYINPUT110), .ZN(n664) );
  NOR2_X1 U733 ( .A1(n665), .A2(n664), .ZN(n669) );
  NOR2_X1 U734 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U735 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U736 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U737 ( .A(KEYINPUT111), .B(n672), .Z(n673) );
  NOR2_X1 U738 ( .A1(n674), .A2(n673), .ZN(n677) );
  XOR2_X1 U739 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n675) );
  XNOR2_X1 U740 ( .A(KEYINPUT52), .B(n675), .ZN(n676) );
  XNOR2_X1 U741 ( .A(n677), .B(n676), .ZN(n680) );
  NAND2_X1 U742 ( .A1(n678), .A2(G952), .ZN(n679) );
  NOR2_X1 U743 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U744 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U745 ( .A(n683), .B(KEYINPUT114), .ZN(n685) );
  NAND2_X1 U746 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U747 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U748 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n691) );
  XNOR2_X1 U749 ( .A(n689), .B(KEYINPUT117), .ZN(n690) );
  XNOR2_X1 U750 ( .A(n691), .B(n690), .ZN(n693) );
  XOR2_X1 U751 ( .A(n693), .B(n692), .Z(n694) );
  NOR2_X1 U752 ( .A1(n703), .A2(n694), .ZN(G54) );
  XOR2_X1 U753 ( .A(KEYINPUT118), .B(KEYINPUT59), .Z(n695) );
  INV_X1 U754 ( .A(KEYINPUT121), .ZN(n698) );
  XNOR2_X1 U755 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U756 ( .A1(n703), .A2(n702), .ZN(G66) );
  XNOR2_X1 U757 ( .A(KEYINPUT124), .B(n704), .ZN(n705) );
  NOR2_X1 U758 ( .A1(n706), .A2(n705), .ZN(n716) );
  NOR2_X1 U759 ( .A1(G953), .A2(n707), .ZN(n714) );
  XOR2_X1 U760 ( .A(KEYINPUT122), .B(KEYINPUT61), .Z(n709) );
  NAND2_X1 U761 ( .A1(G224), .A2(G953), .ZN(n708) );
  XNOR2_X1 U762 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X1 U763 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U764 ( .A(KEYINPUT123), .B(n712), .Z(n713) );
  NOR2_X1 U765 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U766 ( .A(n716), .B(n715), .Z(n717) );
  XOR2_X1 U767 ( .A(KEYINPUT125), .B(n717), .Z(G69) );
  XNOR2_X1 U768 ( .A(n719), .B(n718), .ZN(n723) );
  XNOR2_X1 U769 ( .A(G227), .B(n723), .ZN(n720) );
  NAND2_X1 U770 ( .A1(n720), .A2(G900), .ZN(n721) );
  XNOR2_X1 U771 ( .A(n721), .B(KEYINPUT126), .ZN(n722) );
  NAND2_X1 U772 ( .A1(n722), .A2(G953), .ZN(n728) );
  XNOR2_X1 U773 ( .A(n724), .B(n723), .ZN(n726) );
  NAND2_X1 U774 ( .A1(n726), .A2(n384), .ZN(n727) );
  NAND2_X1 U775 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U776 ( .A(KEYINPUT127), .B(n729), .Z(G72) );
  XNOR2_X1 U777 ( .A(n730), .B(G122), .ZN(G24) );
  XOR2_X1 U778 ( .A(G119), .B(n731), .Z(G21) );
  XOR2_X1 U779 ( .A(G137), .B(n732), .Z(G39) );
  XOR2_X1 U780 ( .A(G131), .B(n733), .Z(G33) );
endmodule

