

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572;

  XOR2_X1 U319 ( .A(n386), .B(n385), .Z(n287) );
  XNOR2_X1 U320 ( .A(KEYINPUT118), .B(KEYINPUT54), .ZN(n434) );
  XNOR2_X1 U321 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U322 ( .A(n387), .B(n287), .ZN(n388) );
  XNOR2_X1 U323 ( .A(n389), .B(n388), .ZN(n561) );
  NOR2_X1 U324 ( .A1(n515), .A2(n438), .ZN(n551) );
  XNOR2_X1 U325 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n439) );
  XNOR2_X1 U326 ( .A(n440), .B(n439), .ZN(G1351GAT) );
  XOR2_X1 U327 ( .A(KEYINPUT78), .B(G176GAT), .Z(n289) );
  XNOR2_X1 U328 ( .A(G169GAT), .B(G120GAT), .ZN(n288) );
  XNOR2_X1 U329 ( .A(n289), .B(n288), .ZN(n293) );
  XOR2_X1 U330 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n291) );
  XNOR2_X1 U331 ( .A(G113GAT), .B(KEYINPUT20), .ZN(n290) );
  XNOR2_X1 U332 ( .A(n291), .B(n290), .ZN(n292) );
  XNOR2_X1 U333 ( .A(n293), .B(n292), .ZN(n305) );
  XOR2_X1 U334 ( .A(KEYINPUT0), .B(G127GAT), .Z(n336) );
  XOR2_X1 U335 ( .A(G190GAT), .B(G134GAT), .Z(n295) );
  XNOR2_X1 U336 ( .A(G43GAT), .B(G99GAT), .ZN(n294) );
  XNOR2_X1 U337 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U338 ( .A(n336), .B(n296), .Z(n298) );
  NAND2_X1 U339 ( .A1(G227GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U340 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U341 ( .A(n299), .B(G71GAT), .Z(n303) );
  XOR2_X1 U342 ( .A(G183GAT), .B(KEYINPUT17), .Z(n301) );
  XNOR2_X1 U343 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n300) );
  XNOR2_X1 U344 ( .A(n301), .B(n300), .ZN(n429) );
  XNOR2_X1 U345 ( .A(G15GAT), .B(n429), .ZN(n302) );
  XNOR2_X1 U346 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U347 ( .A(n305), .B(n304), .ZN(n515) );
  XOR2_X1 U348 ( .A(G148GAT), .B(KEYINPUT22), .Z(n311) );
  XOR2_X1 U349 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n307) );
  XNOR2_X1 U350 ( .A(G22GAT), .B(KEYINPUT82), .ZN(n306) );
  XNOR2_X1 U351 ( .A(n307), .B(n306), .ZN(n309) );
  XNOR2_X1 U352 ( .A(G106GAT), .B(G78GAT), .ZN(n308) );
  XNOR2_X1 U353 ( .A(n308), .B(G204GAT), .ZN(n384) );
  XNOR2_X1 U354 ( .A(n309), .B(n384), .ZN(n310) );
  XNOR2_X1 U355 ( .A(n311), .B(n310), .ZN(n317) );
  XOR2_X1 U356 ( .A(G211GAT), .B(KEYINPUT21), .Z(n313) );
  XNOR2_X1 U357 ( .A(G197GAT), .B(G218GAT), .ZN(n312) );
  XNOR2_X1 U358 ( .A(n313), .B(n312), .ZN(n421) );
  XOR2_X1 U359 ( .A(n421), .B(KEYINPUT81), .Z(n315) );
  NAND2_X1 U360 ( .A1(G228GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U361 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U362 ( .A(n317), .B(n316), .Z(n324) );
  XOR2_X1 U363 ( .A(KEYINPUT3), .B(KEYINPUT84), .Z(n319) );
  XNOR2_X1 U364 ( .A(G162GAT), .B(KEYINPUT2), .ZN(n318) );
  XNOR2_X1 U365 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U366 ( .A(n320), .B(KEYINPUT83), .Z(n322) );
  XNOR2_X1 U367 ( .A(G141GAT), .B(G155GAT), .ZN(n321) );
  XNOR2_X1 U368 ( .A(n322), .B(n321), .ZN(n328) );
  XNOR2_X1 U369 ( .A(G50GAT), .B(n328), .ZN(n323) );
  XNOR2_X1 U370 ( .A(n324), .B(n323), .ZN(n450) );
  XOR2_X1 U371 ( .A(KEYINPUT4), .B(KEYINPUT87), .Z(n326) );
  XNOR2_X1 U372 ( .A(KEYINPUT5), .B(KEYINPUT85), .ZN(n325) );
  XNOR2_X1 U373 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U374 ( .A(n328), .B(n327), .ZN(n340) );
  XOR2_X1 U375 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n330) );
  XNOR2_X1 U376 ( .A(G85GAT), .B(KEYINPUT86), .ZN(n329) );
  XNOR2_X1 U377 ( .A(n330), .B(n329), .ZN(n335) );
  XNOR2_X1 U378 ( .A(G120GAT), .B(G148GAT), .ZN(n331) );
  XNOR2_X1 U379 ( .A(n331), .B(G57GAT), .ZN(n380) );
  XOR2_X1 U380 ( .A(G29GAT), .B(G134GAT), .Z(n353) );
  XOR2_X1 U381 ( .A(n380), .B(n353), .Z(n333) );
  NAND2_X1 U382 ( .A1(G225GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U383 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U384 ( .A(n335), .B(n334), .Z(n338) );
  XOR2_X1 U385 ( .A(G113GAT), .B(G1GAT), .Z(n360) );
  XNOR2_X1 U386 ( .A(n360), .B(n336), .ZN(n337) );
  XNOR2_X1 U387 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U388 ( .A(n340), .B(n339), .ZN(n449) );
  XNOR2_X1 U389 ( .A(KEYINPUT88), .B(n449), .ZN(n499) );
  XOR2_X1 U390 ( .A(KEYINPUT11), .B(KEYINPUT76), .Z(n342) );
  XNOR2_X1 U391 ( .A(G218GAT), .B(KEYINPUT9), .ZN(n341) );
  XNOR2_X1 U392 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U393 ( .A(KEYINPUT65), .B(KEYINPUT10), .Z(n344) );
  XNOR2_X1 U394 ( .A(G162GAT), .B(G106GAT), .ZN(n343) );
  XNOR2_X1 U395 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U396 ( .A(n346), .B(n345), .ZN(n357) );
  XNOR2_X1 U397 ( .A(G99GAT), .B(G85GAT), .ZN(n347) );
  XNOR2_X1 U398 ( .A(n347), .B(KEYINPUT72), .ZN(n383) );
  XOR2_X1 U399 ( .A(G92GAT), .B(n383), .Z(n349) );
  NAND2_X1 U400 ( .A1(G232GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U401 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U402 ( .A(G36GAT), .B(G190GAT), .Z(n419) );
  XOR2_X1 U403 ( .A(n350), .B(n419), .Z(n355) );
  XOR2_X1 U404 ( .A(G43GAT), .B(G50GAT), .Z(n352) );
  XNOR2_X1 U405 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n351) );
  XNOR2_X1 U406 ( .A(n352), .B(n351), .ZN(n371) );
  XNOR2_X1 U407 ( .A(n371), .B(n353), .ZN(n354) );
  XNOR2_X1 U408 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U409 ( .A(n357), .B(n356), .ZN(n538) );
  XOR2_X1 U410 ( .A(G169GAT), .B(G8GAT), .Z(n420) );
  XOR2_X1 U411 ( .A(G22GAT), .B(G15GAT), .Z(n394) );
  XOR2_X1 U412 ( .A(n420), .B(n394), .Z(n359) );
  NAND2_X1 U413 ( .A1(G229GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U414 ( .A(n359), .B(n358), .ZN(n361) );
  XOR2_X1 U415 ( .A(n361), .B(n360), .Z(n369) );
  XOR2_X1 U416 ( .A(G197GAT), .B(G141GAT), .Z(n363) );
  XNOR2_X1 U417 ( .A(G29GAT), .B(G36GAT), .ZN(n362) );
  XNOR2_X1 U418 ( .A(n363), .B(n362), .ZN(n367) );
  XOR2_X1 U419 ( .A(KEYINPUT66), .B(KEYINPUT67), .Z(n365) );
  XNOR2_X1 U420 ( .A(KEYINPUT69), .B(KEYINPUT29), .ZN(n364) );
  XNOR2_X1 U421 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U422 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U423 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U424 ( .A(n370), .B(KEYINPUT68), .Z(n373) );
  XNOR2_X1 U425 ( .A(n371), .B(KEYINPUT30), .ZN(n372) );
  XNOR2_X1 U426 ( .A(n373), .B(n372), .ZN(n556) );
  XOR2_X1 U427 ( .A(KEYINPUT73), .B(KEYINPUT75), .Z(n375) );
  NAND2_X1 U428 ( .A1(G230GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U429 ( .A(n375), .B(n374), .ZN(n378) );
  XOR2_X1 U430 ( .A(KEYINPUT71), .B(KEYINPUT13), .Z(n377) );
  XNOR2_X1 U431 ( .A(G71GAT), .B(KEYINPUT70), .ZN(n376) );
  XNOR2_X1 U432 ( .A(n377), .B(n376), .ZN(n393) );
  XOR2_X1 U433 ( .A(n378), .B(n393), .Z(n382) );
  XNOR2_X1 U434 ( .A(G176GAT), .B(G92GAT), .ZN(n379) );
  XNOR2_X1 U435 ( .A(n379), .B(G64GAT), .ZN(n428) );
  XNOR2_X1 U436 ( .A(n380), .B(n428), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n382), .B(n381), .ZN(n389) );
  XNOR2_X1 U438 ( .A(n384), .B(n383), .ZN(n387) );
  XOR2_X1 U439 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n386) );
  XNOR2_X1 U440 ( .A(KEYINPUT32), .B(KEYINPUT74), .ZN(n385) );
  XOR2_X1 U441 ( .A(n561), .B(KEYINPUT41), .Z(n548) );
  NAND2_X1 U442 ( .A1(n556), .A2(n548), .ZN(n390) );
  XNOR2_X1 U443 ( .A(KEYINPUT46), .B(n390), .ZN(n408) );
  XOR2_X1 U444 ( .A(G57GAT), .B(G211GAT), .Z(n392) );
  XNOR2_X1 U445 ( .A(G183GAT), .B(G127GAT), .ZN(n391) );
  XNOR2_X1 U446 ( .A(n392), .B(n391), .ZN(n407) );
  XOR2_X1 U447 ( .A(n393), .B(G78GAT), .Z(n396) );
  XNOR2_X1 U448 ( .A(n394), .B(G155GAT), .ZN(n395) );
  XNOR2_X1 U449 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U450 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n398) );
  NAND2_X1 U451 ( .A1(G231GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U452 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U453 ( .A(n400), .B(n399), .Z(n405) );
  XOR2_X1 U454 ( .A(KEYINPUT77), .B(G64GAT), .Z(n402) );
  XNOR2_X1 U455 ( .A(G1GAT), .B(G8GAT), .ZN(n401) );
  XNOR2_X1 U456 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U457 ( .A(n403), .B(KEYINPUT14), .ZN(n404) );
  XNOR2_X1 U458 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U459 ( .A(n407), .B(n406), .Z(n456) );
  NAND2_X1 U460 ( .A1(n408), .A2(n456), .ZN(n409) );
  NOR2_X1 U461 ( .A1(n538), .A2(n409), .ZN(n411) );
  XNOR2_X1 U462 ( .A(KEYINPUT47), .B(KEYINPUT110), .ZN(n410) );
  XNOR2_X1 U463 ( .A(n411), .B(n410), .ZN(n417) );
  XOR2_X1 U464 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n413) );
  INV_X1 U465 ( .A(n456), .ZN(n564) );
  XNOR2_X1 U466 ( .A(KEYINPUT36), .B(n538), .ZN(n567) );
  NAND2_X1 U467 ( .A1(n564), .A2(n567), .ZN(n412) );
  XNOR2_X1 U468 ( .A(n413), .B(n412), .ZN(n415) );
  NOR2_X1 U469 ( .A1(n556), .A2(n561), .ZN(n414) );
  NAND2_X1 U470 ( .A1(n415), .A2(n414), .ZN(n416) );
  NAND2_X1 U471 ( .A1(n417), .A2(n416), .ZN(n418) );
  XNOR2_X1 U472 ( .A(KEYINPUT48), .B(n418), .ZN(n528) );
  XNOR2_X1 U473 ( .A(n420), .B(n419), .ZN(n433) );
  XOR2_X1 U474 ( .A(n421), .B(KEYINPUT77), .Z(n423) );
  NAND2_X1 U475 ( .A1(G226GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U476 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U477 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n425) );
  XNOR2_X1 U478 ( .A(G204GAT), .B(KEYINPUT91), .ZN(n424) );
  XNOR2_X1 U479 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U480 ( .A(n427), .B(n426), .Z(n431) );
  XNOR2_X1 U481 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U482 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U483 ( .A(n433), .B(n432), .ZN(n502) );
  NAND2_X1 U484 ( .A1(n528), .A2(n502), .ZN(n435) );
  NOR2_X1 U485 ( .A1(n499), .A2(n436), .ZN(n554) );
  NAND2_X1 U486 ( .A1(n450), .A2(n554), .ZN(n437) );
  XOR2_X1 U487 ( .A(KEYINPUT55), .B(n437), .Z(n438) );
  NAND2_X1 U488 ( .A1(n551), .A2(n538), .ZN(n440) );
  XNOR2_X1 U489 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n461) );
  INV_X1 U490 ( .A(n515), .ZN(n505) );
  NAND2_X1 U491 ( .A1(n502), .A2(n505), .ZN(n441) );
  NAND2_X1 U492 ( .A1(n450), .A2(n441), .ZN(n442) );
  XNOR2_X1 U493 ( .A(KEYINPUT25), .B(n442), .ZN(n447) );
  NOR2_X1 U494 ( .A1(n450), .A2(n505), .ZN(n444) );
  XNOR2_X1 U495 ( .A(KEYINPUT94), .B(KEYINPUT26), .ZN(n443) );
  XNOR2_X1 U496 ( .A(n444), .B(n443), .ZN(n553) );
  XNOR2_X1 U497 ( .A(n502), .B(KEYINPUT27), .ZN(n451) );
  NAND2_X1 U498 ( .A1(n553), .A2(n451), .ZN(n445) );
  XNOR2_X1 U499 ( .A(KEYINPUT95), .B(n445), .ZN(n446) );
  NOR2_X1 U500 ( .A1(n447), .A2(n446), .ZN(n448) );
  NOR2_X1 U501 ( .A1(n449), .A2(n448), .ZN(n455) );
  XOR2_X1 U502 ( .A(n450), .B(KEYINPUT28), .Z(n508) );
  NAND2_X1 U503 ( .A1(n499), .A2(n451), .ZN(n530) );
  NOR2_X1 U504 ( .A1(n508), .A2(n530), .ZN(n513) );
  XOR2_X1 U505 ( .A(n513), .B(KEYINPUT92), .Z(n452) );
  NOR2_X1 U506 ( .A1(n505), .A2(n452), .ZN(n453) );
  XOR2_X1 U507 ( .A(KEYINPUT93), .B(n453), .Z(n454) );
  NOR2_X1 U508 ( .A1(n455), .A2(n454), .ZN(n467) );
  NOR2_X1 U509 ( .A1(n538), .A2(n456), .ZN(n457) );
  XOR2_X1 U510 ( .A(KEYINPUT16), .B(n457), .Z(n458) );
  NOR2_X1 U511 ( .A1(n467), .A2(n458), .ZN(n459) );
  XOR2_X1 U512 ( .A(KEYINPUT96), .B(n459), .Z(n483) );
  INV_X1 U513 ( .A(n556), .ZN(n482) );
  OR2_X1 U514 ( .A1(n561), .A2(n482), .ZN(n471) );
  NOR2_X1 U515 ( .A1(n483), .A2(n471), .ZN(n465) );
  NAND2_X1 U516 ( .A1(n465), .A2(n499), .ZN(n460) );
  XNOR2_X1 U517 ( .A(n461), .B(n460), .ZN(G1324GAT) );
  NAND2_X1 U518 ( .A1(n465), .A2(n502), .ZN(n462) );
  XNOR2_X1 U519 ( .A(n462), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U520 ( .A(G15GAT), .B(KEYINPUT35), .Z(n464) );
  NAND2_X1 U521 ( .A1(n465), .A2(n505), .ZN(n463) );
  XNOR2_X1 U522 ( .A(n464), .B(n463), .ZN(G1326GAT) );
  NAND2_X1 U523 ( .A1(n465), .A2(n508), .ZN(n466) );
  XNOR2_X1 U524 ( .A(n466), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U525 ( .A(KEYINPUT97), .B(KEYINPUT37), .Z(n470) );
  NOR2_X1 U526 ( .A1(n467), .A2(n564), .ZN(n468) );
  NAND2_X1 U527 ( .A1(n468), .A2(n567), .ZN(n469) );
  XOR2_X1 U528 ( .A(n470), .B(n469), .Z(n498) );
  OR2_X1 U529 ( .A1(n498), .A2(n471), .ZN(n473) );
  XOR2_X1 U530 ( .A(KEYINPUT38), .B(KEYINPUT98), .Z(n472) );
  XNOR2_X1 U531 ( .A(n473), .B(n472), .ZN(n480) );
  NAND2_X1 U532 ( .A1(n480), .A2(n499), .ZN(n475) );
  XOR2_X1 U533 ( .A(G29GAT), .B(KEYINPUT39), .Z(n474) );
  XNOR2_X1 U534 ( .A(n475), .B(n474), .ZN(G1328GAT) );
  XOR2_X1 U535 ( .A(G36GAT), .B(KEYINPUT99), .Z(n477) );
  NAND2_X1 U536 ( .A1(n480), .A2(n502), .ZN(n476) );
  XNOR2_X1 U537 ( .A(n477), .B(n476), .ZN(G1329GAT) );
  NAND2_X1 U538 ( .A1(n505), .A2(n480), .ZN(n478) );
  XNOR2_X1 U539 ( .A(n478), .B(KEYINPUT40), .ZN(n479) );
  XNOR2_X1 U540 ( .A(G43GAT), .B(n479), .ZN(G1330GAT) );
  NAND2_X1 U541 ( .A1(n480), .A2(n508), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n481), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U543 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n487) );
  XOR2_X1 U544 ( .A(KEYINPUT102), .B(KEYINPUT101), .Z(n485) );
  NAND2_X1 U545 ( .A1(n548), .A2(n482), .ZN(n497) );
  NOR2_X1 U546 ( .A1(n483), .A2(n497), .ZN(n493) );
  NAND2_X1 U547 ( .A1(n493), .A2(n499), .ZN(n484) );
  XNOR2_X1 U548 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U549 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U550 ( .A(KEYINPUT100), .B(n488), .ZN(G1332GAT) );
  XOR2_X1 U551 ( .A(G64GAT), .B(KEYINPUT103), .Z(n490) );
  NAND2_X1 U552 ( .A1(n493), .A2(n502), .ZN(n489) );
  XNOR2_X1 U553 ( .A(n490), .B(n489), .ZN(G1333GAT) );
  NAND2_X1 U554 ( .A1(n505), .A2(n493), .ZN(n491) );
  XNOR2_X1 U555 ( .A(n491), .B(KEYINPUT104), .ZN(n492) );
  XNOR2_X1 U556 ( .A(G71GAT), .B(n492), .ZN(G1334GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT43), .B(KEYINPUT105), .Z(n495) );
  NAND2_X1 U558 ( .A1(n493), .A2(n508), .ZN(n494) );
  XNOR2_X1 U559 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U560 ( .A(G78GAT), .B(n496), .Z(G1335GAT) );
  NOR2_X1 U561 ( .A1(n498), .A2(n497), .ZN(n509) );
  NAND2_X1 U562 ( .A1(n509), .A2(n499), .ZN(n500) );
  XNOR2_X1 U563 ( .A(KEYINPUT106), .B(n500), .ZN(n501) );
  XNOR2_X1 U564 ( .A(G85GAT), .B(n501), .ZN(G1336GAT) );
  XOR2_X1 U565 ( .A(G92GAT), .B(KEYINPUT107), .Z(n504) );
  NAND2_X1 U566 ( .A1(n509), .A2(n502), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n504), .B(n503), .ZN(G1337GAT) );
  NAND2_X1 U568 ( .A1(n505), .A2(n509), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n506), .B(KEYINPUT108), .ZN(n507) );
  XNOR2_X1 U570 ( .A(G99GAT), .B(n507), .ZN(G1338GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT44), .B(KEYINPUT109), .Z(n511) );
  NAND2_X1 U572 ( .A1(n509), .A2(n508), .ZN(n510) );
  XNOR2_X1 U573 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U574 ( .A(G106GAT), .B(n512), .ZN(G1339GAT) );
  XOR2_X1 U575 ( .A(G113GAT), .B(KEYINPUT111), .Z(n517) );
  NAND2_X1 U576 ( .A1(n528), .A2(n513), .ZN(n514) );
  NOR2_X1 U577 ( .A1(n515), .A2(n514), .ZN(n524) );
  NAND2_X1 U578 ( .A1(n524), .A2(n556), .ZN(n516) );
  XNOR2_X1 U579 ( .A(n517), .B(n516), .ZN(G1340GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT112), .B(KEYINPUT49), .Z(n519) );
  NAND2_X1 U581 ( .A1(n524), .A2(n548), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U583 ( .A(G120GAT), .B(n520), .ZN(G1341GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT113), .B(KEYINPUT50), .Z(n522) );
  NAND2_X1 U585 ( .A1(n524), .A2(n564), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U587 ( .A(G127GAT), .B(n523), .ZN(G1342GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT51), .B(KEYINPUT114), .Z(n526) );
  NAND2_X1 U589 ( .A1(n524), .A2(n538), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U591 ( .A(G134GAT), .B(n527), .ZN(G1343GAT) );
  NAND2_X1 U592 ( .A1(n528), .A2(n553), .ZN(n529) );
  NOR2_X1 U593 ( .A1(n530), .A2(n529), .ZN(n539) );
  NAND2_X1 U594 ( .A1(n539), .A2(n556), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n531), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n533) );
  XNOR2_X1 U597 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U599 ( .A(KEYINPUT53), .B(n534), .Z(n536) );
  NAND2_X1 U600 ( .A1(n539), .A2(n548), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n536), .B(n535), .ZN(G1345GAT) );
  NAND2_X1 U602 ( .A1(n564), .A2(n539), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n537), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U604 ( .A(G162GAT), .B(KEYINPUT117), .Z(n541) );
  NAND2_X1 U605 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(G1347GAT) );
  NAND2_X1 U607 ( .A1(n551), .A2(n556), .ZN(n544) );
  XOR2_X1 U608 ( .A(G169GAT), .B(KEYINPUT119), .Z(n542) );
  XNOR2_X1 U609 ( .A(KEYINPUT120), .B(n542), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(G1348GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n546) );
  XNOR2_X1 U612 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U614 ( .A(KEYINPUT121), .B(n547), .Z(n550) );
  NAND2_X1 U615 ( .A1(n551), .A2(n548), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(G1349GAT) );
  NAND2_X1 U617 ( .A1(n564), .A2(n551), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n552), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U619 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U620 ( .A(KEYINPUT123), .B(n555), .ZN(n568) );
  NAND2_X1 U621 ( .A1(n568), .A2(n556), .ZN(n560) );
  XOR2_X1 U622 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n558) );
  XNOR2_X1 U623 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(G1352GAT) );
  XOR2_X1 U626 ( .A(G204GAT), .B(KEYINPUT61), .Z(n563) );
  NAND2_X1 U627 ( .A1(n568), .A2(n561), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(G1353GAT) );
  XOR2_X1 U629 ( .A(G211GAT), .B(KEYINPUT125), .Z(n566) );
  NAND2_X1 U630 ( .A1(n568), .A2(n564), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(G1354GAT) );
  XNOR2_X1 U632 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n572) );
  XOR2_X1 U633 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n570) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n572), .B(n571), .ZN(G1355GAT) );
endmodule

