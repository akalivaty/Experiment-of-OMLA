//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0 1 0 0 1 0 1 1 1 0 1 0 0 1 1 0 1 1 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n819, new_n820, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973;
  INV_X1    g000(.A(G43gat), .ZN(new_n202));
  INV_X1    g001(.A(G50gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT15), .ZN(new_n205));
  NAND2_X1  g004(.A1(G43gat), .A2(G50gat), .ZN(new_n206));
  AND3_X1   g005(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n205), .B1(new_n204), .B2(new_n206), .ZN(new_n208));
  INV_X1    g007(.A(G29gat), .ZN(new_n209));
  INV_X1    g008(.A(G36gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(new_n210), .A3(KEYINPUT14), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT14), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n212), .B1(G29gat), .B2(G36gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NOR3_X1   g013(.A1(new_n207), .A2(new_n208), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT87), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n209), .A2(KEYINPUT85), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT85), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G29gat), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n216), .B1(new_n220), .B2(new_n210), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n210), .B1(new_n217), .B2(new_n219), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT87), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n215), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n208), .B1(new_n222), .B2(new_n214), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT86), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI211_X1 g026(.A(KEYINPUT86), .B(new_n208), .C1(new_n222), .C2(new_n214), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n224), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT17), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n224), .B(KEYINPUT17), .C1(new_n227), .C2(new_n229), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT8), .ZN(new_n234));
  NAND2_X1  g033(.A1(G99gat), .A2(G106gat), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n234), .B1(new_n235), .B2(KEYINPUT97), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT97), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n237), .A2(G99gat), .A3(G106gat), .ZN(new_n238));
  INV_X1    g037(.A(G85gat), .ZN(new_n239));
  INV_X1    g038(.A(G92gat), .ZN(new_n240));
  AOI22_X1  g039(.A1(new_n236), .A2(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT7), .ZN(new_n242));
  OAI211_X1 g041(.A(KEYINPUT96), .B(new_n242), .C1(new_n239), .C2(new_n240), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT96), .B1(new_n239), .B2(new_n240), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT96), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n245), .A2(G85gat), .A3(G92gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n244), .A2(new_n246), .A3(KEYINPUT7), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n241), .A2(new_n243), .A3(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(G99gat), .B(G106gat), .Z(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n249), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n241), .A2(new_n251), .A3(new_n243), .A4(new_n247), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n232), .A2(new_n233), .A3(new_n253), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n250), .A2(new_n252), .ZN(new_n255));
  AND2_X1   g054(.A1(G232gat), .A2(G233gat), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n255), .A2(new_n230), .B1(KEYINPUT41), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G190gat), .B(G218gat), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT98), .ZN(new_n260));
  OR2_X1    g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G134gat), .B(G162gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n259), .A2(new_n260), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n256), .A2(KEYINPUT41), .ZN(new_n266));
  XOR2_X1   g065(.A(new_n265), .B(new_n266), .Z(new_n267));
  INV_X1    g066(.A(new_n263), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n258), .A2(new_n268), .A3(new_n261), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n264), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n267), .B1(new_n264), .B2(new_n269), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G22gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(G15gat), .ZN(new_n275));
  INV_X1    g074(.A(G15gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G22gat), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT88), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n275), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(G1gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G15gat), .B(G22gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n282), .A2(new_n278), .A3(G1gat), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT16), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n281), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(G8gat), .ZN(new_n287));
  AOI22_X1  g086(.A1(new_n279), .A2(new_n280), .B1(new_n282), .B2(new_n284), .ZN(new_n288));
  INV_X1    g087(.A(G8gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n288), .A2(new_n289), .A3(new_n283), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n292));
  OR2_X1    g091(.A1(new_n292), .A2(KEYINPUT94), .ZN(new_n293));
  XOR2_X1   g092(.A(G57gat), .B(G64gat), .Z(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(KEYINPUT94), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(G71gat), .B(G78gat), .Z(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n297), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n299), .A2(new_n293), .A3(new_n294), .A4(new_n295), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n291), .B1(KEYINPUT21), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G183gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n303), .B(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT95), .B(KEYINPUT21), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n305), .B(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G127gat), .B(G155gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(G231gat), .A2(G233gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G211gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n313), .B(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n310), .B(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G120gat), .B(G148gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(G176gat), .ZN(new_n318));
  INV_X1    g117(.A(G204gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G230gat), .A2(G233gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n253), .A2(new_n301), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT99), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n250), .A2(new_n298), .A3(new_n300), .A4(new_n252), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n253), .A2(KEYINPUT99), .A3(new_n301), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT10), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT100), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n255), .A2(new_n328), .A3(KEYINPUT10), .A4(new_n302), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT10), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT100), .B1(new_n324), .B2(new_n330), .ZN(new_n331));
  AND2_X1   g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n321), .B1(new_n327), .B2(new_n332), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n325), .A2(new_n326), .ZN(new_n334));
  INV_X1    g133(.A(new_n321), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n320), .B1(new_n333), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n333), .A2(new_n336), .A3(new_n320), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT101), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT101), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n333), .A2(new_n340), .A3(new_n336), .A4(new_n320), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n337), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n273), .A2(new_n316), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT93), .ZN(new_n344));
  NAND2_X1  g143(.A1(G227gat), .A2(G233gat), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(G113gat), .ZN(new_n347));
  INV_X1    g146(.A(G120gat), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT1), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n349), .B1(new_n347), .B2(new_n348), .ZN(new_n350));
  XOR2_X1   g149(.A(G127gat), .B(G134gat), .Z(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT66), .ZN(new_n353));
  INV_X1    g152(.A(G190gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n304), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n355), .B(new_n356), .C1(new_n357), .C2(KEYINPUT65), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n357), .A2(KEYINPUT65), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(G169gat), .A2(G176gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT23), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT23), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n363), .B1(G169gat), .B2(G176gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(G169gat), .A2(G176gat), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n362), .A2(KEYINPUT25), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n353), .B1(new_n360), .B2(new_n366), .ZN(new_n367));
  OR2_X1    g166(.A1(new_n357), .A2(KEYINPUT65), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n355), .A2(new_n356), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n357), .A2(KEYINPUT65), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n366), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n371), .A2(new_n372), .A3(KEYINPUT66), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n367), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT25), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n362), .A2(new_n365), .A3(new_n364), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n355), .A2(new_n356), .ZN(new_n377));
  OAI22_X1  g176(.A1(new_n376), .A2(KEYINPUT64), .B1(new_n357), .B2(new_n377), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n376), .A2(KEYINPUT64), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n375), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n365), .ZN(new_n381));
  INV_X1    g180(.A(new_n361), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n381), .B1(new_n382), .B2(KEYINPUT26), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT26), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n361), .A2(new_n384), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n383), .A2(new_n385), .B1(G183gat), .B2(G190gat), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT27), .B(G183gat), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n388), .A2(KEYINPUT28), .A3(new_n354), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT68), .ZN(new_n390));
  NAND2_X1  g189(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n391));
  AOI21_X1  g190(.A(G190gat), .B1(new_n391), .B2(KEYINPUT27), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT27), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n393), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n394));
  AOI211_X1 g193(.A(new_n390), .B(KEYINPUT28), .C1(new_n392), .C2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n391), .A2(KEYINPUT27), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n396), .A2(new_n394), .A3(new_n354), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT28), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT68), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n389), .B1(new_n395), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT69), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n387), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI211_X1 g201(.A(KEYINPUT69), .B(new_n389), .C1(new_n395), .C2(new_n399), .ZN(new_n403));
  AOI221_X4 g202(.A(new_n352), .B1(new_n374), .B2(new_n380), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n350), .A2(new_n351), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n350), .A2(new_n351), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n400), .A2(new_n401), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n408), .A2(new_n403), .A3(new_n386), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n374), .A2(new_n380), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n407), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n346), .B1(new_n404), .B2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G15gat), .B(G43gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(G71gat), .B(G99gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT33), .ZN(new_n416));
  OR2_X1    g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n412), .A2(KEYINPUT32), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT71), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT71), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n412), .A2(new_n420), .A3(KEYINPUT32), .A4(new_n417), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT70), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n409), .A2(new_n410), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n352), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n409), .A2(new_n407), .A3(new_n410), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n345), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n423), .B1(new_n427), .B2(KEYINPUT33), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n415), .B1(new_n412), .B2(KEYINPUT32), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n412), .A2(KEYINPUT70), .A3(new_n416), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n422), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n425), .A2(new_n345), .A3(new_n426), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT72), .ZN(new_n434));
  XNOR2_X1  g233(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n435));
  OR2_X1    g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n435), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n432), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n422), .A2(new_n431), .A3(new_n436), .A4(new_n437), .ZN(new_n440));
  XNOR2_X1  g239(.A(G155gat), .B(G162gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(G141gat), .B(G148gat), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT2), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n441), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(G155gat), .ZN(new_n446));
  INV_X1    g245(.A(G162gat), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT2), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT75), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT75), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n450), .B(KEYINPUT2), .C1(new_n446), .C2(new_n447), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n449), .A2(new_n441), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(G148gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(G141gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(KEYINPUT74), .B(G141gat), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n454), .B1(new_n455), .B2(new_n453), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n445), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(G197gat), .B(G204gat), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT22), .ZN(new_n459));
  INV_X1    g258(.A(G218gat), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n459), .B1(new_n314), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  XOR2_X1   g261(.A(G211gat), .B(G218gat), .Z(new_n463));
  XNOR2_X1  g262(.A(new_n462), .B(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT29), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT3), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n457), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n441), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n469), .B1(KEYINPUT2), .B2(new_n442), .ZN(new_n470));
  INV_X1    g269(.A(new_n456), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n449), .A2(new_n441), .A3(new_n451), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n467), .B(new_n470), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n464), .B1(new_n473), .B2(new_n465), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT79), .B1(new_n468), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n475), .A2(G228gat), .A3(G233gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(G228gat), .A2(G233gat), .ZN(new_n477));
  OAI211_X1 g276(.A(KEYINPUT79), .B(new_n477), .C1(new_n468), .C2(new_n474), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(G22gat), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT80), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n476), .A2(new_n274), .A3(new_n478), .ZN(new_n482));
  XNOR2_X1  g281(.A(G78gat), .B(G106gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n483), .B(KEYINPUT31), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n484), .B(new_n203), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n480), .A2(new_n481), .A3(new_n482), .A4(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n482), .A2(KEYINPUT80), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n488), .A2(new_n485), .B1(new_n480), .B2(new_n482), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n439), .A2(new_n440), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT76), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n492), .B1(new_n457), .B2(new_n407), .ZN(new_n493));
  NAND2_X1  g292(.A1(G225gat), .A2(G233gat), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n496), .A2(new_n352), .A3(KEYINPUT76), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n493), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n457), .A2(new_n407), .B1(KEYINPUT4), .B2(new_n494), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n457), .A2(KEYINPUT4), .A3(new_n407), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n457), .A2(new_n467), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n473), .A2(new_n352), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n498), .A2(new_n499), .B1(new_n503), .B2(new_n494), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT5), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT4), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n506), .B1(new_n496), .B2(new_n352), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n507), .B(new_n500), .C1(new_n501), .C2(new_n502), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n494), .A2(new_n505), .ZN(new_n509));
  OAI22_X1  g308(.A1(new_n504), .A2(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G1gat), .B(G29gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(KEYINPUT0), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(G57gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(new_n239), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT6), .ZN(new_n517));
  OAI221_X1 g316(.A(new_n514), .B1(new_n508), .B2(new_n509), .C1(new_n504), .C2(new_n505), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT78), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n510), .A2(new_n520), .A3(KEYINPUT6), .A4(new_n515), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n498), .A2(new_n499), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n503), .A2(new_n494), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n505), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n508), .A2(new_n509), .ZN(new_n525));
  OAI211_X1 g324(.A(KEYINPUT6), .B(new_n515), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT78), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n519), .A2(new_n521), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(G226gat), .A2(G233gat), .ZN(new_n529));
  AOI22_X1  g328(.A1(new_n409), .A2(new_n410), .B1(new_n465), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n529), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n531), .B(new_n464), .C1(new_n424), .C2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n464), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n424), .A2(new_n532), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n534), .B1(new_n535), .B2(new_n530), .ZN(new_n536));
  XNOR2_X1  g335(.A(G8gat), .B(G36gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(G64gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(new_n240), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n533), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT30), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n533), .A2(new_n536), .A3(KEYINPUT30), .A4(new_n539), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n533), .A2(new_n536), .ZN(new_n544));
  INV_X1    g343(.A(new_n539), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n542), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n547), .A2(KEYINPUT35), .ZN(new_n548));
  NOR3_X1   g347(.A1(new_n491), .A2(new_n528), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT83), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n491), .A2(new_n550), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n527), .A2(new_n521), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n516), .A2(KEYINPUT77), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n524), .A2(new_n525), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT6), .B1(new_n554), .B2(new_n514), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT77), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n510), .A2(new_n556), .A3(new_n515), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n553), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n552), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n547), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n439), .A2(KEYINPUT83), .A3(new_n490), .A4(new_n440), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n551), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n549), .B1(new_n564), .B2(KEYINPUT35), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n544), .A2(KEYINPUT37), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT37), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n533), .A2(new_n567), .A3(new_n536), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n545), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT38), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT82), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n533), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n544), .A2(new_n572), .A3(KEYINPUT37), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n539), .A2(KEYINPUT38), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n571), .A2(new_n567), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n573), .B(new_n574), .C1(new_n544), .C2(new_n575), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n528), .A2(new_n570), .A3(new_n540), .A4(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n488), .A2(new_n485), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n480), .A2(new_n482), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(new_n486), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT40), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n508), .A2(new_n495), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n493), .A2(new_n497), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n494), .B1(new_n496), .B2(new_n352), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n583), .B(KEYINPUT39), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT39), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n508), .A2(new_n587), .A3(new_n495), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n586), .A2(new_n514), .A3(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n516), .B1(new_n582), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n582), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT81), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n589), .A2(KEYINPUT81), .A3(new_n582), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n590), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n581), .B1(new_n595), .B2(new_n547), .ZN(new_n596));
  AOI22_X1  g395(.A1(new_n577), .A2(new_n596), .B1(new_n561), .B2(new_n581), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n439), .A2(new_n440), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT36), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n439), .A2(KEYINPUT36), .A3(new_n440), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n565), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n230), .A2(new_n291), .ZN(new_n605));
  NAND2_X1  g404(.A1(G229gat), .A2(G233gat), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n287), .A2(KEYINPUT89), .A3(new_n290), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n221), .A2(new_n223), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n225), .A2(new_n226), .ZN(new_n609));
  AOI22_X1  g408(.A1(new_n608), .A2(new_n215), .B1(new_n609), .B2(new_n228), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n607), .B1(new_n610), .B2(KEYINPUT17), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT89), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n286), .A2(G8gat), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n289), .B1(new_n288), .B2(new_n283), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n233), .A2(new_n615), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n605), .B(new_n606), .C1(new_n611), .C2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n605), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n230), .A2(new_n291), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n606), .B(KEYINPUT13), .Z(new_n622));
  AOI22_X1  g421(.A1(new_n618), .A2(KEYINPUT18), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n617), .A2(KEYINPUT90), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT18), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n232), .A2(new_n607), .A3(new_n233), .A4(new_n615), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT90), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n626), .A2(new_n627), .A3(new_n605), .A4(new_n606), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n624), .A2(new_n625), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n623), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT91), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n622), .B1(new_n619), .B2(new_n620), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n631), .B(new_n632), .C1(new_n617), .C2(new_n625), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n634));
  XNOR2_X1  g433(.A(G113gat), .B(G141gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G169gat), .B(G197gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT12), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n630), .A2(new_n633), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n633), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n641), .A2(new_n623), .A3(new_n629), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n640), .A2(KEYINPUT92), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(KEYINPUT92), .B1(new_n640), .B2(new_n642), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n344), .B1(new_n604), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n645), .ZN(new_n647));
  OAI211_X1 g446(.A(KEYINPUT93), .B(new_n647), .C1(new_n565), .C2(new_n603), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n343), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n559), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g450(.A(KEYINPUT102), .B(G1gat), .Z(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(G1324gat));
  AOI211_X1 g452(.A(new_n560), .B(new_n343), .C1(new_n646), .C2(new_n648), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT16), .B(G8gat), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n654), .A2(KEYINPUT103), .A3(KEYINPUT42), .A4(new_n656), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n649), .A2(KEYINPUT42), .A3(new_n547), .A4(new_n656), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT103), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n649), .A2(new_n547), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n661), .B1(new_n662), .B2(G8gat), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n655), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n657), .B(new_n660), .C1(new_n663), .C2(new_n664), .ZN(G1325gat));
  INV_X1    g464(.A(new_n649), .ZN(new_n666));
  OAI21_X1  g465(.A(G15gat), .B1(new_n666), .B2(new_n602), .ZN(new_n667));
  INV_X1    g466(.A(new_n598), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n649), .A2(new_n276), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(G1326gat));
  NAND2_X1  g469(.A1(new_n649), .A2(new_n581), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT43), .B(G22gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1327gat));
  NAND2_X1  g472(.A1(new_n646), .A2(new_n648), .ZN(new_n674));
  INV_X1    g473(.A(new_n342), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n675), .A2(new_n273), .A3(new_n316), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n674), .A2(new_n650), .A3(new_n220), .A4(new_n676), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n677), .A2(KEYINPUT45), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(KEYINPUT45), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n630), .B(new_n641), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n316), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n681), .A2(new_n682), .A3(new_n342), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n272), .B1(new_n565), .B2(new_n603), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT44), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n686), .B(new_n272), .C1(new_n565), .C2(new_n603), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n683), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n688), .A2(new_n650), .ZN(new_n689));
  OAI22_X1  g488(.A1(new_n678), .A2(new_n679), .B1(new_n220), .B2(new_n689), .ZN(G1328gat));
  NAND4_X1  g489(.A1(new_n674), .A2(new_n210), .A3(new_n547), .A4(new_n676), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT46), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n688), .A2(new_n547), .ZN(new_n695));
  OAI22_X1  g494(.A1(new_n693), .A2(new_n694), .B1(new_n210), .B2(new_n695), .ZN(G1329gat));
  INV_X1    g495(.A(KEYINPUT47), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n674), .A2(new_n202), .A3(new_n668), .A4(new_n676), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n602), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n202), .B1(new_n688), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n697), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n688), .A2(new_n700), .ZN(new_n703));
  OAI211_X1 g502(.A(KEYINPUT47), .B(new_n698), .C1(new_n703), .C2(new_n202), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(G1330gat));
  INV_X1    g504(.A(KEYINPUT48), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n674), .A2(new_n203), .A3(new_n581), .A4(new_n676), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n203), .B1(new_n688), .B2(new_n581), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n706), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n688), .A2(new_n581), .ZN(new_n711));
  OAI211_X1 g510(.A(KEYINPUT48), .B(new_n707), .C1(new_n711), .C2(new_n203), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(G1331gat));
  INV_X1    g512(.A(KEYINPUT104), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n680), .A2(new_n675), .A3(new_n316), .A4(new_n273), .ZN(new_n715));
  OR3_X1    g514(.A1(new_n604), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n714), .B1(new_n604), .B2(new_n715), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n650), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g520(.A(KEYINPUT49), .B(G64gat), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n719), .A2(new_n547), .A3(new_n722), .ZN(new_n723));
  OAI22_X1  g522(.A1(new_n718), .A2(new_n560), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(G1333gat));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n598), .B(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n716), .A2(new_n717), .A3(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(G71gat), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n700), .A2(G71gat), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n718), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT50), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n729), .A2(new_n730), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT50), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n735), .B(new_n736), .C1(new_n718), .C2(new_n732), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n734), .A2(new_n737), .ZN(G1334gat));
  NAND2_X1  g537(.A1(new_n719), .A2(new_n581), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(G78gat), .ZN(G1335gat));
  OR2_X1    g539(.A1(new_n565), .A2(new_n603), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n681), .A2(new_n316), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n741), .A2(KEYINPUT51), .A3(new_n272), .A4(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT51), .ZN(new_n744));
  INV_X1    g543(.A(new_n742), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n684), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n342), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n747), .A2(new_n239), .A3(new_n650), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n742), .A2(new_n675), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n749), .B1(new_n685), .B2(new_n687), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n750), .A2(new_n650), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n748), .B1(new_n239), .B2(new_n751), .ZN(G1336gat));
  NOR2_X1   g551(.A1(new_n560), .A2(G92gat), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT52), .B1(new_n747), .B2(new_n753), .ZN(new_n754));
  AOI211_X1 g553(.A(new_n560), .B(new_n749), .C1(new_n685), .C2(new_n687), .ZN(new_n755));
  OAI21_X1  g554(.A(G92gat), .B1(new_n755), .B2(KEYINPUT106), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n750), .A2(KEYINPUT106), .A3(new_n547), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n754), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n753), .ZN(new_n759));
  AOI211_X1 g558(.A(new_n342), .B(new_n759), .C1(new_n743), .C2(new_n746), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n240), .B1(new_n750), .B2(new_n547), .ZN(new_n761));
  OAI21_X1  g560(.A(KEYINPUT52), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n758), .A2(new_n762), .ZN(G1337gat));
  AOI21_X1  g562(.A(G99gat), .B1(new_n747), .B2(new_n668), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n700), .A2(G99gat), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n764), .B1(new_n750), .B2(new_n765), .ZN(G1338gat));
  INV_X1    g565(.A(G106gat), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n747), .A2(new_n767), .A3(new_n581), .ZN(new_n768));
  XNOR2_X1  g567(.A(KEYINPUT107), .B(KEYINPUT53), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n750), .A2(new_n581), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n768), .B(new_n769), .C1(new_n767), .C2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n769), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n581), .A2(new_n767), .ZN(new_n773));
  AOI211_X1 g572(.A(new_n342), .B(new_n773), .C1(new_n743), .C2(new_n746), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n767), .B1(new_n750), .B2(new_n581), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n772), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n771), .A2(new_n776), .ZN(G1339gat));
  NOR2_X1   g576(.A1(new_n343), .A2(new_n681), .ZN(new_n778));
  INV_X1    g577(.A(new_n638), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n621), .A2(new_n622), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n606), .B1(new_n626), .B2(new_n605), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n782), .B1(new_n630), .B2(new_n639), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT108), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n783), .B(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n329), .A2(new_n331), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n335), .B(new_n787), .C1(new_n334), .C2(KEYINPUT10), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n788), .A2(KEYINPUT54), .A3(new_n333), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT54), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n790), .B(new_n321), .C1(new_n327), .C2(new_n332), .ZN(new_n791));
  INV_X1    g590(.A(new_n320), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n786), .B1(new_n789), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n339), .A2(new_n341), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n788), .A2(new_n333), .A3(KEYINPUT54), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n796), .A2(KEYINPUT55), .A3(new_n792), .A4(new_n791), .ZN(new_n797));
  AND4_X1   g596(.A1(new_n272), .A2(new_n794), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n785), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n342), .A2(new_n783), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n794), .A2(new_n795), .A3(new_n797), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n800), .B1(new_n801), .B2(new_n681), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n799), .B1(new_n802), .B2(new_n272), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n778), .B1(new_n803), .B2(new_n682), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n804), .A2(new_n559), .ZN(new_n805));
  INV_X1    g604(.A(new_n551), .ZN(new_n806));
  INV_X1    g605(.A(new_n563), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n806), .A2(new_n547), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(G113gat), .B1(new_n810), .B2(new_n681), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n804), .A2(new_n581), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n812), .A2(new_n650), .A3(new_n668), .A4(new_n560), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n813), .A2(new_n347), .A3(new_n645), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n811), .A2(new_n814), .ZN(G1340gat));
  AOI21_X1  g614(.A(G120gat), .B1(new_n810), .B2(new_n675), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n813), .A2(new_n348), .A3(new_n342), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n816), .A2(new_n817), .ZN(G1341gat));
  OAI21_X1  g617(.A(G127gat), .B1(new_n813), .B2(new_n682), .ZN(new_n819));
  OR2_X1    g618(.A1(new_n682), .A2(G127gat), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n819), .B1(new_n809), .B2(new_n820), .ZN(G1342gat));
  OR2_X1    g620(.A1(new_n273), .A2(G134gat), .ZN(new_n822));
  XOR2_X1   g621(.A(KEYINPUT109), .B(KEYINPUT56), .Z(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  OR3_X1    g623(.A1(new_n809), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(G134gat), .B1(new_n813), .B2(new_n273), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n824), .B1(new_n809), .B2(new_n822), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(KEYINPUT110), .ZN(G1343gat));
  AOI211_X1 g628(.A(new_n559), .B(new_n547), .C1(new_n600), .C2(new_n601), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n831), .B1(new_n804), .B2(new_n490), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n581), .A2(KEYINPUT57), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n795), .A2(new_n797), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT111), .B1(new_n789), .B2(new_n793), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT111), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n796), .A2(new_n836), .A3(new_n792), .A4(new_n791), .ZN(new_n837));
  XOR2_X1   g636(.A(KEYINPUT112), .B(KEYINPUT55), .Z(new_n838));
  NAND3_X1  g637(.A1(new_n835), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n834), .B(new_n839), .C1(new_n643), .C2(new_n644), .ZN(new_n840));
  INV_X1    g639(.A(new_n800), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n272), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n799), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n682), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n778), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n833), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT113), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n832), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AOI211_X1 g647(.A(KEYINPUT113), .B(new_n833), .C1(new_n844), .C2(new_n845), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n830), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n455), .B1(new_n850), .B2(new_n645), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n700), .A2(new_n547), .A3(new_n490), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n805), .A2(new_n852), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n853), .A2(G141gat), .A3(new_n645), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  XNOR2_X1  g654(.A(KEYINPUT114), .B(KEYINPUT58), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n851), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT58), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n681), .B(new_n830), .C1(new_n848), .C2(new_n849), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n854), .B1(new_n859), .B2(new_n455), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n857), .B1(new_n858), .B2(new_n860), .ZN(G1344gat));
  NOR2_X1   g660(.A1(new_n490), .A2(KEYINPUT57), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n647), .A2(new_n343), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n863), .B1(new_n844), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n794), .A2(new_n795), .A3(new_n797), .ZN(new_n866));
  OAI22_X1  g665(.A1(new_n866), .A2(new_n680), .B1(new_n342), .B2(new_n783), .ZN(new_n867));
  AOI22_X1  g666(.A1(new_n867), .A2(new_n273), .B1(new_n785), .B2(new_n798), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n845), .B1(new_n868), .B2(new_n316), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n831), .B1(new_n869), .B2(new_n581), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n830), .A2(KEYINPUT115), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n830), .A2(KEYINPUT115), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n342), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n453), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n877));
  OR3_X1    g676(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n877), .B(G148gat), .C1(new_n850), .C2(new_n342), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n876), .B1(new_n875), .B2(new_n877), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n853), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(new_n453), .A3(new_n675), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(new_n883), .ZN(G1345gat));
  OAI21_X1  g683(.A(G155gat), .B1(new_n850), .B2(new_n682), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n882), .A2(new_n446), .A3(new_n316), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(G1346gat));
  OAI211_X1 g686(.A(new_n272), .B(new_n830), .C1(new_n848), .C2(new_n849), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(G162gat), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n882), .A2(new_n447), .A3(new_n272), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n889), .A2(KEYINPUT117), .A3(new_n890), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(G1347gat));
  NAND2_X1  g694(.A1(new_n559), .A2(new_n547), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n806), .A2(new_n807), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n869), .A2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(G169gat), .B1(new_n899), .B2(new_n681), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n727), .A2(new_n896), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n812), .A2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n647), .A2(G169gat), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n900), .B1(new_n903), .B2(new_n904), .ZN(G1348gat));
  AOI21_X1  g704(.A(G176gat), .B1(new_n899), .B2(new_n675), .ZN(new_n906));
  XOR2_X1   g705(.A(new_n906), .B(KEYINPUT118), .Z(new_n907));
  NAND3_X1  g706(.A1(new_n903), .A2(G176gat), .A3(new_n675), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n907), .A2(new_n908), .ZN(G1349gat));
  NAND2_X1  g708(.A1(new_n316), .A2(new_n388), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT119), .B1(new_n898), .B2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT119), .ZN(new_n912));
  INV_X1    g711(.A(new_n910), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n869), .A2(new_n897), .A3(new_n912), .A4(new_n913), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n869), .A2(new_n901), .A3(new_n490), .A4(new_n316), .ZN(new_n915));
  AOI22_X1  g714(.A1(new_n911), .A2(new_n914), .B1(G183gat), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT120), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(KEYINPUT60), .B1(new_n916), .B2(KEYINPUT120), .ZN(new_n919));
  OAI21_X1  g718(.A(KEYINPUT121), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n916), .A2(KEYINPUT120), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n921), .A2(new_n922), .A3(KEYINPUT60), .A4(new_n917), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT60), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n916), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n920), .A2(new_n923), .A3(new_n925), .ZN(G1350gat));
  OAI21_X1  g725(.A(G190gat), .B1(new_n902), .B2(new_n273), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n928), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n898), .A2(G190gat), .A3(new_n273), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT122), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n929), .A2(new_n930), .A3(new_n932), .ZN(G1351gat));
  INV_X1    g732(.A(G197gat), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n844), .A2(new_n864), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n862), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n937));
  OAI21_X1  g736(.A(KEYINPUT57), .B1(new_n804), .B2(new_n490), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(KEYINPUT124), .B1(new_n865), .B2(new_n870), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n700), .A2(new_n896), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n939), .A2(new_n940), .A3(new_n647), .A4(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n934), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n944), .B1(new_n943), .B2(new_n942), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n700), .A2(new_n490), .ZN(new_n946));
  INV_X1    g745(.A(new_n896), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n946), .A2(new_n869), .A3(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n949), .A2(new_n934), .A3(new_n681), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT123), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n945), .A2(new_n951), .ZN(G1352gat));
  NAND4_X1  g751(.A1(new_n939), .A2(new_n940), .A3(new_n675), .A4(new_n941), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(G204gat), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n948), .A2(G204gat), .A3(new_n342), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT62), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(KEYINPUT126), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT126), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n954), .A2(new_n959), .A3(new_n956), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(G1353gat));
  NAND3_X1  g760(.A1(new_n949), .A2(new_n314), .A3(new_n316), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n871), .A2(new_n316), .A3(new_n941), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n963), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n964));
  AOI21_X1  g763(.A(KEYINPUT63), .B1(new_n963), .B2(G211gat), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(G1354gat));
  NAND4_X1  g765(.A1(new_n939), .A2(new_n940), .A3(new_n272), .A4(new_n941), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(G218gat), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n949), .A2(new_n460), .A3(new_n272), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(KEYINPUT127), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT127), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n968), .A2(new_n972), .A3(new_n969), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n971), .A2(new_n973), .ZN(G1355gat));
endmodule


