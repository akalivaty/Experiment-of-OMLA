

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725;

  NOR2_X1 U370 ( .A1(n675), .A2(n694), .ZN(n368) );
  NOR2_X1 U371 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U372 ( .A(n347), .B(n693), .ZN(n695) );
  XNOR2_X1 U373 ( .A(n673), .B(n674), .ZN(n675) );
  AND2_X1 U374 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U375 ( .A1(n591), .A2(n590), .ZN(n595) );
  OR2_X1 U376 ( .A1(n633), .A2(G902), .ZN(n395) );
  XNOR2_X1 U377 ( .A(n463), .B(n415), .ZN(n389) );
  NAND2_X1 U378 ( .A1(n348), .A2(G217), .ZN(n347) );
  XNOR2_X2 U379 ( .A(n582), .B(KEYINPUT6), .ZN(n574) );
  INV_X2 U380 ( .A(G128), .ZN(n385) );
  XNOR2_X2 U381 ( .A(n410), .B(n373), .ZN(n390) );
  XNOR2_X1 U382 ( .A(n634), .B(KEYINPUT2), .ZN(n636) );
  XNOR2_X1 U383 ( .A(n387), .B(KEYINPUT39), .ZN(n611) );
  NAND2_X1 U384 ( .A1(n372), .A2(n370), .ZN(n614) );
  XNOR2_X1 U385 ( .A(n395), .B(G472), .ZN(n589) );
  XNOR2_X1 U386 ( .A(n386), .B(n439), .ZN(n571) );
  INV_X2 U387 ( .A(G122), .ZN(n365) );
  NOR2_X1 U388 ( .A1(n723), .A2(n557), .ZN(n558) );
  NOR2_X1 U389 ( .A1(n636), .A2(n635), .ZN(n348) );
  NOR2_X1 U390 ( .A1(n636), .A2(n635), .ZN(n349) );
  BUF_X1 U391 ( .A(n577), .Z(n350) );
  NOR2_X1 U392 ( .A1(n636), .A2(n635), .ZN(n691) );
  OR2_X1 U393 ( .A1(n571), .A2(n492), .ZN(n553) );
  NAND2_X1 U394 ( .A1(n378), .A2(n376), .ZN(n375) );
  AND2_X1 U395 ( .A1(n377), .A2(G469), .ZN(n376) );
  INV_X1 U396 ( .A(G902), .ZN(n377) );
  AND2_X1 U397 ( .A1(n381), .A2(n380), .ZN(n379) );
  NAND2_X1 U398 ( .A1(n382), .A2(G902), .ZN(n380) );
  INV_X1 U399 ( .A(G469), .ZN(n382) );
  NOR2_X1 U400 ( .A1(n719), .A2(n725), .ZN(n608) );
  XNOR2_X1 U401 ( .A(n404), .B(n443), .ZN(n403) );
  AND2_X1 U402 ( .A1(n450), .A2(G210), .ZN(n404) );
  XNOR2_X1 U403 ( .A(n402), .B(n401), .ZN(n400) );
  INV_X1 U404 ( .A(KEYINPUT5), .ZN(n401) );
  XNOR2_X1 U405 ( .A(KEYINPUT87), .B(KEYINPUT70), .ZN(n402) );
  XNOR2_X1 U406 ( .A(n389), .B(n416), .ZN(n374) );
  XNOR2_X1 U407 ( .A(G131), .B(G134), .ZN(n416) );
  OR2_X1 U408 ( .A1(G237), .A2(G902), .ZN(n486) );
  XNOR2_X1 U409 ( .A(G902), .B(KEYINPUT15), .ZN(n635) );
  XNOR2_X1 U410 ( .A(n374), .B(G146), .ZN(n447) );
  XNOR2_X1 U411 ( .A(n704), .B(n405), .ZN(n670) );
  XNOR2_X1 U412 ( .A(n407), .B(n406), .ZN(n405) );
  XNOR2_X1 U413 ( .A(n412), .B(n483), .ZN(n406) );
  XNOR2_X1 U414 ( .A(n389), .B(n484), .ZN(n407) );
  XNOR2_X1 U415 ( .A(n487), .B(n362), .ZN(n606) );
  INV_X1 U416 ( .A(KEYINPUT97), .ZN(n592) );
  XNOR2_X1 U417 ( .A(n584), .B(n585), .ZN(n586) );
  INV_X1 U418 ( .A(KEYINPUT22), .ZN(n373) );
  AND2_X1 U419 ( .A1(n538), .A2(n572), .ZN(n539) );
  NAND2_X1 U420 ( .A1(n369), .A2(n425), .ZN(n372) );
  AND2_X1 U421 ( .A1(n375), .A2(KEYINPUT1), .ZN(n371) );
  INV_X1 U422 ( .A(G953), .ZN(n711) );
  NOR2_X1 U423 ( .A1(G952), .A2(n711), .ZN(n694) );
  NAND2_X1 U424 ( .A1(n351), .A2(n364), .ZN(n363) );
  NOR2_X1 U425 ( .A1(n598), .A2(n654), .ZN(n599) );
  XNOR2_X1 U426 ( .A(G125), .B(G146), .ZN(n482) );
  NAND2_X1 U427 ( .A1(G234), .A2(G237), .ZN(n517) );
  XNOR2_X1 U428 ( .A(KEYINPUT83), .B(KEYINPUT81), .ZN(n481) );
  AND2_X1 U429 ( .A1(G224), .A2(n711), .ZN(n412) );
  INV_X1 U430 ( .A(n668), .ZN(n620) );
  NAND2_X1 U431 ( .A1(n504), .A2(n615), .ZN(n503) );
  XNOR2_X1 U432 ( .A(n383), .B(n360), .ZN(n530) );
  NAND2_X1 U433 ( .A1(n384), .A2(n391), .ZN(n383) );
  XNOR2_X1 U434 ( .A(n488), .B(KEYINPUT95), .ZN(n384) );
  XNOR2_X1 U435 ( .A(n403), .B(n400), .ZN(n444) );
  XOR2_X1 U436 ( .A(KEYINPUT23), .B(KEYINPUT85), .Z(n431) );
  XNOR2_X1 U437 ( .A(KEYINPUT77), .B(KEYINPUT8), .ZN(n433) );
  XOR2_X1 U438 ( .A(KEYINPUT73), .B(G104), .Z(n418) );
  XNOR2_X1 U439 ( .A(n394), .B(KEYINPUT30), .ZN(n590) );
  NOR2_X1 U440 ( .A1(n553), .A2(n369), .ZN(n593) );
  XNOR2_X1 U441 ( .A(n409), .B(n408), .ZN(n704) );
  XNOR2_X1 U442 ( .A(n480), .B(n474), .ZN(n408) );
  XOR2_X1 U443 ( .A(KEYINPUT69), .B(KEYINPUT16), .Z(n474) );
  XNOR2_X1 U444 ( .A(n396), .B(KEYINPUT118), .ZN(n626) );
  NAND2_X1 U445 ( .A1(n397), .A2(n357), .ZN(n396) );
  NAND2_X1 U446 ( .A1(n352), .A2(n625), .ZN(n397) );
  XNOR2_X1 U447 ( .A(n393), .B(n361), .ZN(n719) );
  XNOR2_X1 U448 ( .A(n399), .B(n398), .ZN(n725) );
  INV_X1 U449 ( .A(KEYINPUT40), .ZN(n398) );
  XNOR2_X1 U450 ( .A(KEYINPUT32), .B(n544), .ZN(n724) );
  NOR2_X1 U451 ( .A1(n605), .A2(n388), .ZN(n655) );
  NOR2_X1 U452 ( .A1(n685), .A2(n694), .ZN(n366) );
  XNOR2_X1 U453 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X1 U454 ( .A(n676), .B(n367), .ZN(n679) );
  XNOR2_X1 U455 ( .A(n678), .B(n677), .ZN(n367) );
  OR2_X1 U456 ( .A1(n604), .A2(n603), .ZN(n351) );
  AND2_X1 U457 ( .A1(n624), .A2(n413), .ZN(n352) );
  XOR2_X1 U458 ( .A(n424), .B(n423), .Z(n353) );
  XOR2_X1 U459 ( .A(G113), .B(G101), .Z(n354) );
  XOR2_X1 U460 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n355) );
  AND2_X1 U461 ( .A1(G210), .A2(n486), .ZN(n356) );
  AND2_X1 U462 ( .A1(n521), .A2(n520), .ZN(n357) );
  AND2_X1 U463 ( .A1(n504), .A2(n595), .ZN(n358) );
  AND2_X1 U464 ( .A1(n379), .A2(n375), .ZN(n359) );
  XOR2_X1 U465 ( .A(KEYINPUT33), .B(KEYINPUT67), .Z(n360) );
  XNOR2_X1 U466 ( .A(KEYINPUT100), .B(KEYINPUT42), .ZN(n361) );
  XOR2_X1 U467 ( .A(KEYINPUT99), .B(KEYINPUT41), .Z(n362) );
  NOR2_X1 U468 ( .A1(n600), .A2(n363), .ZN(n610) );
  INV_X1 U469 ( .A(n665), .ZN(n364) );
  NAND2_X1 U470 ( .A1(n571), .A2(n572), .ZN(n573) );
  XNOR2_X1 U471 ( .A(n432), .B(n431), .ZN(n436) );
  XNOR2_X2 U472 ( .A(n365), .B(G104), .ZN(n476) );
  NOR2_X2 U473 ( .A1(n582), .A2(n541), .ZN(n650) );
  XNOR2_X1 U474 ( .A(n366), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U475 ( .A1(n639), .A2(n694), .ZN(n642) );
  INV_X1 U476 ( .A(n574), .ZN(n391) );
  XNOR2_X1 U477 ( .A(n368), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U478 ( .A(n353), .B(n447), .ZN(n678) );
  NAND2_X1 U479 ( .A1(n379), .A2(n375), .ZN(n369) );
  NAND2_X1 U480 ( .A1(n371), .A2(n379), .ZN(n370) );
  AND2_X1 U481 ( .A1(n390), .A2(n580), .ZN(n540) );
  AND2_X1 U482 ( .A1(n390), .A2(n574), .ZN(n543) );
  XNOR2_X1 U483 ( .A(n374), .B(KEYINPUT125), .ZN(n709) );
  INV_X1 U484 ( .A(n678), .ZN(n378) );
  NAND2_X1 U485 ( .A1(n678), .A2(n382), .ZN(n381) );
  NAND2_X1 U486 ( .A1(n530), .A2(n554), .ZN(n532) );
  XNOR2_X2 U487 ( .A(n385), .B(G143), .ZN(n463) );
  NOR2_X1 U488 ( .A1(n693), .A2(G902), .ZN(n386) );
  INV_X1 U489 ( .A(n553), .ZN(n489) );
  NAND2_X1 U490 ( .A1(n594), .A2(n595), .ZN(n607) );
  NAND2_X1 U491 ( .A1(n594), .A2(n358), .ZN(n387) );
  NOR2_X2 U492 ( .A1(n388), .A2(n529), .ZN(n411) );
  XNOR2_X2 U493 ( .A(n577), .B(n528), .ZN(n388) );
  NAND2_X1 U494 ( .A1(n390), .A2(n549), .ZN(n550) );
  INV_X1 U495 ( .A(n392), .ZN(n618) );
  NAND2_X1 U496 ( .A1(n392), .A2(n615), .ZN(n527) );
  XNOR2_X2 U497 ( .A(n485), .B(n356), .ZN(n392) );
  XNOR2_X1 U498 ( .A(n618), .B(KEYINPUT38), .ZN(n504) );
  NAND2_X1 U499 ( .A1(n596), .A2(n392), .ZN(n597) );
  XNOR2_X1 U500 ( .A(n478), .B(n475), .ZN(n409) );
  NOR2_X1 U501 ( .A1(n606), .A2(n605), .ZN(n393) );
  NAND2_X1 U502 ( .A1(n589), .A2(n615), .ZN(n394) );
  NAND2_X1 U503 ( .A1(n611), .A2(n659), .ZN(n399) );
  NAND2_X1 U504 ( .A1(n554), .A2(n539), .ZN(n410) );
  XNOR2_X2 U505 ( .A(n411), .B(KEYINPUT0), .ZN(n554) );
  NAND2_X1 U506 ( .A1(n543), .A2(n542), .ZN(n544) );
  OR2_X1 U507 ( .A1(n623), .A2(KEYINPUT2), .ZN(n413) );
  AND2_X1 U508 ( .A1(n609), .A2(n610), .ZN(n414) );
  INV_X1 U509 ( .A(KEYINPUT4), .ZN(n415) );
  BUF_X1 U510 ( .A(n475), .Z(n445) );
  INV_X1 U511 ( .A(KEYINPUT72), .ZN(n419) );
  NOR2_X1 U512 ( .A1(n720), .A2(n620), .ZN(n621) );
  XNOR2_X1 U513 ( .A(n420), .B(n419), .ZN(n421) );
  INV_X1 U514 ( .A(KEYINPUT79), .ZN(n526) );
  XNOR2_X1 U515 ( .A(n436), .B(n435), .ZN(n438) );
  XNOR2_X1 U516 ( .A(n422), .B(n421), .ZN(n423) );
  INV_X1 U517 ( .A(KEYINPUT19), .ZN(n528) );
  INV_X1 U518 ( .A(KEYINPUT63), .ZN(n640) );
  INV_X1 U519 ( .A(KEYINPUT53), .ZN(n627) );
  XNOR2_X1 U520 ( .A(n640), .B(KEYINPUT104), .ZN(n641) );
  XOR2_X2 U521 ( .A(KEYINPUT71), .B(G110), .Z(n477) );
  XOR2_X1 U522 ( .A(G137), .B(G140), .Z(n437) );
  XNOR2_X1 U523 ( .A(n477), .B(n437), .ZN(n424) );
  XNOR2_X1 U524 ( .A(G101), .B(G107), .ZN(n417) );
  XNOR2_X1 U525 ( .A(n418), .B(n417), .ZN(n422) );
  NAND2_X1 U526 ( .A1(G227), .A2(n711), .ZN(n420) );
  INV_X1 U527 ( .A(KEYINPUT1), .ZN(n425) );
  XOR2_X1 U528 ( .A(KEYINPUT25), .B(KEYINPUT86), .Z(n428) );
  NAND2_X1 U529 ( .A1(G234), .A2(n635), .ZN(n426) );
  XNOR2_X1 U530 ( .A(KEYINPUT20), .B(n426), .ZN(n440) );
  NAND2_X1 U531 ( .A1(G217), .A2(n440), .ZN(n427) );
  XNOR2_X1 U532 ( .A(n428), .B(n427), .ZN(n439) );
  XOR2_X1 U533 ( .A(KEYINPUT24), .B(G128), .Z(n430) );
  XNOR2_X1 U534 ( .A(G119), .B(G110), .ZN(n429) );
  XNOR2_X1 U535 ( .A(n430), .B(n429), .ZN(n432) );
  NAND2_X1 U536 ( .A1(n711), .A2(G234), .ZN(n434) );
  XNOR2_X1 U537 ( .A(n434), .B(n433), .ZN(n467) );
  NAND2_X1 U538 ( .A1(G221), .A2(n467), .ZN(n435) );
  XNOR2_X1 U539 ( .A(KEYINPUT10), .B(n482), .ZN(n455) );
  XNOR2_X1 U540 ( .A(n437), .B(n455), .ZN(n708) );
  XNOR2_X1 U541 ( .A(n438), .B(n708), .ZN(n693) );
  NAND2_X1 U542 ( .A1(G221), .A2(n440), .ZN(n441) );
  XOR2_X1 U543 ( .A(KEYINPUT21), .B(n441), .Z(n572) );
  INV_X1 U544 ( .A(n572), .ZN(n492) );
  NAND2_X1 U545 ( .A1(n614), .A2(n489), .ZN(n488) );
  XNOR2_X1 U546 ( .A(KEYINPUT3), .B(G119), .ZN(n442) );
  XNOR2_X1 U547 ( .A(n354), .B(n442), .ZN(n475) );
  NOR2_X1 U548 ( .A1(G953), .A2(G237), .ZN(n450) );
  XNOR2_X1 U549 ( .A(G116), .B(G137), .ZN(n443) );
  XNOR2_X1 U550 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U551 ( .A(n447), .B(n446), .ZN(n633) );
  BUF_X1 U552 ( .A(n589), .Z(n582) );
  INV_X1 U553 ( .A(n530), .ZN(n511) );
  XNOR2_X1 U554 ( .A(KEYINPUT13), .B(KEYINPUT90), .ZN(n461) );
  XOR2_X1 U555 ( .A(KEYINPUT89), .B(KEYINPUT12), .Z(n449) );
  XNOR2_X1 U556 ( .A(G143), .B(G140), .ZN(n448) );
  XNOR2_X1 U557 ( .A(n449), .B(n448), .ZN(n454) );
  XOR2_X1 U558 ( .A(KEYINPUT11), .B(KEYINPUT88), .Z(n452) );
  NAND2_X1 U559 ( .A1(n450), .A2(G214), .ZN(n451) );
  XNOR2_X1 U560 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U561 ( .A(n454), .B(n453), .ZN(n459) );
  XOR2_X1 U562 ( .A(n455), .B(G131), .Z(n457) );
  XNOR2_X1 U563 ( .A(n476), .B(G113), .ZN(n456) );
  XNOR2_X1 U564 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U565 ( .A(n459), .B(n458), .ZN(n680) );
  NOR2_X1 U566 ( .A1(G902), .A2(n680), .ZN(n460) );
  XNOR2_X1 U567 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U568 ( .A(G475), .B(n462), .ZN(n533) );
  XOR2_X1 U569 ( .A(G116), .B(G107), .Z(n479) );
  XNOR2_X1 U570 ( .A(n479), .B(KEYINPUT91), .ZN(n466) );
  XNOR2_X1 U571 ( .A(G122), .B(n463), .ZN(n464) );
  XNOR2_X1 U572 ( .A(n464), .B(G134), .ZN(n465) );
  XNOR2_X1 U573 ( .A(n466), .B(n465), .ZN(n471) );
  XOR2_X1 U574 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n469) );
  NAND2_X1 U575 ( .A1(G217), .A2(n467), .ZN(n468) );
  XNOR2_X1 U576 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U577 ( .A(n471), .B(n470), .ZN(n688) );
  NOR2_X1 U578 ( .A1(G902), .A2(n688), .ZN(n473) );
  XNOR2_X1 U579 ( .A(KEYINPUT92), .B(G478), .ZN(n472) );
  XNOR2_X1 U580 ( .A(n473), .B(n472), .ZN(n502) );
  INV_X1 U581 ( .A(n502), .ZN(n534) );
  NOR2_X1 U582 ( .A1(n533), .A2(n534), .ZN(n538) );
  INV_X1 U583 ( .A(n538), .ZN(n507) );
  XNOR2_X1 U584 ( .A(n477), .B(n476), .ZN(n478) );
  INV_X1 U585 ( .A(n479), .ZN(n480) );
  XNOR2_X1 U586 ( .A(n355), .B(n481), .ZN(n484) );
  INV_X1 U587 ( .A(n482), .ZN(n483) );
  NAND2_X1 U588 ( .A1(n670), .A2(n635), .ZN(n485) );
  NAND2_X1 U589 ( .A1(G214), .A2(n486), .ZN(n615) );
  NOR2_X1 U590 ( .A1(n507), .A2(n503), .ZN(n487) );
  OR2_X1 U591 ( .A1(n511), .A2(n606), .ZN(n521) );
  INV_X1 U592 ( .A(n582), .ZN(n495) );
  NOR2_X1 U593 ( .A1(n495), .A2(n488), .ZN(n551) );
  XOR2_X1 U594 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n491) );
  INV_X1 U595 ( .A(n614), .ZN(n580) );
  NAND2_X1 U596 ( .A1(n580), .A2(n553), .ZN(n490) );
  XNOR2_X1 U597 ( .A(n491), .B(n490), .ZN(n498) );
  NAND2_X1 U598 ( .A1(n492), .A2(n571), .ZN(n494) );
  XNOR2_X1 U599 ( .A(KEYINPUT49), .B(KEYINPUT113), .ZN(n493) );
  XNOR2_X1 U600 ( .A(n494), .B(n493), .ZN(n496) );
  NAND2_X1 U601 ( .A1(n496), .A2(n495), .ZN(n497) );
  NOR2_X1 U602 ( .A1(n498), .A2(n497), .ZN(n499) );
  NOR2_X1 U603 ( .A1(n551), .A2(n499), .ZN(n500) );
  XOR2_X1 U604 ( .A(KEYINPUT51), .B(n500), .Z(n501) );
  NOR2_X1 U605 ( .A1(n606), .A2(n501), .ZN(n514) );
  NOR2_X1 U606 ( .A1(n502), .A2(n533), .ZN(n661) );
  NAND2_X1 U607 ( .A1(n533), .A2(n502), .ZN(n575) );
  INV_X1 U608 ( .A(n575), .ZN(n659) );
  NOR2_X1 U609 ( .A1(n661), .A2(n659), .ZN(n601) );
  NOR2_X1 U610 ( .A1(n601), .A2(n503), .ZN(n509) );
  NOR2_X1 U611 ( .A1(n504), .A2(n615), .ZN(n505) );
  XOR2_X1 U612 ( .A(KEYINPUT115), .B(n505), .Z(n506) );
  NOR2_X1 U613 ( .A1(n507), .A2(n506), .ZN(n508) );
  NOR2_X1 U614 ( .A1(n509), .A2(n508), .ZN(n510) );
  NOR2_X1 U615 ( .A1(n511), .A2(n510), .ZN(n512) );
  XNOR2_X1 U616 ( .A(n512), .B(KEYINPUT116), .ZN(n513) );
  NOR2_X1 U617 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U618 ( .A(n515), .B(KEYINPUT117), .ZN(n516) );
  XNOR2_X1 U619 ( .A(n516), .B(KEYINPUT52), .ZN(n519) );
  XNOR2_X1 U620 ( .A(n517), .B(KEYINPUT14), .ZN(n523) );
  NAND2_X1 U621 ( .A1(G952), .A2(n523), .ZN(n518) );
  XOR2_X1 U622 ( .A(KEYINPUT84), .B(n518), .Z(n522) );
  NAND2_X1 U623 ( .A1(n519), .A2(n522), .ZN(n520) );
  INV_X1 U624 ( .A(KEYINPUT2), .ZN(n566) );
  AND2_X1 U625 ( .A1(n711), .A2(n522), .ZN(n570) );
  AND2_X1 U626 ( .A1(G953), .A2(n523), .ZN(n524) );
  NAND2_X1 U627 ( .A1(G902), .A2(n524), .ZN(n568) );
  NOR2_X1 U628 ( .A1(G898), .A2(n568), .ZN(n525) );
  NOR2_X1 U629 ( .A1(n570), .A2(n525), .ZN(n529) );
  XNOR2_X2 U630 ( .A(n527), .B(n526), .ZN(n577) );
  XOR2_X1 U631 ( .A(KEYINPUT34), .B(KEYINPUT74), .Z(n531) );
  XNOR2_X1 U632 ( .A(n532), .B(n531), .ZN(n536) );
  AND2_X1 U633 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U634 ( .A(n535), .B(KEYINPUT96), .ZN(n596) );
  NAND2_X1 U635 ( .A1(n536), .A2(n596), .ZN(n537) );
  XNOR2_X1 U636 ( .A(n537), .B(KEYINPUT35), .ZN(n721) );
  NAND2_X1 U637 ( .A1(n540), .A2(n571), .ZN(n541) );
  NOR2_X1 U638 ( .A1(n721), .A2(n650), .ZN(n545) );
  AND2_X1 U639 ( .A1(n571), .A2(n614), .ZN(n542) );
  NAND2_X1 U640 ( .A1(n545), .A2(n724), .ZN(n547) );
  INV_X1 U641 ( .A(KEYINPUT68), .ZN(n559) );
  NOR2_X1 U642 ( .A1(n559), .A2(KEYINPUT44), .ZN(n546) );
  XNOR2_X1 U643 ( .A(n547), .B(n546), .ZN(n563) );
  NOR2_X1 U644 ( .A1(n571), .A2(n614), .ZN(n548) );
  AND2_X1 U645 ( .A1(n574), .A2(n548), .ZN(n549) );
  XNOR2_X1 U646 ( .A(n550), .B(KEYINPUT93), .ZN(n723) );
  NAND2_X1 U647 ( .A1(n554), .A2(n551), .ZN(n552) );
  XNOR2_X1 U648 ( .A(n552), .B(KEYINPUT31), .ZN(n662) );
  NAND2_X1 U649 ( .A1(n593), .A2(n554), .ZN(n555) );
  NOR2_X1 U650 ( .A1(n582), .A2(n555), .ZN(n645) );
  NOR2_X1 U651 ( .A1(n662), .A2(n645), .ZN(n556) );
  NOR2_X1 U652 ( .A1(n601), .A2(n556), .ZN(n557) );
  XNOR2_X1 U653 ( .A(KEYINPUT94), .B(n558), .ZN(n561) );
  NAND2_X1 U654 ( .A1(n559), .A2(KEYINPUT44), .ZN(n560) );
  AND2_X1 U655 ( .A1(n561), .A2(n560), .ZN(n562) );
  NAND2_X1 U656 ( .A1(n563), .A2(n562), .ZN(n565) );
  XOR2_X1 U657 ( .A(KEYINPUT45), .B(KEYINPUT64), .Z(n564) );
  XNOR2_X2 U658 ( .A(n565), .B(n564), .ZN(n697) );
  NAND2_X1 U659 ( .A1(n566), .A2(n697), .ZN(n567) );
  XNOR2_X1 U660 ( .A(n567), .B(KEYINPUT78), .ZN(n625) );
  NOR2_X1 U661 ( .A1(G900), .A2(n568), .ZN(n569) );
  NOR2_X1 U662 ( .A1(n570), .A2(n569), .ZN(n591) );
  NOR2_X1 U663 ( .A1(n591), .A2(n573), .ZN(n583) );
  NOR2_X1 U664 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U665 ( .A1(n583), .A2(n576), .ZN(n613) );
  NOR2_X1 U666 ( .A1(n613), .A2(n350), .ZN(n578) );
  XOR2_X1 U667 ( .A(KEYINPUT36), .B(n578), .Z(n579) );
  NOR2_X1 U668 ( .A1(n580), .A2(n579), .ZN(n665) );
  NAND2_X1 U669 ( .A1(n601), .A2(KEYINPUT47), .ZN(n581) );
  XNOR2_X1 U670 ( .A(n581), .B(KEYINPUT76), .ZN(n588) );
  XOR2_X1 U671 ( .A(KEYINPUT98), .B(KEYINPUT28), .Z(n585) );
  NAND2_X1 U672 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U673 ( .A1(n359), .A2(n586), .ZN(n605) );
  INV_X1 U674 ( .A(n655), .ZN(n602) );
  NAND2_X1 U675 ( .A1(n602), .A2(KEYINPUT47), .ZN(n587) );
  NAND2_X1 U676 ( .A1(n588), .A2(n587), .ZN(n598) );
  XNOR2_X1 U677 ( .A(n593), .B(n592), .ZN(n594) );
  NOR2_X1 U678 ( .A1(n607), .A2(n597), .ZN(n654) );
  XNOR2_X1 U679 ( .A(KEYINPUT75), .B(n599), .ZN(n600) );
  OR2_X1 U680 ( .A1(n602), .A2(n601), .ZN(n604) );
  XNOR2_X1 U681 ( .A(KEYINPUT66), .B(KEYINPUT47), .ZN(n603) );
  XNOR2_X1 U682 ( .A(n608), .B(KEYINPUT46), .ZN(n609) );
  XNOR2_X1 U683 ( .A(n414), .B(KEYINPUT48), .ZN(n622) );
  NAND2_X1 U684 ( .A1(n661), .A2(n611), .ZN(n612) );
  XNOR2_X1 U685 ( .A(KEYINPUT101), .B(n612), .ZN(n720) );
  NOR2_X1 U686 ( .A1(n614), .A2(n613), .ZN(n616) );
  NAND2_X1 U687 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U688 ( .A(n617), .B(KEYINPUT43), .ZN(n619) );
  NAND2_X1 U689 ( .A1(n619), .A2(n618), .ZN(n668) );
  INV_X1 U690 ( .A(n623), .ZN(n710) );
  NOR2_X2 U691 ( .A1(n697), .A2(n710), .ZN(n634) );
  NAND2_X1 U692 ( .A1(KEYINPUT2), .A2(n634), .ZN(n624) );
  NOR2_X1 U693 ( .A1(G953), .A2(n626), .ZN(n629) );
  XNOR2_X1 U694 ( .A(n627), .B(KEYINPUT119), .ZN(n628) );
  XNOR2_X1 U695 ( .A(n629), .B(n628), .ZN(G75) );
  XOR2_X1 U696 ( .A(KEYINPUT103), .B(KEYINPUT82), .Z(n631) );
  XNOR2_X1 U697 ( .A(KEYINPUT102), .B(KEYINPUT62), .ZN(n630) );
  XNOR2_X1 U698 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U699 ( .A(n633), .B(n632), .ZN(n638) );
  NAND2_X1 U700 ( .A1(G472), .A2(n349), .ZN(n637) );
  XNOR2_X1 U701 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U702 ( .A(n642), .B(n641), .ZN(G57) );
  XOR2_X1 U703 ( .A(G104), .B(KEYINPUT105), .Z(n644) );
  NAND2_X1 U704 ( .A1(n645), .A2(n659), .ZN(n643) );
  XNOR2_X1 U705 ( .A(n644), .B(n643), .ZN(G6) );
  XNOR2_X1 U706 ( .A(G107), .B(KEYINPUT27), .ZN(n649) );
  XOR2_X1 U707 ( .A(KEYINPUT106), .B(KEYINPUT26), .Z(n647) );
  NAND2_X1 U708 ( .A1(n645), .A2(n661), .ZN(n646) );
  XNOR2_X1 U709 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U710 ( .A(n649), .B(n648), .ZN(G9) );
  XNOR2_X1 U711 ( .A(n650), .B(G110), .ZN(n651) );
  XNOR2_X1 U712 ( .A(n651), .B(KEYINPUT107), .ZN(G12) );
  XOR2_X1 U713 ( .A(G128), .B(KEYINPUT29), .Z(n653) );
  NAND2_X1 U714 ( .A1(n655), .A2(n661), .ZN(n652) );
  XNOR2_X1 U715 ( .A(n653), .B(n652), .ZN(G30) );
  XOR2_X1 U716 ( .A(G143), .B(n654), .Z(G45) );
  XOR2_X1 U717 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n657) );
  NAND2_X1 U718 ( .A1(n655), .A2(n659), .ZN(n656) );
  XNOR2_X1 U719 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U720 ( .A(G146), .B(n658), .ZN(G48) );
  NAND2_X1 U721 ( .A1(n662), .A2(n659), .ZN(n660) );
  XNOR2_X1 U722 ( .A(n660), .B(G113), .ZN(G15) );
  NAND2_X1 U723 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U724 ( .A(n663), .B(KEYINPUT110), .ZN(n664) );
  XNOR2_X1 U725 ( .A(G116), .B(n664), .ZN(G18) );
  XOR2_X1 U726 ( .A(KEYINPUT37), .B(KEYINPUT111), .Z(n667) );
  XNOR2_X1 U727 ( .A(G125), .B(n665), .ZN(n666) );
  XNOR2_X1 U728 ( .A(n667), .B(n666), .ZN(G27) );
  XNOR2_X1 U729 ( .A(G140), .B(KEYINPUT112), .ZN(n669) );
  XNOR2_X1 U730 ( .A(n669), .B(n668), .ZN(G42) );
  XNOR2_X1 U731 ( .A(KEYINPUT55), .B(KEYINPUT80), .ZN(n672) );
  XNOR2_X1 U732 ( .A(n670), .B(KEYINPUT54), .ZN(n671) );
  XNOR2_X1 U733 ( .A(n672), .B(n671), .ZN(n674) );
  NAND2_X1 U734 ( .A1(n691), .A2(G210), .ZN(n673) );
  XOR2_X1 U735 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n677) );
  NAND2_X1 U736 ( .A1(n348), .A2(G469), .ZN(n676) );
  NOR2_X1 U737 ( .A1(n694), .A2(n679), .ZN(G54) );
  NAND2_X1 U738 ( .A1(n691), .A2(G475), .ZN(n684) );
  INV_X1 U739 ( .A(n680), .ZN(n682) );
  XOR2_X1 U740 ( .A(KEYINPUT59), .B(KEYINPUT65), .Z(n681) );
  XNOR2_X1 U741 ( .A(n684), .B(n683), .ZN(n685) );
  XOR2_X1 U742 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n687) );
  NAND2_X1 U743 ( .A1(n349), .A2(G478), .ZN(n686) );
  XNOR2_X1 U744 ( .A(n687), .B(n686), .ZN(n689) );
  XNOR2_X1 U745 ( .A(n689), .B(n688), .ZN(n690) );
  NOR2_X1 U746 ( .A1(n694), .A2(n690), .ZN(G63) );
  XNOR2_X1 U747 ( .A(n696), .B(KEYINPUT122), .ZN(G66) );
  NOR2_X1 U748 ( .A1(G953), .A2(n697), .ZN(n698) );
  XNOR2_X1 U749 ( .A(KEYINPUT123), .B(n698), .ZN(n702) );
  NAND2_X1 U750 ( .A1(G953), .A2(G224), .ZN(n699) );
  XNOR2_X1 U751 ( .A(KEYINPUT61), .B(n699), .ZN(n700) );
  NAND2_X1 U752 ( .A1(n700), .A2(G898), .ZN(n701) );
  NAND2_X1 U753 ( .A1(n702), .A2(n701), .ZN(n706) );
  NOR2_X1 U754 ( .A1(G898), .A2(n711), .ZN(n703) );
  NOR2_X1 U755 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U756 ( .A(n706), .B(n705), .ZN(n707) );
  XNOR2_X1 U757 ( .A(KEYINPUT124), .B(n707), .ZN(G69) );
  XOR2_X1 U758 ( .A(n709), .B(n708), .Z(n713) );
  XNOR2_X1 U759 ( .A(n713), .B(n710), .ZN(n712) );
  NAND2_X1 U760 ( .A1(n712), .A2(n711), .ZN(n718) );
  XNOR2_X1 U761 ( .A(G227), .B(n713), .ZN(n714) );
  NAND2_X1 U762 ( .A1(n714), .A2(G900), .ZN(n715) );
  XNOR2_X1 U763 ( .A(KEYINPUT126), .B(n715), .ZN(n716) );
  NAND2_X1 U764 ( .A1(n716), .A2(G953), .ZN(n717) );
  NAND2_X1 U765 ( .A1(n718), .A2(n717), .ZN(G72) );
  XOR2_X1 U766 ( .A(G137), .B(n719), .Z(G39) );
  XOR2_X1 U767 ( .A(G134), .B(n720), .Z(G36) );
  XNOR2_X1 U768 ( .A(n721), .B(G122), .ZN(n722) );
  XNOR2_X1 U769 ( .A(n722), .B(KEYINPUT127), .ZN(G24) );
  XOR2_X1 U770 ( .A(n723), .B(G101), .Z(G3) );
  XNOR2_X1 U771 ( .A(n724), .B(G119), .ZN(G21) );
  XOR2_X1 U772 ( .A(n725), .B(G131), .Z(G33) );
endmodule

