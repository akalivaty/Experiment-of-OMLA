

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U552 ( .A1(G2104), .A2(G2105), .ZN(n527) );
  INV_X1 U553 ( .A(G651), .ZN(n544) );
  NOR2_X1 U554 ( .A1(n731), .A2(n990), .ZN(n699) );
  NOR2_X1 U555 ( .A1(n737), .A2(n736), .ZN(n739) );
  INV_X2 U556 ( .A(G2105), .ZN(n522) );
  AND2_X1 U557 ( .A1(n694), .A2(n693), .ZN(n788) );
  NOR2_X2 U558 ( .A1(n653), .A2(n544), .ZN(n659) );
  NOR2_X1 U559 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U560 ( .A(n553), .B(KEYINPUT91), .ZN(n556) );
  BUF_X1 U561 ( .A(n618), .Z(n899) );
  XNOR2_X1 U562 ( .A(n527), .B(n526), .ZN(n618) );
  INV_X1 U563 ( .A(KEYINPUT17), .ZN(n526) );
  NOR2_X1 U564 ( .A1(n581), .A2(n580), .ZN(n583) );
  NOR2_X1 U565 ( .A1(G543), .A2(n544), .ZN(n538) );
  NOR2_X1 U566 ( .A1(G543), .A2(G651), .ZN(n542) );
  INV_X1 U567 ( .A(KEYINPUT66), .ZN(n528) );
  NAND2_X1 U568 ( .A1(n525), .A2(n518), .ZN(n535) );
  XNOR2_X2 U569 ( .A(n538), .B(n537), .ZN(n584) );
  XNOR2_X2 U570 ( .A(n529), .B(n528), .ZN(n558) );
  NAND2_X1 U571 ( .A1(n763), .A2(n762), .ZN(n516) );
  OR2_X1 U572 ( .A1(n521), .A2(n785), .ZN(n517) );
  XOR2_X1 U573 ( .A(n524), .B(n523), .Z(n518) );
  XOR2_X1 U574 ( .A(n562), .B(n561), .Z(n519) );
  AND2_X1 U575 ( .A1(n935), .A2(n830), .ZN(n520) );
  NAND2_X1 U576 ( .A1(G8), .A2(n743), .ZN(n521) );
  AND2_X1 U577 ( .A1(n731), .A2(G1341), .ZN(n696) );
  INV_X1 U578 ( .A(n731), .ZN(n712) );
  INV_X1 U579 ( .A(KEYINPUT29), .ZN(n722) );
  XNOR2_X1 U580 ( .A(KEYINPUT99), .B(KEYINPUT31), .ZN(n738) );
  INV_X1 U581 ( .A(n930), .ZN(n762) );
  NOR2_X1 U582 ( .A1(n712), .A2(n730), .ZN(n757) );
  INV_X1 U583 ( .A(KEYINPUT32), .ZN(n752) );
  NAND2_X2 U584 ( .A1(n788), .A2(n695), .ZN(n731) );
  BUF_X1 U585 ( .A(n731), .Z(n743) );
  NOR2_X1 U586 ( .A1(n767), .A2(n521), .ZN(n774) );
  INV_X1 U587 ( .A(KEYINPUT1), .ZN(n536) );
  INV_X1 U588 ( .A(KEYINPUT104), .ZN(n782) );
  XNOR2_X1 U589 ( .A(n536), .B(KEYINPUT68), .ZN(n537) );
  NAND2_X1 U590 ( .A1(n618), .A2(G138), .ZN(n553) );
  NOR2_X1 U591 ( .A1(n818), .A2(n520), .ZN(n819) );
  XNOR2_X1 U592 ( .A(n595), .B(KEYINPUT15), .ZN(n697) );
  NOR2_X2 U593 ( .A1(G2104), .A2(n522), .ZN(n904) );
  BUF_X1 U594 ( .A(n697), .Z(n933) );
  INV_X1 U595 ( .A(KEYINPUT67), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n533), .B(n532), .ZN(n534) );
  NOR2_X2 U597 ( .A1(n535), .A2(n534), .ZN(G160) );
  NAND2_X1 U598 ( .A1(G125), .A2(n904), .ZN(n525) );
  XOR2_X1 U599 ( .A(KEYINPUT23), .B(KEYINPUT65), .Z(n524) );
  AND2_X4 U600 ( .A1(n522), .A2(G2104), .ZN(n615) );
  NAND2_X1 U601 ( .A1(G101), .A2(n615), .ZN(n523) );
  NAND2_X1 U602 ( .A1(n618), .A2(G137), .ZN(n531) );
  NAND2_X1 U603 ( .A1(G2104), .A2(G2105), .ZN(n529) );
  NAND2_X1 U604 ( .A1(n558), .A2(G113), .ZN(n530) );
  NAND2_X1 U605 ( .A1(n531), .A2(n530), .ZN(n533) );
  XOR2_X1 U606 ( .A(KEYINPUT0), .B(G543), .Z(n653) );
  NOR2_X2 U607 ( .A1(G651), .A2(n653), .ZN(n663) );
  NAND2_X1 U608 ( .A1(n663), .A2(G51), .ZN(n540) );
  NAND2_X1 U609 ( .A1(G63), .A2(n584), .ZN(n539) );
  NAND2_X1 U610 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U611 ( .A(KEYINPUT6), .B(n541), .ZN(n549) );
  XNOR2_X2 U612 ( .A(n542), .B(KEYINPUT64), .ZN(n656) );
  NAND2_X1 U613 ( .A1(G89), .A2(n656), .ZN(n543) );
  XNOR2_X1 U614 ( .A(n543), .B(KEYINPUT4), .ZN(n546) );
  NAND2_X1 U615 ( .A1(G76), .A2(n659), .ZN(n545) );
  NAND2_X1 U616 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U617 ( .A(n547), .B(KEYINPUT5), .Z(n548) );
  NOR2_X1 U618 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U619 ( .A(KEYINPUT7), .B(n550), .Z(n552) );
  XOR2_X1 U620 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n551) );
  XNOR2_X1 U621 ( .A(n552), .B(n551), .ZN(G168) );
  XOR2_X1 U622 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U623 ( .A1(n615), .A2(G102), .ZN(n554) );
  XOR2_X1 U624 ( .A(KEYINPUT90), .B(n554), .Z(n555) );
  XNOR2_X1 U625 ( .A(n557), .B(KEYINPUT92), .ZN(n563) );
  NAND2_X1 U626 ( .A1(G126), .A2(n904), .ZN(n560) );
  NAND2_X1 U627 ( .A1(G114), .A2(n558), .ZN(n559) );
  NAND2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n562) );
  INV_X1 U629 ( .A(KEYINPUT89), .ZN(n561) );
  NAND2_X1 U630 ( .A1(n563), .A2(n519), .ZN(n694) );
  INV_X1 U631 ( .A(n694), .ZN(G164) );
  NAND2_X1 U632 ( .A1(n663), .A2(G52), .ZN(n565) );
  NAND2_X1 U633 ( .A1(G64), .A2(n584), .ZN(n564) );
  NAND2_X1 U634 ( .A1(n565), .A2(n564), .ZN(n570) );
  NAND2_X1 U635 ( .A1(n659), .A2(G77), .ZN(n567) );
  NAND2_X1 U636 ( .A1(G90), .A2(n656), .ZN(n566) );
  NAND2_X1 U637 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U638 ( .A(KEYINPUT9), .B(n568), .Z(n569) );
  NOR2_X1 U639 ( .A1(n570), .A2(n569), .ZN(G171) );
  AND2_X1 U640 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U641 ( .A(G57), .ZN(G237) );
  INV_X1 U642 ( .A(G132), .ZN(G219) );
  INV_X1 U643 ( .A(G82), .ZN(G220) );
  NAND2_X1 U644 ( .A1(G7), .A2(G661), .ZN(n571) );
  XNOR2_X1 U645 ( .A(n571), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U646 ( .A(G223), .ZN(n846) );
  NAND2_X1 U647 ( .A1(n846), .A2(G567), .ZN(n572) );
  XOR2_X1 U648 ( .A(KEYINPUT11), .B(n572), .Z(G234) );
  XOR2_X1 U649 ( .A(KEYINPUT72), .B(KEYINPUT14), .Z(n574) );
  NAND2_X1 U650 ( .A1(G56), .A2(n584), .ZN(n573) );
  XNOR2_X1 U651 ( .A(n574), .B(n573), .ZN(n581) );
  XNOR2_X1 U652 ( .A(KEYINPUT13), .B(KEYINPUT73), .ZN(n579) );
  NAND2_X1 U653 ( .A1(G81), .A2(n656), .ZN(n575) );
  XNOR2_X1 U654 ( .A(n575), .B(KEYINPUT12), .ZN(n577) );
  NAND2_X1 U655 ( .A1(G68), .A2(n659), .ZN(n576) );
  NAND2_X1 U656 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U657 ( .A(n579), .B(n578), .ZN(n580) );
  NAND2_X1 U658 ( .A1(n663), .A2(G43), .ZN(n582) );
  NAND2_X1 U659 ( .A1(n583), .A2(n582), .ZN(n937) );
  INV_X1 U660 ( .A(G860), .ZN(n608) );
  OR2_X1 U661 ( .A1(n937), .A2(n608), .ZN(G153) );
  INV_X1 U662 ( .A(G171), .ZN(G301) );
  NAND2_X1 U663 ( .A1(G868), .A2(G301), .ZN(n597) );
  NAND2_X1 U664 ( .A1(G66), .A2(n584), .ZN(n585) );
  XNOR2_X1 U665 ( .A(n585), .B(KEYINPUT74), .ZN(n587) );
  NAND2_X1 U666 ( .A1(G92), .A2(n656), .ZN(n586) );
  NAND2_X1 U667 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U668 ( .A(n588), .B(KEYINPUT75), .ZN(n594) );
  NAND2_X1 U669 ( .A1(G79), .A2(n659), .ZN(n589) );
  XOR2_X1 U670 ( .A(KEYINPUT76), .B(n589), .Z(n592) );
  NAND2_X1 U671 ( .A1(G54), .A2(n663), .ZN(n590) );
  XNOR2_X1 U672 ( .A(KEYINPUT77), .B(n590), .ZN(n591) );
  NOR2_X1 U673 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U674 ( .A1(n594), .A2(n593), .ZN(n595) );
  OR2_X1 U675 ( .A1(n933), .A2(G868), .ZN(n596) );
  NAND2_X1 U676 ( .A1(n597), .A2(n596), .ZN(G284) );
  NAND2_X1 U677 ( .A1(n584), .A2(G65), .ZN(n598) );
  XNOR2_X1 U678 ( .A(n598), .B(KEYINPUT70), .ZN(n601) );
  NAND2_X1 U679 ( .A1(n656), .A2(G91), .ZN(n599) );
  XOR2_X1 U680 ( .A(KEYINPUT69), .B(n599), .Z(n600) );
  NAND2_X1 U681 ( .A1(n601), .A2(n600), .ZN(n605) );
  NAND2_X1 U682 ( .A1(G78), .A2(n659), .ZN(n603) );
  NAND2_X1 U683 ( .A1(G53), .A2(n663), .ZN(n602) );
  NAND2_X1 U684 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U685 ( .A1(n605), .A2(n604), .ZN(n927) );
  XNOR2_X1 U686 ( .A(n927), .B(KEYINPUT71), .ZN(G299) );
  NAND2_X1 U687 ( .A1(G868), .A2(G286), .ZN(n607) );
  INV_X1 U688 ( .A(G868), .ZN(n674) );
  NAND2_X1 U689 ( .A1(n674), .A2(G299), .ZN(n606) );
  NAND2_X1 U690 ( .A1(n607), .A2(n606), .ZN(G297) );
  NAND2_X1 U691 ( .A1(n608), .A2(G559), .ZN(n609) );
  NAND2_X1 U692 ( .A1(n609), .A2(n933), .ZN(n610) );
  XNOR2_X1 U693 ( .A(n610), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U694 ( .A1(G868), .A2(n937), .ZN(n613) );
  NAND2_X1 U695 ( .A1(G868), .A2(n933), .ZN(n611) );
  NOR2_X1 U696 ( .A1(G559), .A2(n611), .ZN(n612) );
  NOR2_X1 U697 ( .A1(n613), .A2(n612), .ZN(G282) );
  NAND2_X1 U698 ( .A1(n904), .A2(G123), .ZN(n614) );
  XNOR2_X1 U699 ( .A(n614), .B(KEYINPUT18), .ZN(n617) );
  NAND2_X1 U700 ( .A1(G99), .A2(n615), .ZN(n616) );
  NAND2_X1 U701 ( .A1(n617), .A2(n616), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n899), .A2(G135), .ZN(n620) );
  NAND2_X1 U703 ( .A1(G111), .A2(n558), .ZN(n619) );
  NAND2_X1 U704 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U705 ( .A1(n622), .A2(n621), .ZN(n1014) );
  XOR2_X1 U706 ( .A(n1014), .B(G2096), .Z(n623) );
  NOR2_X1 U707 ( .A1(G2100), .A2(n623), .ZN(n624) );
  XOR2_X1 U708 ( .A(KEYINPUT80), .B(n624), .Z(G156) );
  XNOR2_X1 U709 ( .A(n937), .B(KEYINPUT81), .ZN(n626) );
  NAND2_X1 U710 ( .A1(n933), .A2(G559), .ZN(n625) );
  XOR2_X1 U711 ( .A(n626), .B(n625), .Z(n671) );
  NOR2_X1 U712 ( .A1(n671), .A2(G860), .ZN(n635) );
  NAND2_X1 U713 ( .A1(n659), .A2(G80), .ZN(n628) );
  NAND2_X1 U714 ( .A1(G67), .A2(n584), .ZN(n627) );
  NAND2_X1 U715 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U716 ( .A1(G93), .A2(n656), .ZN(n629) );
  XNOR2_X1 U717 ( .A(KEYINPUT83), .B(n629), .ZN(n630) );
  NOR2_X1 U718 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U719 ( .A1(n663), .A2(G55), .ZN(n632) );
  NAND2_X1 U720 ( .A1(n633), .A2(n632), .ZN(n673) );
  XOR2_X1 U721 ( .A(n673), .B(KEYINPUT82), .Z(n634) );
  XNOR2_X1 U722 ( .A(n635), .B(n634), .ZN(G145) );
  AND2_X1 U723 ( .A1(G60), .A2(n584), .ZN(n639) );
  NAND2_X1 U724 ( .A1(n659), .A2(G72), .ZN(n637) );
  NAND2_X1 U725 ( .A1(G85), .A2(n656), .ZN(n636) );
  NAND2_X1 U726 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U727 ( .A1(n639), .A2(n638), .ZN(n641) );
  NAND2_X1 U728 ( .A1(n663), .A2(G47), .ZN(n640) );
  NAND2_X1 U729 ( .A1(n641), .A2(n640), .ZN(G290) );
  NAND2_X1 U730 ( .A1(n659), .A2(G75), .ZN(n643) );
  NAND2_X1 U731 ( .A1(G88), .A2(n656), .ZN(n642) );
  NAND2_X1 U732 ( .A1(n643), .A2(n642), .ZN(n647) );
  NAND2_X1 U733 ( .A1(n663), .A2(G50), .ZN(n645) );
  NAND2_X1 U734 ( .A1(G62), .A2(n584), .ZN(n644) );
  NAND2_X1 U735 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U736 ( .A1(n647), .A2(n646), .ZN(G166) );
  NAND2_X1 U737 ( .A1(G651), .A2(G74), .ZN(n648) );
  XNOR2_X1 U738 ( .A(n648), .B(KEYINPUT84), .ZN(n650) );
  NAND2_X1 U739 ( .A1(G49), .A2(n663), .ZN(n649) );
  NAND2_X1 U740 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U741 ( .A(KEYINPUT85), .B(n651), .Z(n652) );
  NOR2_X1 U742 ( .A1(n584), .A2(n652), .ZN(n655) );
  NAND2_X1 U743 ( .A1(n653), .A2(G87), .ZN(n654) );
  NAND2_X1 U744 ( .A1(n655), .A2(n654), .ZN(G288) );
  NAND2_X1 U745 ( .A1(G61), .A2(n584), .ZN(n658) );
  NAND2_X1 U746 ( .A1(G86), .A2(n656), .ZN(n657) );
  NAND2_X1 U747 ( .A1(n658), .A2(n657), .ZN(n662) );
  NAND2_X1 U748 ( .A1(n659), .A2(G73), .ZN(n660) );
  XOR2_X1 U749 ( .A(KEYINPUT2), .B(n660), .Z(n661) );
  NOR2_X1 U750 ( .A1(n662), .A2(n661), .ZN(n665) );
  NAND2_X1 U751 ( .A1(n663), .A2(G48), .ZN(n664) );
  NAND2_X1 U752 ( .A1(n665), .A2(n664), .ZN(G305) );
  XNOR2_X1 U753 ( .A(KEYINPUT19), .B(G290), .ZN(n670) );
  XOR2_X1 U754 ( .A(G288), .B(G299), .Z(n666) );
  XNOR2_X1 U755 ( .A(n673), .B(n666), .ZN(n667) );
  XNOR2_X1 U756 ( .A(G166), .B(n667), .ZN(n668) );
  XNOR2_X1 U757 ( .A(n668), .B(G305), .ZN(n669) );
  XNOR2_X1 U758 ( .A(n670), .B(n669), .ZN(n915) );
  XOR2_X1 U759 ( .A(n671), .B(n915), .Z(n672) );
  NAND2_X1 U760 ( .A1(n672), .A2(G868), .ZN(n676) );
  NAND2_X1 U761 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U762 ( .A1(n676), .A2(n675), .ZN(G295) );
  NAND2_X1 U763 ( .A1(G2078), .A2(G2084), .ZN(n677) );
  XOR2_X1 U764 ( .A(KEYINPUT20), .B(n677), .Z(n678) );
  NAND2_X1 U765 ( .A1(G2090), .A2(n678), .ZN(n679) );
  XNOR2_X1 U766 ( .A(n679), .B(KEYINPUT87), .ZN(n681) );
  XOR2_X1 U767 ( .A(KEYINPUT21), .B(KEYINPUT86), .Z(n680) );
  XNOR2_X1 U768 ( .A(n681), .B(n680), .ZN(n682) );
  NAND2_X1 U769 ( .A1(n682), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U770 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U771 ( .A1(G220), .A2(G219), .ZN(n683) );
  XOR2_X1 U772 ( .A(KEYINPUT22), .B(n683), .Z(n684) );
  NOR2_X1 U773 ( .A1(G218), .A2(n684), .ZN(n685) );
  NAND2_X1 U774 ( .A1(G96), .A2(n685), .ZN(n853) );
  AND2_X1 U775 ( .A1(G2106), .A2(n853), .ZN(n690) );
  NAND2_X1 U776 ( .A1(G108), .A2(G120), .ZN(n686) );
  NOR2_X1 U777 ( .A1(G237), .A2(n686), .ZN(n687) );
  NAND2_X1 U778 ( .A1(G69), .A2(n687), .ZN(n852) );
  NAND2_X1 U779 ( .A1(G567), .A2(n852), .ZN(n688) );
  XOR2_X1 U780 ( .A(KEYINPUT88), .B(n688), .Z(n689) );
  NOR2_X1 U781 ( .A1(n690), .A2(n689), .ZN(G319) );
  INV_X1 U782 ( .A(G319), .ZN(n692) );
  NAND2_X1 U783 ( .A1(G661), .A2(G483), .ZN(n691) );
  NOR2_X1 U784 ( .A1(n692), .A2(n691), .ZN(n851) );
  NAND2_X1 U785 ( .A1(n851), .A2(G36), .ZN(G176) );
  XNOR2_X1 U786 ( .A(KEYINPUT93), .B(G166), .ZN(G303) );
  INV_X1 U787 ( .A(G1384), .ZN(n693) );
  NAND2_X1 U788 ( .A1(G160), .A2(G40), .ZN(n787) );
  INV_X1 U789 ( .A(n787), .ZN(n695) );
  NOR2_X1 U790 ( .A1(n696), .A2(n937), .ZN(n706) );
  AND2_X1 U791 ( .A1(n706), .A2(n697), .ZN(n700) );
  INV_X1 U792 ( .A(G1996), .ZN(n990) );
  INV_X1 U793 ( .A(KEYINPUT26), .ZN(n698) );
  XNOR2_X1 U794 ( .A(n699), .B(n698), .ZN(n707) );
  NAND2_X1 U795 ( .A1(n700), .A2(n707), .ZN(n704) );
  NOR2_X1 U796 ( .A1(n712), .A2(G1348), .ZN(n702) );
  NOR2_X1 U797 ( .A1(G2067), .A2(n743), .ZN(n701) );
  NOR2_X1 U798 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U799 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U800 ( .A(n705), .B(KEYINPUT98), .ZN(n710) );
  AND2_X1 U801 ( .A1(n707), .A2(n706), .ZN(n708) );
  OR2_X1 U802 ( .A1(n708), .A2(n933), .ZN(n709) );
  NAND2_X1 U803 ( .A1(n710), .A2(n709), .ZN(n716) );
  NAND2_X1 U804 ( .A1(n712), .A2(G2072), .ZN(n711) );
  XNOR2_X1 U805 ( .A(n711), .B(KEYINPUT27), .ZN(n714) );
  INV_X1 U806 ( .A(G1956), .ZN(n955) );
  NOR2_X1 U807 ( .A1(n955), .A2(n712), .ZN(n713) );
  NOR2_X1 U808 ( .A1(n714), .A2(n713), .ZN(n717) );
  NAND2_X1 U809 ( .A1(n927), .A2(n717), .ZN(n715) );
  NAND2_X1 U810 ( .A1(n716), .A2(n715), .ZN(n721) );
  NOR2_X1 U811 ( .A1(n717), .A2(n927), .ZN(n719) );
  INV_X1 U812 ( .A(KEYINPUT28), .ZN(n718) );
  XNOR2_X1 U813 ( .A(n719), .B(n718), .ZN(n720) );
  NAND2_X1 U814 ( .A1(n721), .A2(n720), .ZN(n723) );
  XNOR2_X1 U815 ( .A(n723), .B(n722), .ZN(n728) );
  XNOR2_X1 U816 ( .A(G2078), .B(KEYINPUT25), .ZN(n989) );
  NOR2_X1 U817 ( .A1(n743), .A2(n989), .ZN(n725) );
  AND2_X1 U818 ( .A1(n743), .A2(G1961), .ZN(n724) );
  NOR2_X1 U819 ( .A1(n725), .A2(n724), .ZN(n735) );
  AND2_X1 U820 ( .A1(G171), .A2(n735), .ZN(n726) );
  XNOR2_X1 U821 ( .A(n726), .B(KEYINPUT97), .ZN(n727) );
  NAND2_X1 U822 ( .A1(n728), .A2(n727), .ZN(n741) );
  INV_X1 U823 ( .A(G8), .ZN(n729) );
  OR2_X1 U824 ( .A1(n729), .A2(G1966), .ZN(n730) );
  NOR2_X1 U825 ( .A1(G2084), .A2(n731), .ZN(n755) );
  NOR2_X1 U826 ( .A1(n757), .A2(n755), .ZN(n732) );
  NAND2_X1 U827 ( .A1(n732), .A2(G8), .ZN(n733) );
  XNOR2_X1 U828 ( .A(KEYINPUT30), .B(n733), .ZN(n734) );
  NOR2_X1 U829 ( .A1(n734), .A2(G168), .ZN(n737) );
  NOR2_X1 U830 ( .A1(G171), .A2(n735), .ZN(n736) );
  XNOR2_X1 U831 ( .A(n739), .B(n738), .ZN(n740) );
  NAND2_X1 U832 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U833 ( .A(n742), .B(KEYINPUT100), .ZN(n754) );
  NAND2_X1 U834 ( .A1(n754), .A2(G286), .ZN(n748) );
  NOR2_X1 U835 ( .A1(G1971), .A2(n521), .ZN(n745) );
  NOR2_X1 U836 ( .A1(G2090), .A2(n743), .ZN(n744) );
  NOR2_X1 U837 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U838 ( .A1(n746), .A2(G303), .ZN(n747) );
  NAND2_X1 U839 ( .A1(n748), .A2(n747), .ZN(n750) );
  INV_X1 U840 ( .A(KEYINPUT101), .ZN(n749) );
  XNOR2_X1 U841 ( .A(n750), .B(n749), .ZN(n751) );
  NAND2_X1 U842 ( .A1(n751), .A2(G8), .ZN(n753) );
  XNOR2_X1 U843 ( .A(n753), .B(n752), .ZN(n760) );
  NAND2_X1 U844 ( .A1(G8), .A2(n755), .ZN(n756) );
  NAND2_X1 U845 ( .A1(n754), .A2(n756), .ZN(n758) );
  NOR2_X1 U846 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X2 U847 ( .A1(n760), .A2(n759), .ZN(n768) );
  NOR2_X1 U848 ( .A1(G1971), .A2(G303), .ZN(n761) );
  XOR2_X1 U849 ( .A(n761), .B(KEYINPUT102), .Z(n763) );
  NOR2_X1 U850 ( .A1(G1976), .A2(G288), .ZN(n930) );
  OR2_X1 U851 ( .A1(n768), .A2(n516), .ZN(n764) );
  NAND2_X1 U852 ( .A1(G1976), .A2(G288), .ZN(n934) );
  NAND2_X1 U853 ( .A1(n764), .A2(n934), .ZN(n766) );
  INV_X1 U854 ( .A(KEYINPUT103), .ZN(n765) );
  XNOR2_X1 U855 ( .A(n766), .B(n765), .ZN(n767) );
  INV_X1 U856 ( .A(n768), .ZN(n771) );
  NOR2_X1 U857 ( .A1(G2090), .A2(G303), .ZN(n769) );
  NAND2_X1 U858 ( .A1(G8), .A2(n769), .ZN(n770) );
  NAND2_X1 U859 ( .A1(n771), .A2(n770), .ZN(n772) );
  AND2_X1 U860 ( .A1(n772), .A2(n521), .ZN(n779) );
  OR2_X1 U861 ( .A1(KEYINPUT33), .A2(n779), .ZN(n773) );
  NOR2_X1 U862 ( .A1(n774), .A2(n773), .ZN(n781) );
  NAND2_X1 U863 ( .A1(n930), .A2(KEYINPUT33), .ZN(n775) );
  NOR2_X1 U864 ( .A1(n775), .A2(n521), .ZN(n777) );
  XOR2_X1 U865 ( .A(G1981), .B(G305), .Z(n944) );
  INV_X1 U866 ( .A(n944), .ZN(n776) );
  NOR2_X1 U867 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U868 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n783) );
  XNOR2_X1 U870 ( .A(n783), .B(n782), .ZN(n786) );
  NOR2_X1 U871 ( .A1(G1981), .A2(G305), .ZN(n784) );
  XOR2_X1 U872 ( .A(n784), .B(KEYINPUT24), .Z(n785) );
  NAND2_X1 U873 ( .A1(n786), .A2(n517), .ZN(n820) );
  NOR2_X1 U874 ( .A1(n788), .A2(n787), .ZN(n830) );
  XOR2_X1 U875 ( .A(KEYINPUT96), .B(KEYINPUT36), .Z(n800) );
  NAND2_X1 U876 ( .A1(G128), .A2(n904), .ZN(n790) );
  NAND2_X1 U877 ( .A1(G116), .A2(n558), .ZN(n789) );
  NAND2_X1 U878 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U879 ( .A(KEYINPUT35), .B(n791), .Z(n798) );
  XNOR2_X1 U880 ( .A(KEYINPUT94), .B(KEYINPUT95), .ZN(n795) );
  NAND2_X1 U881 ( .A1(G104), .A2(n615), .ZN(n793) );
  NAND2_X1 U882 ( .A1(G140), .A2(n899), .ZN(n792) );
  NAND2_X1 U883 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U884 ( .A(n795), .B(n794), .ZN(n796) );
  XOR2_X1 U885 ( .A(n796), .B(KEYINPUT34), .Z(n797) );
  NOR2_X1 U886 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U887 ( .A(n800), .B(n799), .Z(n883) );
  XNOR2_X1 U888 ( .A(KEYINPUT37), .B(G2067), .ZN(n828) );
  NOR2_X1 U889 ( .A1(n883), .A2(n828), .ZN(n1013) );
  NAND2_X1 U890 ( .A1(n830), .A2(n1013), .ZN(n826) );
  NAND2_X1 U891 ( .A1(G119), .A2(n904), .ZN(n802) );
  NAND2_X1 U892 ( .A1(G131), .A2(n899), .ZN(n801) );
  NAND2_X1 U893 ( .A1(n802), .A2(n801), .ZN(n806) );
  NAND2_X1 U894 ( .A1(n615), .A2(G95), .ZN(n804) );
  NAND2_X1 U895 ( .A1(G107), .A2(n558), .ZN(n803) );
  NAND2_X1 U896 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U897 ( .A1(n806), .A2(n805), .ZN(n882) );
  INV_X1 U898 ( .A(G1991), .ZN(n872) );
  NOR2_X1 U899 ( .A1(n882), .A2(n872), .ZN(n815) );
  NAND2_X1 U900 ( .A1(G129), .A2(n904), .ZN(n808) );
  NAND2_X1 U901 ( .A1(G141), .A2(n899), .ZN(n807) );
  NAND2_X1 U902 ( .A1(n808), .A2(n807), .ZN(n811) );
  NAND2_X1 U903 ( .A1(n615), .A2(G105), .ZN(n809) );
  XOR2_X1 U904 ( .A(KEYINPUT38), .B(n809), .Z(n810) );
  NOR2_X1 U905 ( .A1(n811), .A2(n810), .ZN(n813) );
  NAND2_X1 U906 ( .A1(G117), .A2(n558), .ZN(n812) );
  NAND2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n881) );
  AND2_X1 U908 ( .A1(G1996), .A2(n881), .ZN(n814) );
  NOR2_X1 U909 ( .A1(n815), .A2(n814), .ZN(n1007) );
  INV_X1 U910 ( .A(n830), .ZN(n816) );
  NOR2_X1 U911 ( .A1(n1007), .A2(n816), .ZN(n823) );
  INV_X1 U912 ( .A(n823), .ZN(n817) );
  NAND2_X1 U913 ( .A1(n826), .A2(n817), .ZN(n818) );
  XNOR2_X1 U914 ( .A(G1986), .B(G290), .ZN(n935) );
  NAND2_X1 U915 ( .A1(n820), .A2(n819), .ZN(n833) );
  NOR2_X1 U916 ( .A1(G1996), .A2(n881), .ZN(n1010) );
  NOR2_X1 U917 ( .A1(G1986), .A2(G290), .ZN(n821) );
  AND2_X1 U918 ( .A1(n872), .A2(n882), .ZN(n1015) );
  NOR2_X1 U919 ( .A1(n821), .A2(n1015), .ZN(n822) );
  NOR2_X1 U920 ( .A1(n823), .A2(n822), .ZN(n824) );
  NOR2_X1 U921 ( .A1(n1010), .A2(n824), .ZN(n825) );
  XNOR2_X1 U922 ( .A(n825), .B(KEYINPUT39), .ZN(n827) );
  NAND2_X1 U923 ( .A1(n827), .A2(n826), .ZN(n829) );
  NAND2_X1 U924 ( .A1(n883), .A2(n828), .ZN(n1018) );
  NAND2_X1 U925 ( .A1(n829), .A2(n1018), .ZN(n831) );
  NAND2_X1 U926 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U927 ( .A1(n833), .A2(n832), .ZN(n835) );
  XOR2_X1 U928 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n834) );
  XNOR2_X1 U929 ( .A(n835), .B(n834), .ZN(G329) );
  XNOR2_X1 U930 ( .A(G2454), .B(G2446), .ZN(n844) );
  XNOR2_X1 U931 ( .A(G2430), .B(G2443), .ZN(n842) );
  XOR2_X1 U932 ( .A(G2435), .B(KEYINPUT106), .Z(n837) );
  XNOR2_X1 U933 ( .A(G2451), .B(G2438), .ZN(n836) );
  XNOR2_X1 U934 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U935 ( .A(n838), .B(G2427), .Z(n840) );
  XNOR2_X1 U936 ( .A(G1341), .B(G1348), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n842), .B(n841), .ZN(n843) );
  XNOR2_X1 U939 ( .A(n844), .B(n843), .ZN(n845) );
  NAND2_X1 U940 ( .A1(n845), .A2(G14), .ZN(n922) );
  XNOR2_X1 U941 ( .A(KEYINPUT107), .B(n922), .ZN(G401) );
  NAND2_X1 U942 ( .A1(G2106), .A2(n846), .ZN(G217) );
  INV_X1 U943 ( .A(G661), .ZN(n848) );
  NAND2_X1 U944 ( .A1(G2), .A2(G15), .ZN(n847) );
  NOR2_X1 U945 ( .A1(n848), .A2(n847), .ZN(n849) );
  XOR2_X1 U946 ( .A(KEYINPUT108), .B(n849), .Z(G259) );
  NAND2_X1 U947 ( .A1(G3), .A2(G1), .ZN(n850) );
  NAND2_X1 U948 ( .A1(n851), .A2(n850), .ZN(G188) );
  XNOR2_X1 U949 ( .A(G120), .B(KEYINPUT109), .ZN(G236) );
  INV_X1 U951 ( .A(G108), .ZN(G238) );
  INV_X1 U952 ( .A(G96), .ZN(G221) );
  NOR2_X1 U953 ( .A1(n853), .A2(n852), .ZN(G325) );
  INV_X1 U954 ( .A(G325), .ZN(G261) );
  XOR2_X1 U955 ( .A(G2096), .B(KEYINPUT43), .Z(n855) );
  XNOR2_X1 U956 ( .A(G2090), .B(G2678), .ZN(n854) );
  XNOR2_X1 U957 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U958 ( .A(n856), .B(KEYINPUT110), .Z(n858) );
  XNOR2_X1 U959 ( .A(G2067), .B(G2072), .ZN(n857) );
  XNOR2_X1 U960 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U961 ( .A(KEYINPUT42), .B(G2100), .Z(n860) );
  XNOR2_X1 U962 ( .A(G2078), .B(G2084), .ZN(n859) );
  XNOR2_X1 U963 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U964 ( .A(n862), .B(n861), .ZN(G227) );
  XOR2_X1 U965 ( .A(G1971), .B(G1961), .Z(n864) );
  XNOR2_X1 U966 ( .A(G1996), .B(G1956), .ZN(n863) );
  XNOR2_X1 U967 ( .A(n864), .B(n863), .ZN(n868) );
  XOR2_X1 U968 ( .A(G1976), .B(G1966), .Z(n866) );
  XNOR2_X1 U969 ( .A(G1986), .B(G1981), .ZN(n865) );
  XNOR2_X1 U970 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U971 ( .A(n868), .B(n867), .Z(n870) );
  XNOR2_X1 U972 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n869) );
  XNOR2_X1 U973 ( .A(n870), .B(n869), .ZN(n871) );
  XNOR2_X1 U974 ( .A(G2474), .B(n871), .ZN(n873) );
  XNOR2_X1 U975 ( .A(n873), .B(n872), .ZN(G229) );
  NAND2_X1 U976 ( .A1(n904), .A2(G124), .ZN(n874) );
  XNOR2_X1 U977 ( .A(n874), .B(KEYINPUT44), .ZN(n876) );
  NAND2_X1 U978 ( .A1(G100), .A2(n615), .ZN(n875) );
  NAND2_X1 U979 ( .A1(n876), .A2(n875), .ZN(n880) );
  NAND2_X1 U980 ( .A1(n899), .A2(G136), .ZN(n878) );
  NAND2_X1 U981 ( .A1(G112), .A2(n558), .ZN(n877) );
  NAND2_X1 U982 ( .A1(n878), .A2(n877), .ZN(n879) );
  NOR2_X1 U983 ( .A1(n880), .A2(n879), .ZN(G162) );
  XNOR2_X1 U984 ( .A(n882), .B(n881), .ZN(n885) );
  XNOR2_X1 U985 ( .A(G160), .B(n883), .ZN(n884) );
  XNOR2_X1 U986 ( .A(n885), .B(n884), .ZN(n898) );
  XOR2_X1 U987 ( .A(KEYINPUT112), .B(KEYINPUT46), .Z(n887) );
  XNOR2_X1 U988 ( .A(G162), .B(KEYINPUT48), .ZN(n886) );
  XNOR2_X1 U989 ( .A(n887), .B(n886), .ZN(n896) );
  NAND2_X1 U990 ( .A1(G130), .A2(n904), .ZN(n889) );
  NAND2_X1 U991 ( .A1(G118), .A2(n558), .ZN(n888) );
  NAND2_X1 U992 ( .A1(n889), .A2(n888), .ZN(n894) );
  NAND2_X1 U993 ( .A1(G106), .A2(n615), .ZN(n891) );
  NAND2_X1 U994 ( .A1(G142), .A2(n899), .ZN(n890) );
  NAND2_X1 U995 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U996 ( .A(n892), .B(KEYINPUT45), .Z(n893) );
  NOR2_X1 U997 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U998 ( .A(n896), .B(n895), .Z(n897) );
  XOR2_X1 U999 ( .A(n898), .B(n897), .Z(n912) );
  NAND2_X1 U1000 ( .A1(G103), .A2(n615), .ZN(n901) );
  NAND2_X1 U1001 ( .A1(G139), .A2(n899), .ZN(n900) );
  NAND2_X1 U1002 ( .A1(n901), .A2(n900), .ZN(n902) );
  XOR2_X1 U1003 ( .A(KEYINPUT113), .B(n902), .Z(n910) );
  NAND2_X1 U1004 ( .A1(G115), .A2(n558), .ZN(n903) );
  XNOR2_X1 U1005 ( .A(KEYINPUT115), .B(n903), .ZN(n907) );
  NAND2_X1 U1006 ( .A1(n904), .A2(G127), .ZN(n905) );
  XOR2_X1 U1007 ( .A(KEYINPUT114), .B(n905), .Z(n906) );
  NOR2_X1 U1008 ( .A1(n907), .A2(n906), .ZN(n908) );
  XNOR2_X1 U1009 ( .A(n908), .B(KEYINPUT47), .ZN(n909) );
  NOR2_X1 U1010 ( .A1(n910), .A2(n909), .ZN(n1019) );
  XNOR2_X1 U1011 ( .A(n1019), .B(n1014), .ZN(n911) );
  XNOR2_X1 U1012 ( .A(n912), .B(n911), .ZN(n913) );
  XNOR2_X1 U1013 ( .A(n913), .B(G164), .ZN(n914) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n914), .ZN(G395) );
  XNOR2_X1 U1015 ( .A(n933), .B(G286), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(G171), .B(n915), .ZN(n916) );
  XNOR2_X1 U1017 ( .A(n916), .B(n937), .ZN(n917) );
  XNOR2_X1 U1018 ( .A(n918), .B(n917), .ZN(n919) );
  NOR2_X1 U1019 ( .A1(G37), .A2(n919), .ZN(G397) );
  NOR2_X1 U1020 ( .A1(G227), .A2(G229), .ZN(n921) );
  XNOR2_X1 U1021 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n920) );
  XNOR2_X1 U1022 ( .A(n921), .B(n920), .ZN(n924) );
  NAND2_X1 U1023 ( .A1(G319), .A2(n922), .ZN(n923) );
  NOR2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n926) );
  NOR2_X1 U1025 ( .A1(G395), .A2(G397), .ZN(n925) );
  NAND2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(G225) );
  INV_X1 U1027 ( .A(G225), .ZN(G308) );
  INV_X1 U1028 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1029 ( .A(G16), .B(KEYINPUT56), .ZN(n952) );
  XNOR2_X1 U1030 ( .A(G171), .B(G1961), .ZN(n929) );
  XNOR2_X1 U1031 ( .A(n927), .B(G1956), .ZN(n928) );
  NAND2_X1 U1032 ( .A1(n929), .A2(n928), .ZN(n932) );
  XNOR2_X1 U1033 ( .A(KEYINPUT124), .B(n930), .ZN(n931) );
  NOR2_X1 U1034 ( .A1(n932), .A2(n931), .ZN(n950) );
  XNOR2_X1 U1035 ( .A(n933), .B(G1348), .ZN(n943) );
  INV_X1 U1036 ( .A(n934), .ZN(n936) );
  NOR2_X1 U1037 ( .A1(n936), .A2(n935), .ZN(n939) );
  XOR2_X1 U1038 ( .A(G1341), .B(n937), .Z(n938) );
  NAND2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n941) );
  XNOR2_X1 U1040 ( .A(G1971), .B(G303), .ZN(n940) );
  NOR2_X1 U1041 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1042 ( .A1(n943), .A2(n942), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(G1966), .B(G168), .ZN(n945) );
  NAND2_X1 U1044 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1045 ( .A(KEYINPUT57), .B(n946), .Z(n947) );
  NOR2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n980) );
  INV_X1 U1049 ( .A(G16), .ZN(n978) );
  XNOR2_X1 U1050 ( .A(G1966), .B(G21), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(G5), .B(G1961), .ZN(n953) );
  NOR2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n966) );
  XOR2_X1 U1053 ( .A(G1341), .B(G19), .Z(n957) );
  XNOR2_X1 U1054 ( .A(n955), .B(G20), .ZN(n956) );
  NAND2_X1 U1055 ( .A1(n957), .A2(n956), .ZN(n963) );
  XOR2_X1 U1056 ( .A(G1981), .B(G6), .Z(n961) );
  XOR2_X1 U1057 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n958) );
  XNOR2_X1 U1058 ( .A(G4), .B(n958), .ZN(n959) );
  XNOR2_X1 U1059 ( .A(n959), .B(G1348), .ZN(n960) );
  NAND2_X1 U1060 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1061 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1062 ( .A(n964), .B(KEYINPUT60), .ZN(n965) );
  NAND2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n974) );
  XNOR2_X1 U1064 ( .A(G1971), .B(G22), .ZN(n968) );
  XNOR2_X1 U1065 ( .A(G23), .B(G1976), .ZN(n967) );
  NOR2_X1 U1066 ( .A1(n968), .A2(n967), .ZN(n971) );
  XOR2_X1 U1067 ( .A(G1986), .B(KEYINPUT126), .Z(n969) );
  XNOR2_X1 U1068 ( .A(G24), .B(n969), .ZN(n970) );
  NAND2_X1 U1069 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1070 ( .A(KEYINPUT58), .B(n972), .ZN(n973) );
  NOR2_X1 U1071 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1072 ( .A(n975), .B(KEYINPUT61), .Z(n976) );
  XNOR2_X1 U1073 ( .A(KEYINPUT127), .B(n976), .ZN(n977) );
  NAND2_X1 U1074 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n1036) );
  XNOR2_X1 U1076 ( .A(G2084), .B(G34), .ZN(n981) );
  XNOR2_X1 U1077 ( .A(n981), .B(KEYINPUT54), .ZN(n1001) );
  XNOR2_X1 U1078 ( .A(G2090), .B(G35), .ZN(n998) );
  XNOR2_X1 U1079 ( .A(G25), .B(G1991), .ZN(n982) );
  XNOR2_X1 U1080 ( .A(n982), .B(KEYINPUT119), .ZN(n988) );
  XOR2_X1 U1081 ( .A(G2072), .B(G33), .Z(n983) );
  NAND2_X1 U1082 ( .A1(n983), .A2(G28), .ZN(n986) );
  XNOR2_X1 U1083 ( .A(KEYINPUT120), .B(G2067), .ZN(n984) );
  XNOR2_X1 U1084 ( .A(G26), .B(n984), .ZN(n985) );
  NOR2_X1 U1085 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1086 ( .A1(n988), .A2(n987), .ZN(n995) );
  XOR2_X1 U1087 ( .A(n989), .B(G27), .Z(n992) );
  XOR2_X1 U1088 ( .A(n990), .B(G32), .Z(n991) );
  NOR2_X1 U1089 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1090 ( .A(n993), .B(KEYINPUT121), .ZN(n994) );
  NOR2_X1 U1091 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1092 ( .A(KEYINPUT53), .B(n996), .ZN(n997) );
  NOR2_X1 U1093 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1094 ( .A(KEYINPUT122), .B(n999), .Z(n1000) );
  NOR2_X1 U1095 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1096 ( .A(KEYINPUT55), .B(n1002), .ZN(n1004) );
  INV_X1 U1097 ( .A(G29), .ZN(n1003) );
  NAND2_X1 U1098 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1099 ( .A1(n1005), .A2(G11), .ZN(n1006) );
  XNOR2_X1 U1100 ( .A(n1006), .B(KEYINPUT123), .ZN(n1034) );
  XNOR2_X1 U1101 ( .A(G160), .B(G2084), .ZN(n1008) );
  NAND2_X1 U1102 ( .A1(n1008), .A2(n1007), .ZN(n1028) );
  XOR2_X1 U1103 ( .A(G2090), .B(G162), .Z(n1009) );
  NOR2_X1 U1104 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1105 ( .A(n1011), .B(KEYINPUT51), .ZN(n1012) );
  NOR2_X1 U1106 ( .A1(n1013), .A2(n1012), .ZN(n1026) );
  NOR2_X1 U1107 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1108 ( .A(KEYINPUT117), .B(n1016), .Z(n1017) );
  NAND2_X1 U1109 ( .A1(n1018), .A2(n1017), .ZN(n1024) );
  XOR2_X1 U1110 ( .A(G2072), .B(n1019), .Z(n1021) );
  XOR2_X1 U1111 ( .A(G164), .B(G2078), .Z(n1020) );
  NOR2_X1 U1112 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1113 ( .A(KEYINPUT50), .B(n1022), .Z(n1023) );
  NOR2_X1 U1114 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1115 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1116 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1117 ( .A(KEYINPUT52), .B(n1029), .Z(n1030) );
  NOR2_X1 U1118 ( .A1(KEYINPUT55), .A2(n1030), .ZN(n1031) );
  XOR2_X1 U1119 ( .A(KEYINPUT118), .B(n1031), .Z(n1032) );
  NAND2_X1 U1120 ( .A1(n1032), .A2(G29), .ZN(n1033) );
  NAND2_X1 U1121 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NOR2_X1 U1122 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XNOR2_X1 U1123 ( .A(n1037), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1124 ( .A(G311), .ZN(G150) );
endmodule

