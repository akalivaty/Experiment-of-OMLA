//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 1 0 1 1 1 1 1 1 1 0 0 0 1 1 0 0 1 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 1 0 0 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n458));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(G137), .A3(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n459), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  AND3_X1   g041(.A1(new_n464), .A2(KEYINPUT68), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g042(.A(KEYINPUT68), .B1(new_n464), .B2(new_n466), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n460), .A2(new_n461), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n469), .A2(new_n475), .ZN(G160));
  AOI21_X1  g051(.A(new_n463), .B1(new_n460), .B2(new_n461), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n480));
  INV_X1    g055(.A(G136), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n462), .A2(new_n463), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n478), .B(new_n480), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  NAND3_X1  g059(.A1(new_n462), .A2(G126), .A3(G2105), .ZN(new_n485));
  OR2_X1    g060(.A1(G102), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n463), .A2(G138), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT4), .B1(new_n471), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n462), .A2(new_n491), .A3(G138), .A4(new_n463), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n488), .B1(new_n490), .B2(new_n492), .ZN(G164));
  NAND2_X1  g068(.A1(G50), .A2(G543), .ZN(new_n494));
  INV_X1    g069(.A(G543), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT70), .B1(new_n495), .B2(KEYINPUT5), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT70), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n497), .A2(new_n498), .A3(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n501), .B1(new_n498), .B2(G543), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n495), .A2(KEYINPUT69), .A3(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G88), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n494), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(G75), .A2(G543), .ZN(new_n510));
  XOR2_X1   g085(.A(new_n510), .B(KEYINPUT71), .Z(new_n511));
  INV_X1    g086(.A(G62), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n505), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n509), .A2(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  INV_X1    g091(.A(G51), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n518));
  AND2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n524), .A2(KEYINPUT72), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n521), .A2(new_n526), .A3(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(KEYINPUT73), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT73), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n521), .A2(new_n526), .A3(new_n529), .A4(G543), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n517), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n500), .A2(new_n504), .A3(G89), .A4(new_n508), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n500), .A2(new_n504), .A3(G63), .A4(G651), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n531), .A2(new_n536), .ZN(G168));
  AOI22_X1  g112(.A1(new_n496), .A2(new_n499), .B1(new_n502), .B2(new_n503), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n538), .A2(G90), .A3(new_n508), .ZN(new_n539));
  AND2_X1   g114(.A1(G77), .A2(G543), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n540), .B1(new_n538), .B2(G64), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n539), .B1(new_n541), .B2(new_n523), .ZN(new_n542));
  INV_X1    g117(.A(G52), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n543), .B1(new_n528), .B2(new_n530), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n542), .A2(new_n544), .ZN(G171));
  NAND2_X1  g120(.A1(new_n528), .A2(new_n530), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G43), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n500), .A2(new_n504), .A3(G56), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AND3_X1   g125(.A1(new_n500), .A2(new_n504), .A3(new_n508), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n550), .A2(G651), .B1(new_n551), .B2(G81), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  NAND4_X1  g134(.A1(new_n521), .A2(new_n526), .A3(G53), .A4(G543), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n551), .A2(G91), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n505), .A2(KEYINPUT74), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT74), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n538), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n566), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n567));
  OAI211_X1 g142(.A(new_n561), .B(new_n562), .C1(new_n567), .C2(new_n523), .ZN(G299));
  INV_X1    g143(.A(G171), .ZN(G301));
  INV_X1    g144(.A(G168), .ZN(G286));
  NAND2_X1  g145(.A1(new_n551), .A2(G87), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n538), .B2(G74), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n495), .B1(new_n508), .B2(new_n518), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n573), .A2(G49), .A3(new_n526), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n571), .A2(new_n572), .A3(new_n574), .ZN(G288));
  AND2_X1   g150(.A1(new_n538), .A2(G86), .ZN(new_n576));
  AND2_X1   g151(.A1(G48), .A2(G543), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n508), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n505), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n578), .A2(new_n582), .ZN(G305));
  NAND2_X1  g158(.A1(new_n546), .A2(G47), .ZN(new_n584));
  NAND2_X1  g159(.A1(G72), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G60), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n505), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n587), .A2(G651), .B1(G85), .B2(new_n551), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n584), .A2(new_n588), .ZN(G290));
  INV_X1    g164(.A(G868), .ZN(new_n590));
  NOR2_X1   g165(.A1(G301), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n538), .A2(G92), .A3(new_n508), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n551), .A2(KEYINPUT10), .A3(G92), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n594), .A2(new_n595), .B1(new_n546), .B2(G54), .ZN(new_n596));
  INV_X1    g171(.A(G66), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n597), .B1(new_n563), .B2(new_n565), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(G651), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT75), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n591), .B1(new_n603), .B2(new_n590), .ZN(G284));
  AOI21_X1  g179(.A(new_n591), .B1(new_n603), .B2(new_n590), .ZN(G321));
  NAND2_X1  g180(.A1(G286), .A2(G868), .ZN(new_n606));
  AND3_X1   g181(.A1(new_n500), .A2(new_n504), .A3(new_n564), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n564), .B1(new_n500), .B2(new_n504), .ZN(new_n608));
  OAI21_X1  g183(.A(G65), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(G78), .A2(G543), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n523), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n560), .B(KEYINPUT9), .Z(new_n612));
  INV_X1    g187(.A(new_n562), .ZN(new_n613));
  NOR3_X1   g188(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n606), .B1(new_n614), .B2(G868), .ZN(G297));
  XNOR2_X1  g190(.A(G297), .B(KEYINPUT76), .ZN(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n603), .B1(new_n617), .B2(G860), .ZN(G148));
  NAND2_X1  g193(.A1(new_n603), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  OAI22_X1  g195(.A1(new_n620), .A2(KEYINPUT77), .B1(G868), .B2(new_n554), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(KEYINPUT77), .B2(new_n620), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT78), .Z(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n462), .A2(new_n465), .ZN(new_n625));
  XOR2_X1   g200(.A(KEYINPUT79), .B(KEYINPUT12), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  INV_X1    g203(.A(G2100), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n477), .A2(G123), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n463), .A2(G111), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  INV_X1    g209(.A(G135), .ZN(new_n635));
  OAI221_X1 g210(.A(new_n632), .B1(new_n633), .B2(new_n634), .C1(new_n635), .C2(new_n482), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND3_X1  g212(.A1(new_n630), .A2(new_n631), .A3(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(G2427), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G1341), .B(G1348), .Z(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n644), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n649), .B(new_n650), .Z(new_n651));
  OR2_X1    g226(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n648), .A2(new_n651), .ZN(new_n653));
  AND3_X1   g228(.A1(new_n652), .A2(G14), .A3(new_n653), .ZN(G401));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  XNOR2_X1  g230(.A(G2072), .B(G2078), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT18), .Z(new_n659));
  AOI21_X1  g234(.A(new_n657), .B1(new_n656), .B2(KEYINPUT81), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n660), .B1(KEYINPUT81), .B2(new_n656), .ZN(new_n661));
  INV_X1    g236(.A(new_n655), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n656), .B(KEYINPUT17), .Z(new_n663));
  INV_X1    g238(.A(new_n657), .ZN(new_n664));
  OAI211_X1 g239(.A(new_n661), .B(new_n662), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n663), .A2(new_n664), .A3(new_n655), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n659), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2096), .B(G2100), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G227));
  XOR2_X1   g244(.A(G1956), .B(G2474), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT82), .ZN(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n673), .A2(KEYINPUT83), .ZN(new_n674));
  XOR2_X1   g249(.A(G1971), .B(G1976), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(KEYINPUT83), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT20), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n671), .A2(new_n672), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(new_n673), .B2(new_n676), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT84), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n676), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1991), .B(G1996), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(G229));
  INV_X1    g267(.A(G16), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G6), .ZN(new_n694));
  INV_X1    g269(.A(G305), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n694), .B1(new_n695), .B2(new_n693), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT32), .B(G1981), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT86), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n696), .B(new_n698), .Z(new_n699));
  NAND2_X1  g274(.A1(new_n693), .A2(G22), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G166), .B2(new_n693), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(G1971), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n693), .A2(G23), .ZN(new_n703));
  INV_X1    g278(.A(G288), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(new_n693), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT33), .B(G1976), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n705), .B(new_n706), .Z(new_n707));
  NOR3_X1   g282(.A1(new_n699), .A2(new_n702), .A3(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT34), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n693), .A2(G24), .ZN(new_n712));
  INV_X1    g287(.A(G290), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(new_n693), .ZN(new_n714));
  INV_X1    g289(.A(G1986), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G25), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT85), .Z(new_n719));
  NAND2_X1  g294(.A1(new_n477), .A2(G119), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n463), .A2(G107), .ZN(new_n721));
  OAI21_X1  g296(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n722));
  INV_X1    g297(.A(G131), .ZN(new_n723));
  OAI221_X1 g298(.A(new_n720), .B1(new_n721), .B2(new_n722), .C1(new_n723), .C2(new_n482), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n719), .B1(new_n724), .B2(G29), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT35), .B(G1991), .Z(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n725), .B(new_n727), .ZN(new_n728));
  NAND4_X1  g303(.A1(new_n710), .A2(new_n711), .A3(new_n716), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT36), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n693), .A2(G20), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT23), .Z(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G299), .B2(G16), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G1956), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT25), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n462), .A2(G127), .ZN(new_n737));
  NAND2_X1  g312(.A1(G115), .A2(G2104), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n463), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(new_n482), .ZN(new_n740));
  AOI211_X1 g315(.A(new_n736), .B(new_n739), .C1(G139), .C2(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n741), .A2(new_n717), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n717), .B2(G33), .ZN(new_n743));
  INV_X1    g318(.A(G2072), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT91), .Z(new_n746));
  NAND2_X1  g321(.A1(new_n717), .A2(G27), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G164), .B2(new_n717), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT96), .Z(new_n749));
  OR2_X1    g324(.A1(new_n749), .A2(G2078), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT24), .B(G34), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(new_n717), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT90), .ZN(new_n753));
  INV_X1    g328(.A(G160), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n753), .B1(new_n754), .B2(new_n717), .ZN(new_n755));
  INV_X1    g330(.A(G2084), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n749), .A2(G2078), .ZN(new_n758));
  NAND4_X1  g333(.A1(new_n746), .A2(new_n750), .A3(new_n757), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n717), .A2(G32), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n477), .A2(G129), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n465), .A2(G105), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G141), .B2(new_n740), .ZN(new_n764));
  NAND3_X1  g339(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT92), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT26), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT93), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n760), .B1(new_n769), .B2(new_n717), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT27), .B(G1996), .ZN(new_n772));
  INV_X1    g347(.A(G1961), .ZN(new_n773));
  NOR2_X1   g348(.A1(G171), .A2(new_n693), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G5), .B2(new_n693), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n771), .A2(new_n772), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n772), .B2(new_n771), .ZN(new_n777));
  INV_X1    g352(.A(G28), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n778), .A2(KEYINPUT30), .ZN(new_n779));
  AOI21_X1  g354(.A(G29), .B1(new_n778), .B2(KEYINPUT30), .ZN(new_n780));
  OR2_X1    g355(.A1(KEYINPUT31), .A2(G11), .ZN(new_n781));
  NAND2_X1  g356(.A1(KEYINPUT31), .A2(G11), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n779), .A2(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(G29), .A2(G35), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G162), .B2(G29), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT97), .B(KEYINPUT29), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G2090), .ZN(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  OAI221_X1 g363(.A(new_n783), .B1(new_n717), .B2(new_n636), .C1(new_n785), .C2(new_n788), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n785), .A2(new_n788), .ZN(new_n790));
  AOI211_X1 g365(.A(new_n789), .B(new_n790), .C1(new_n743), .C2(new_n744), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n693), .A2(G21), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G168), .B2(new_n693), .ZN(new_n793));
  OAI221_X1 g368(.A(new_n791), .B1(G1966), .B2(new_n793), .C1(new_n756), .C2(new_n755), .ZN(new_n794));
  NOR3_X1   g369(.A1(new_n759), .A2(new_n777), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n793), .A2(G1966), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT94), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n775), .A2(new_n773), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT95), .ZN(new_n799));
  AND4_X1   g374(.A1(new_n734), .A2(new_n795), .A3(new_n797), .A4(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n603), .A2(new_n693), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G4), .B2(new_n693), .ZN(new_n802));
  INV_X1    g377(.A(G1348), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n717), .A2(G26), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT28), .Z(new_n806));
  OR2_X1    g381(.A1(G104), .A2(G2105), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n807), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT88), .Z(new_n809));
  AOI22_X1  g384(.A1(new_n740), .A2(G140), .B1(G128), .B2(new_n477), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n806), .B1(new_n811), .B2(G29), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G2067), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n802), .A2(new_n803), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n693), .A2(G19), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n554), .B2(new_n693), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT87), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G1341), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n804), .A2(new_n813), .A3(new_n814), .A4(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT89), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n730), .A2(new_n800), .A3(new_n820), .ZN(G150));
  INV_X1    g396(.A(G150), .ZN(G311));
  INV_X1    g397(.A(KEYINPUT39), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n603), .A2(G559), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT38), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n551), .A2(G81), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n538), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n827), .B2(new_n523), .ZN(new_n828));
  INV_X1    g403(.A(G43), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(new_n528), .B2(new_n530), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT98), .B(G93), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n538), .A2(new_n508), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(G80), .A2(G543), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n538), .B2(G67), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n832), .B1(new_n835), .B2(new_n523), .ZN(new_n836));
  INV_X1    g411(.A(G55), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(new_n528), .B2(new_n530), .ZN(new_n838));
  OAI22_X1  g413(.A1(new_n828), .A2(new_n830), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n529), .B1(new_n573), .B2(new_n526), .ZN(new_n840));
  INV_X1    g415(.A(new_n530), .ZN(new_n841));
  OAI21_X1  g416(.A(G55), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AND4_X1   g417(.A1(new_n504), .A2(new_n500), .A3(new_n508), .A4(new_n831), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n500), .A2(new_n504), .A3(G67), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(new_n833), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n843), .B1(new_n845), .B2(G651), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n547), .A2(new_n552), .A3(new_n842), .A4(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n839), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n825), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT38), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n824), .B(new_n850), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n839), .A2(new_n847), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n823), .B1(new_n849), .B2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(G860), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n851), .A2(new_n852), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n825), .A2(new_n848), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n857), .A2(new_n858), .A3(KEYINPUT39), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT99), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n857), .A2(new_n858), .A3(KEYINPUT99), .A4(KEYINPUT39), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n856), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n842), .A2(new_n846), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(G860), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT37), .ZN(new_n866));
  OAI21_X1  g441(.A(KEYINPUT100), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n868));
  INV_X1    g443(.A(new_n866), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n861), .A2(new_n862), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n868), .B(new_n869), .C1(new_n870), .C2(new_n856), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n867), .A2(new_n871), .ZN(G145));
  XNOR2_X1  g447(.A(new_n811), .B(G164), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n477), .A2(G130), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n463), .A2(G118), .ZN(new_n875));
  OAI21_X1  g450(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n740), .A2(KEYINPUT101), .A3(G142), .ZN(new_n877));
  AOI21_X1  g452(.A(KEYINPUT101), .B1(new_n740), .B2(G142), .ZN(new_n878));
  OAI221_X1 g453(.A(new_n874), .B1(new_n875), .B2(new_n876), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n873), .B(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n724), .B(new_n627), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n880), .B(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n769), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n741), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n884), .B1(new_n768), .B2(new_n741), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n882), .B(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(G160), .B(G162), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n636), .ZN(new_n888));
  AOI21_X1  g463(.A(G37), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n889), .B1(new_n888), .B2(new_n886), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT40), .ZN(G395));
  AOI21_X1  g466(.A(KEYINPUT105), .B1(new_n864), .B2(new_n590), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n848), .B(KEYINPUT102), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n619), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n619), .A2(new_n893), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n897), .B1(new_n614), .B2(new_n602), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT103), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n614), .A2(new_n602), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n594), .A2(new_n595), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n546), .A2(G54), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(G66), .B1(new_n607), .B2(new_n608), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n523), .B1(new_n904), .B2(new_n599), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(KEYINPUT103), .B1(new_n906), .B2(G299), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n898), .B1(new_n900), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n614), .A2(new_n602), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n906), .A2(G299), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n897), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n896), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n899), .B1(new_n614), .B2(new_n602), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n906), .A2(G299), .A3(KEYINPUT103), .ZN(new_n917));
  AOI22_X1  g492(.A1(new_n916), .A2(new_n917), .B1(new_n614), .B2(new_n602), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n894), .A2(new_n895), .A3(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(G290), .B(G303), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n704), .A2(KEYINPUT104), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n923));
  NAND2_X1  g498(.A1(G288), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n695), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n925), .A2(new_n695), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n921), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n928), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n930), .A2(new_n920), .A3(new_n926), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT42), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n929), .A2(new_n931), .A3(KEYINPUT42), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n915), .A2(new_n919), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(G868), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n936), .B1(new_n915), .B2(new_n919), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n892), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n939), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n941), .A2(KEYINPUT105), .A3(G868), .A4(new_n937), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n940), .A2(new_n942), .ZN(G295));
  AND3_X1   g518(.A1(new_n940), .A2(new_n942), .A3(KEYINPUT106), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT106), .B1(new_n940), .B2(new_n942), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(G331));
  INV_X1    g521(.A(new_n932), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n546), .A2(G51), .ZN(new_n948));
  OAI21_X1  g523(.A(G52), .B1(new_n840), .B2(new_n841), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n500), .A2(new_n504), .A3(G64), .ZN(new_n950));
  INV_X1    g525(.A(new_n540), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n952), .A2(G651), .B1(new_n551), .B2(G90), .ZN(new_n953));
  INV_X1    g528(.A(new_n536), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n948), .A2(new_n949), .A3(new_n953), .A4(new_n954), .ZN(new_n955));
  OAI22_X1  g530(.A1(new_n542), .A2(new_n544), .B1(new_n531), .B2(new_n536), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n848), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n839), .A2(new_n847), .A3(new_n955), .A4(new_n956), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n852), .A2(KEYINPUT107), .A3(new_n956), .A4(new_n955), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT109), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n909), .B1(new_n900), .B2(new_n907), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n964), .B1(new_n963), .B2(new_n965), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n898), .A2(new_n910), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(new_n918), .B2(KEYINPUT41), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n958), .A2(new_n971), .A3(new_n960), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n848), .A2(new_n957), .A3(KEYINPUT108), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n970), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n947), .B1(new_n968), .B2(new_n976), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n961), .A2(new_n962), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n913), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n974), .A2(new_n965), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n947), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G37), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT110), .B1(new_n977), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT109), .B1(new_n978), .B2(new_n918), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n963), .A2(new_n965), .A3(new_n964), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n976), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n932), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n989));
  AOI22_X1  g564(.A1(new_n913), .A2(new_n978), .B1(new_n965), .B2(new_n974), .ZN(new_n990));
  AOI21_X1  g565(.A(G37), .B1(new_n990), .B2(new_n947), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n988), .A2(new_n989), .A3(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n984), .A2(KEYINPUT43), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT111), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n984), .A2(KEYINPUT111), .A3(new_n992), .A4(KEYINPUT43), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT44), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n990), .A2(new_n947), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n983), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT43), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n997), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n995), .A2(new_n996), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n988), .A2(new_n1000), .A3(new_n991), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1003), .B1(new_n999), .B2(new_n1000), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n997), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1002), .A2(new_n1005), .ZN(G397));
  NAND2_X1  g581(.A1(new_n490), .A2(new_n492), .ZN(new_n1007));
  INV_X1    g582(.A(new_n488), .ZN(new_n1008));
  AOI21_X1  g583(.A(G1384), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT45), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n474), .B(G40), .C1(new_n467), .C2(new_n468), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G2067), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n811), .B(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n768), .ZN(new_n1017));
  INV_X1    g592(.A(G1996), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1019), .B1(new_n1018), .B2(new_n769), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n724), .B(new_n726), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1020), .B(new_n1021), .C1(new_n715), .C2(new_n713), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n713), .A2(new_n715), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1023), .B(KEYINPUT112), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1014), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT119), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1013), .B1(KEYINPUT45), .B2(new_n1009), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(new_n1009), .B2(KEYINPUT45), .ZN(new_n1029));
  OAI211_X1 g604(.A(KEYINPUT113), .B(new_n1011), .C1(G164), .C2(G1384), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1027), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G1971), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1013), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n1036));
  INV_X1    g611(.A(G1384), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n1033), .A2(new_n1034), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G2090), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n1031), .A2(new_n1032), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G8), .ZN(new_n1042));
  NAND2_X1  g617(.A1(KEYINPUT114), .A2(KEYINPUT55), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1043), .B1(G166), .B2(new_n1042), .ZN(new_n1044));
  XNOR2_X1  g619(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n1045));
  NAND3_X1  g620(.A1(G303), .A2(G8), .A3(new_n1045), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n1041), .A2(new_n1042), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1047), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1048), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(G8), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OAI211_X1 g629(.A(KEYINPUT115), .B(G8), .C1(new_n1010), .C2(new_n1013), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G1981), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n578), .A2(new_n1057), .A3(new_n582), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1057), .B1(new_n578), .B2(new_n582), .ZN(new_n1059));
  OAI21_X1  g634(.A(KEYINPUT49), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(G305), .A2(G1981), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT49), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n578), .A2(new_n1057), .A3(new_n582), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1060), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1056), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n704), .A2(G1976), .ZN(new_n1067));
  INV_X1    g642(.A(G1976), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT52), .B1(G288), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1033), .A2(new_n1009), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT115), .B1(new_n1070), .B2(G8), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1055), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1067), .B(new_n1069), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1066), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1075), .B1(new_n1056), .B2(new_n1067), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(KEYINPUT116), .B(new_n1047), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1027), .A2(new_n1012), .ZN(new_n1079));
  INV_X1    g654(.A(G1966), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT117), .B(G2084), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1039), .A2(new_n1082), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(G168), .A2(G8), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1051), .A2(new_n1077), .A3(new_n1078), .A4(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT63), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1047), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1091), .A2(new_n1092), .A3(G8), .ZN(new_n1093));
  AOI211_X1 g668(.A(new_n1088), .B(new_n1085), .C1(new_n1081), .C2(new_n1083), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1056), .A2(new_n1067), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT52), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1050), .A2(new_n1097), .A3(new_n1073), .A4(new_n1066), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1095), .B1(new_n1098), .B2(KEYINPUT118), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1077), .A2(new_n1100), .A3(new_n1050), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1087), .A2(new_n1088), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1077), .A2(new_n1048), .ZN(new_n1103));
  NOR2_X1   g678(.A1(G288), .A2(G1976), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1066), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1056), .B1(new_n1105), .B2(new_n1058), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1026), .B1(new_n1102), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1050), .A2(new_n1049), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1077), .A2(new_n1109), .A3(new_n1078), .A4(new_n1093), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1086), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1088), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1107), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1114), .A2(KEYINPUT119), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1108), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1033), .A2(new_n1034), .A3(new_n1038), .ZN(new_n1118));
  INV_X1    g693(.A(G1956), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g695(.A(KEYINPUT56), .B(G2072), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1027), .A2(new_n1029), .A3(new_n1030), .A4(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1120), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1124), .B1(new_n1123), .B2(new_n1122), .ZN(new_n1125));
  OAI211_X1 g700(.A(KEYINPUT120), .B(new_n562), .C1(new_n567), .C2(new_n523), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n611), .B2(new_n613), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1126), .A2(new_n1128), .A3(new_n561), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT57), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(new_n1131), .B2(G299), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1130), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1125), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(KEYINPUT61), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT61), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1125), .B(new_n1137), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1118), .A2(new_n803), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n602), .A2(KEYINPUT60), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1033), .A2(new_n1015), .A3(new_n1009), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT123), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1033), .A2(KEYINPUT123), .A3(new_n1015), .A4(new_n1009), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1139), .A2(new_n1140), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT59), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1027), .A2(new_n1018), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1147));
  XOR2_X1   g722(.A(KEYINPUT58), .B(G1341), .Z(new_n1148));
  NAND2_X1  g723(.A1(new_n1070), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1146), .B1(new_n1150), .B2(new_n554), .ZN(new_n1151));
  AOI211_X1 g726(.A(KEYINPUT59), .B(new_n553), .C1(new_n1147), .C2(new_n1149), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1145), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT60), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1139), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(new_n906), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1139), .A2(new_n1143), .A3(new_n1144), .A4(new_n602), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1154), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1153), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1136), .A2(new_n1138), .A3(new_n1159), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1125), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1156), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1161), .B1(new_n1135), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1164));
  AND2_X1   g739(.A1(new_n1027), .A2(new_n1012), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT53), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1166), .A2(G2078), .ZN(new_n1167));
  AOI22_X1  g742(.A1(new_n1165), .A2(new_n1167), .B1(new_n773), .B2(new_n1118), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1166), .B1(new_n1031), .B2(G2078), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(G171), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1170), .A2(G171), .ZN(new_n1173));
  OAI21_X1  g748(.A(KEYINPUT54), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1173), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT54), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1175), .A2(new_n1176), .A3(new_n1171), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1042), .B1(new_n1084), .B2(G168), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(G286), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(KEYINPUT51), .ZN(new_n1182));
  AOI211_X1 g757(.A(KEYINPUT51), .B(new_n1042), .C1(new_n1084), .C2(G168), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1183), .ZN(new_n1184));
  AOI22_X1  g759(.A1(new_n1174), .A2(new_n1177), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1164), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT51), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1187), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1188));
  OR3_X1    g763(.A1(new_n1188), .A2(KEYINPUT62), .A3(new_n1183), .ZN(new_n1189));
  OAI21_X1  g764(.A(KEYINPUT62), .B1(new_n1188), .B2(new_n1183), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1189), .A2(new_n1172), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1110), .B1(new_n1186), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1025), .B1(new_n1117), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT46), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n1196), .B(KEYINPUT124), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1198));
  AOI22_X1  g773(.A1(new_n1195), .A2(new_n1194), .B1(new_n1198), .B2(new_n1014), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n1200), .B(KEYINPUT125), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT47), .ZN(new_n1202));
  OR2_X1    g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1204));
  INV_X1    g779(.A(new_n1014), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n724), .A2(new_n727), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1020), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n809), .A2(new_n1015), .A3(new_n810), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1205), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1205), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1024), .A2(new_n1014), .ZN(new_n1211));
  INV_X1    g786(.A(new_n1211), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1210), .B1(KEYINPUT48), .B2(new_n1212), .ZN(new_n1213));
  OR2_X1    g788(.A1(new_n1212), .A2(KEYINPUT48), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1209), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  AND3_X1   g790(.A1(new_n1203), .A2(new_n1204), .A3(new_n1215), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1193), .A2(new_n1216), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g792(.A(G319), .ZN(new_n1219));
  NOR2_X1   g793(.A1(G227), .A2(new_n1219), .ZN(new_n1220));
  XOR2_X1   g794(.A(new_n1220), .B(KEYINPUT126), .Z(new_n1221));
  NOR2_X1   g795(.A1(new_n1221), .A2(G401), .ZN(new_n1222));
  XNOR2_X1  g796(.A(new_n1222), .B(KEYINPUT127), .ZN(new_n1223));
  NAND4_X1  g797(.A1(new_n691), .A2(new_n890), .A3(new_n1004), .A4(new_n1223), .ZN(G225));
  INV_X1    g798(.A(G225), .ZN(G308));
endmodule


