

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U557 ( .A1(G2104), .A2(n541), .ZN(n880) );
  NOR2_X2 U558 ( .A1(G2105), .A2(G2104), .ZN(n537) );
  XNOR2_X1 U559 ( .A(n702), .B(n701), .ZN(n708) );
  INV_X1 U560 ( .A(KEYINPUT13), .ZN(n558) );
  NOR2_X1 U561 ( .A1(n691), .A2(n954), .ZN(n698) );
  OR2_X1 U562 ( .A1(n898), .A2(n698), .ZN(n699) );
  INV_X1 U563 ( .A(KEYINPUT99), .ZN(n701) );
  BUF_X1 U564 ( .A(n692), .Z(n715) );
  XNOR2_X1 U565 ( .A(n722), .B(KEYINPUT30), .ZN(n723) );
  XNOR2_X1 U566 ( .A(KEYINPUT31), .B(KEYINPUT100), .ZN(n726) );
  XNOR2_X1 U567 ( .A(n727), .B(n726), .ZN(n728) );
  AND2_X1 U568 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X2 U569 ( .A1(n687), .A2(n778), .ZN(n692) );
  NAND2_X1 U570 ( .A1(G8), .A2(n739), .ZN(n802) );
  NOR2_X1 U571 ( .A1(G1384), .A2(G164), .ZN(n683) );
  NOR2_X1 U572 ( .A1(G651), .A2(G543), .ZN(n524) );
  XNOR2_X1 U573 ( .A(n559), .B(n558), .ZN(n563) );
  NOR2_X1 U574 ( .A1(G651), .A2(n652), .ZN(n646) );
  NAND2_X1 U575 ( .A1(n566), .A2(n565), .ZN(n954) );
  XOR2_X1 U576 ( .A(KEYINPUT65), .B(n524), .Z(n636) );
  NAND2_X1 U577 ( .A1(n636), .A2(G89), .ZN(n525) );
  XNOR2_X1 U578 ( .A(n525), .B(KEYINPUT4), .ZN(n527) );
  XOR2_X1 U579 ( .A(G543), .B(KEYINPUT0), .Z(n652) );
  INV_X1 U580 ( .A(G651), .ZN(n529) );
  NOR2_X1 U581 ( .A1(n652), .A2(n529), .ZN(n639) );
  NAND2_X1 U582 ( .A1(G76), .A2(n639), .ZN(n526) );
  NAND2_X1 U583 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U584 ( .A(n528), .B(KEYINPUT5), .ZN(n535) );
  NAND2_X1 U585 ( .A1(G51), .A2(n646), .ZN(n532) );
  NOR2_X1 U586 ( .A1(G543), .A2(n529), .ZN(n530) );
  XOR2_X1 U587 ( .A(KEYINPUT1), .B(n530), .Z(n650) );
  NAND2_X1 U588 ( .A1(G63), .A2(n650), .ZN(n531) );
  NAND2_X1 U589 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U590 ( .A(KEYINPUT6), .B(n533), .Z(n534) );
  NAND2_X1 U591 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U592 ( .A(n536), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X2 U593 ( .A(KEYINPUT17), .B(n537), .Z(n889) );
  NAND2_X1 U594 ( .A1(G138), .A2(n889), .ZN(n539) );
  INV_X1 U595 ( .A(G2104), .ZN(n540) );
  NOR2_X1 U596 ( .A1(G2105), .A2(n540), .ZN(n886) );
  NAND2_X1 U597 ( .A1(G102), .A2(n886), .ZN(n538) );
  NAND2_X1 U598 ( .A1(n539), .A2(n538), .ZN(n545) );
  INV_X1 U599 ( .A(G2105), .ZN(n541) );
  NAND2_X1 U600 ( .A1(G126), .A2(n880), .ZN(n543) );
  NOR2_X1 U601 ( .A1(n541), .A2(n540), .ZN(n882) );
  NAND2_X1 U602 ( .A1(G114), .A2(n882), .ZN(n542) );
  NAND2_X1 U603 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X1 U604 ( .A1(n545), .A2(n544), .ZN(G164) );
  NAND2_X1 U605 ( .A1(G137), .A2(n889), .ZN(n547) );
  NAND2_X1 U606 ( .A1(G113), .A2(n882), .ZN(n546) );
  NAND2_X1 U607 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U608 ( .A(KEYINPUT66), .B(n548), .Z(n550) );
  NAND2_X1 U609 ( .A1(n880), .A2(G125), .ZN(n549) );
  AND2_X1 U610 ( .A1(n550), .A2(n549), .ZN(n686) );
  NAND2_X1 U611 ( .A1(G101), .A2(n886), .ZN(n551) );
  XOR2_X1 U612 ( .A(KEYINPUT23), .B(n551), .Z(n684) );
  AND2_X1 U613 ( .A1(n686), .A2(n684), .ZN(G160) );
  AND2_X1 U614 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U615 ( .A(G57), .ZN(G237) );
  INV_X1 U616 ( .A(G132), .ZN(G219) );
  XOR2_X1 U617 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U618 ( .A1(G7), .A2(G661), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n552), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U620 ( .A(KEYINPUT11), .B(KEYINPUT74), .Z(n554) );
  INV_X1 U621 ( .A(G223), .ZN(n828) );
  NAND2_X1 U622 ( .A1(G567), .A2(n828), .ZN(n553) );
  XNOR2_X1 U623 ( .A(n554), .B(n553), .ZN(G234) );
  NAND2_X1 U624 ( .A1(n636), .A2(G81), .ZN(n555) );
  XNOR2_X1 U625 ( .A(n555), .B(KEYINPUT12), .ZN(n557) );
  NAND2_X1 U626 ( .A1(G68), .A2(n639), .ZN(n556) );
  NAND2_X1 U627 ( .A1(n557), .A2(n556), .ZN(n559) );
  NAND2_X1 U628 ( .A1(G56), .A2(n650), .ZN(n560) );
  XNOR2_X1 U629 ( .A(n560), .B(KEYINPUT75), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n561), .B(KEYINPUT14), .ZN(n562) );
  NOR2_X1 U631 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n564), .B(KEYINPUT76), .ZN(n566) );
  NAND2_X1 U633 ( .A1(G43), .A2(n646), .ZN(n565) );
  INV_X1 U634 ( .A(G860), .ZN(n611) );
  OR2_X1 U635 ( .A1(n954), .A2(n611), .ZN(G153) );
  NAND2_X1 U636 ( .A1(G52), .A2(n646), .ZN(n568) );
  NAND2_X1 U637 ( .A1(G64), .A2(n650), .ZN(n567) );
  NAND2_X1 U638 ( .A1(n568), .A2(n567), .ZN(n573) );
  NAND2_X1 U639 ( .A1(G90), .A2(n636), .ZN(n570) );
  NAND2_X1 U640 ( .A1(G77), .A2(n639), .ZN(n569) );
  NAND2_X1 U641 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U642 ( .A(KEYINPUT9), .B(n571), .Z(n572) );
  NOR2_X1 U643 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U644 ( .A(KEYINPUT70), .B(n574), .Z(G301) );
  NAND2_X1 U645 ( .A1(G301), .A2(G868), .ZN(n584) );
  NAND2_X1 U646 ( .A1(G66), .A2(n650), .ZN(n581) );
  NAND2_X1 U647 ( .A1(G54), .A2(n646), .ZN(n576) );
  NAND2_X1 U648 ( .A1(G92), .A2(n636), .ZN(n575) );
  NAND2_X1 U649 ( .A1(n576), .A2(n575), .ZN(n579) );
  NAND2_X1 U650 ( .A1(G79), .A2(n639), .ZN(n577) );
  XNOR2_X1 U651 ( .A(KEYINPUT77), .B(n577), .ZN(n578) );
  NOR2_X1 U652 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U653 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U654 ( .A(n582), .B(KEYINPUT15), .ZN(n898) );
  INV_X1 U655 ( .A(n898), .ZN(n957) );
  INV_X1 U656 ( .A(G868), .ZN(n664) );
  NAND2_X1 U657 ( .A1(n957), .A2(n664), .ZN(n583) );
  NAND2_X1 U658 ( .A1(n584), .A2(n583), .ZN(G284) );
  NAND2_X1 U659 ( .A1(n639), .A2(G78), .ZN(n587) );
  NAND2_X1 U660 ( .A1(G53), .A2(n646), .ZN(n585) );
  XOR2_X1 U661 ( .A(KEYINPUT71), .B(n585), .Z(n586) );
  NAND2_X1 U662 ( .A1(n587), .A2(n586), .ZN(n591) );
  NAND2_X1 U663 ( .A1(G91), .A2(n636), .ZN(n589) );
  NAND2_X1 U664 ( .A1(G65), .A2(n650), .ZN(n588) );
  NAND2_X1 U665 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U666 ( .A1(n591), .A2(n590), .ZN(n943) );
  XOR2_X1 U667 ( .A(n943), .B(KEYINPUT72), .Z(G299) );
  NOR2_X1 U668 ( .A1(G868), .A2(G299), .ZN(n593) );
  NOR2_X1 U669 ( .A1(G286), .A2(n664), .ZN(n592) );
  NOR2_X1 U670 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U671 ( .A(KEYINPUT78), .B(n594), .ZN(G297) );
  NAND2_X1 U672 ( .A1(n611), .A2(G559), .ZN(n595) );
  NAND2_X1 U673 ( .A1(n595), .A2(n898), .ZN(n596) );
  XNOR2_X1 U674 ( .A(n596), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U675 ( .A1(G868), .A2(n954), .ZN(n599) );
  NAND2_X1 U676 ( .A1(G868), .A2(n898), .ZN(n597) );
  NOR2_X1 U677 ( .A1(G559), .A2(n597), .ZN(n598) );
  NOR2_X1 U678 ( .A1(n599), .A2(n598), .ZN(G282) );
  NAND2_X1 U679 ( .A1(G111), .A2(n882), .ZN(n606) );
  NAND2_X1 U680 ( .A1(G135), .A2(n889), .ZN(n601) );
  NAND2_X1 U681 ( .A1(G99), .A2(n886), .ZN(n600) );
  NAND2_X1 U682 ( .A1(n601), .A2(n600), .ZN(n604) );
  NAND2_X1 U683 ( .A1(n880), .A2(G123), .ZN(n602) );
  XOR2_X1 U684 ( .A(KEYINPUT18), .B(n602), .Z(n603) );
  NOR2_X1 U685 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U686 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U687 ( .A(n607), .B(KEYINPUT79), .ZN(n1008) );
  XNOR2_X1 U688 ( .A(n1008), .B(G2096), .ZN(n609) );
  INV_X1 U689 ( .A(G2100), .ZN(n608) );
  NAND2_X1 U690 ( .A1(n609), .A2(n608), .ZN(G156) );
  NAND2_X1 U691 ( .A1(G559), .A2(n898), .ZN(n610) );
  XOR2_X1 U692 ( .A(n954), .B(n610), .Z(n662) );
  NAND2_X1 U693 ( .A1(n611), .A2(n662), .ZN(n619) );
  NAND2_X1 U694 ( .A1(G93), .A2(n636), .ZN(n613) );
  NAND2_X1 U695 ( .A1(G80), .A2(n639), .ZN(n612) );
  NAND2_X1 U696 ( .A1(n613), .A2(n612), .ZN(n616) );
  NAND2_X1 U697 ( .A1(n646), .A2(G55), .ZN(n614) );
  XOR2_X1 U698 ( .A(KEYINPUT80), .B(n614), .Z(n615) );
  NOR2_X1 U699 ( .A1(n616), .A2(n615), .ZN(n618) );
  NAND2_X1 U700 ( .A1(n650), .A2(G67), .ZN(n617) );
  NAND2_X1 U701 ( .A1(n618), .A2(n617), .ZN(n665) );
  XNOR2_X1 U702 ( .A(n619), .B(n665), .ZN(G145) );
  NAND2_X1 U703 ( .A1(G86), .A2(n636), .ZN(n621) );
  NAND2_X1 U704 ( .A1(G61), .A2(n650), .ZN(n620) );
  NAND2_X1 U705 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U706 ( .A1(n639), .A2(G73), .ZN(n622) );
  XOR2_X1 U707 ( .A(KEYINPUT2), .B(n622), .Z(n623) );
  NOR2_X1 U708 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U709 ( .A1(n646), .A2(G48), .ZN(n625) );
  NAND2_X1 U710 ( .A1(n626), .A2(n625), .ZN(G305) );
  NAND2_X1 U711 ( .A1(n639), .A2(G72), .ZN(n634) );
  NAND2_X1 U712 ( .A1(G47), .A2(n646), .ZN(n627) );
  XNOR2_X1 U713 ( .A(n627), .B(KEYINPUT68), .ZN(n629) );
  NAND2_X1 U714 ( .A1(n650), .A2(G60), .ZN(n628) );
  NAND2_X1 U715 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U716 ( .A1(G85), .A2(n636), .ZN(n630) );
  XNOR2_X1 U717 ( .A(KEYINPUT67), .B(n630), .ZN(n631) );
  NOR2_X1 U718 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U719 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U720 ( .A(KEYINPUT69), .B(n635), .Z(G290) );
  NAND2_X1 U721 ( .A1(G62), .A2(n650), .ZN(n644) );
  NAND2_X1 U722 ( .A1(G50), .A2(n646), .ZN(n638) );
  NAND2_X1 U723 ( .A1(G88), .A2(n636), .ZN(n637) );
  NAND2_X1 U724 ( .A1(n638), .A2(n637), .ZN(n642) );
  NAND2_X1 U725 ( .A1(n639), .A2(G75), .ZN(n640) );
  XOR2_X1 U726 ( .A(KEYINPUT82), .B(n640), .Z(n641) );
  NOR2_X1 U727 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U728 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U729 ( .A(n645), .B(KEYINPUT83), .ZN(G166) );
  NAND2_X1 U730 ( .A1(G49), .A2(n646), .ZN(n648) );
  NAND2_X1 U731 ( .A1(G74), .A2(G651), .ZN(n647) );
  NAND2_X1 U732 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U733 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U734 ( .A(KEYINPUT81), .B(n651), .Z(n654) );
  NAND2_X1 U735 ( .A1(n652), .A2(G87), .ZN(n653) );
  NAND2_X1 U736 ( .A1(n654), .A2(n653), .ZN(G288) );
  XNOR2_X1 U737 ( .A(KEYINPUT19), .B(KEYINPUT84), .ZN(n656) );
  XNOR2_X1 U738 ( .A(G305), .B(KEYINPUT85), .ZN(n655) );
  XNOR2_X1 U739 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U740 ( .A(G299), .B(n657), .ZN(n659) );
  XNOR2_X1 U741 ( .A(G290), .B(G166), .ZN(n658) );
  XNOR2_X1 U742 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U743 ( .A(n660), .B(G288), .ZN(n661) );
  XNOR2_X1 U744 ( .A(n661), .B(n665), .ZN(n897) );
  XNOR2_X1 U745 ( .A(n897), .B(n662), .ZN(n663) );
  NOR2_X1 U746 ( .A1(n664), .A2(n663), .ZN(n667) );
  NOR2_X1 U747 ( .A1(G868), .A2(n665), .ZN(n666) );
  NOR2_X1 U748 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U749 ( .A(KEYINPUT86), .B(n668), .ZN(G295) );
  NAND2_X1 U750 ( .A1(G2084), .A2(G2078), .ZN(n669) );
  XOR2_X1 U751 ( .A(KEYINPUT20), .B(n669), .Z(n670) );
  NAND2_X1 U752 ( .A1(G2090), .A2(n670), .ZN(n671) );
  XNOR2_X1 U753 ( .A(KEYINPUT21), .B(n671), .ZN(n672) );
  NAND2_X1 U754 ( .A1(n672), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U755 ( .A(KEYINPUT73), .B(G82), .ZN(G220) );
  XNOR2_X1 U756 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U757 ( .A1(G219), .A2(G220), .ZN(n674) );
  XNOR2_X1 U758 ( .A(KEYINPUT87), .B(KEYINPUT22), .ZN(n673) );
  XNOR2_X1 U759 ( .A(n674), .B(n673), .ZN(n675) );
  NOR2_X1 U760 ( .A1(n675), .A2(G218), .ZN(n676) );
  NAND2_X1 U761 ( .A1(G96), .A2(n676), .ZN(n834) );
  NAND2_X1 U762 ( .A1(n834), .A2(G2106), .ZN(n681) );
  NAND2_X1 U763 ( .A1(G120), .A2(G108), .ZN(n677) );
  NOR2_X1 U764 ( .A1(G237), .A2(n677), .ZN(n678) );
  NAND2_X1 U765 ( .A1(G69), .A2(n678), .ZN(n833) );
  NAND2_X1 U766 ( .A1(G567), .A2(n833), .ZN(n679) );
  XNOR2_X1 U767 ( .A(KEYINPUT88), .B(n679), .ZN(n680) );
  NAND2_X1 U768 ( .A1(n681), .A2(n680), .ZN(n835) );
  NAND2_X1 U769 ( .A1(G483), .A2(G661), .ZN(n682) );
  NOR2_X1 U770 ( .A1(n835), .A2(n682), .ZN(n832) );
  NAND2_X1 U771 ( .A1(n832), .A2(G36), .ZN(G176) );
  INV_X1 U772 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U773 ( .A(n683), .B(KEYINPUT64), .ZN(n779) );
  INV_X1 U774 ( .A(n779), .ZN(n687) );
  AND2_X1 U775 ( .A1(n684), .A2(G40), .ZN(n685) );
  NAND2_X1 U776 ( .A1(n686), .A2(n685), .ZN(n778) );
  INV_X1 U777 ( .A(n692), .ZN(n739) );
  NOR2_X1 U778 ( .A1(G1966), .A2(n802), .ZN(n730) );
  AND2_X1 U779 ( .A1(n692), .A2(G1996), .ZN(n688) );
  XOR2_X1 U780 ( .A(KEYINPUT26), .B(n688), .Z(n690) );
  NAND2_X1 U781 ( .A1(n739), .A2(G1341), .ZN(n689) );
  NAND2_X1 U782 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U783 ( .A1(n698), .A2(n898), .ZN(n697) );
  AND2_X1 U784 ( .A1(n715), .A2(G2067), .ZN(n693) );
  XOR2_X1 U785 ( .A(n693), .B(KEYINPUT98), .Z(n695) );
  NAND2_X1 U786 ( .A1(n739), .A2(G1348), .ZN(n694) );
  NAND2_X1 U787 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U788 ( .A1(n697), .A2(n696), .ZN(n700) );
  NAND2_X1 U789 ( .A1(n700), .A2(n699), .ZN(n702) );
  XOR2_X1 U790 ( .A(KEYINPUT97), .B(KEYINPUT27), .Z(n704) );
  NAND2_X1 U791 ( .A1(G2072), .A2(n715), .ZN(n703) );
  XNOR2_X1 U792 ( .A(n704), .B(n703), .ZN(n706) );
  INV_X1 U793 ( .A(G1956), .ZN(n978) );
  NOR2_X1 U794 ( .A1(n715), .A2(n978), .ZN(n705) );
  NOR2_X1 U795 ( .A1(n706), .A2(n705), .ZN(n709) );
  NAND2_X1 U796 ( .A1(n709), .A2(n943), .ZN(n707) );
  NAND2_X1 U797 ( .A1(n708), .A2(n707), .ZN(n712) );
  NOR2_X1 U798 ( .A1(n709), .A2(n943), .ZN(n710) );
  XOR2_X1 U799 ( .A(n710), .B(KEYINPUT28), .Z(n711) );
  NAND2_X1 U800 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U801 ( .A(n713), .B(KEYINPUT29), .ZN(n719) );
  XNOR2_X1 U802 ( .A(G2078), .B(KEYINPUT25), .ZN(n925) );
  NAND2_X1 U803 ( .A1(n715), .A2(n925), .ZN(n714) );
  XOR2_X1 U804 ( .A(KEYINPUT96), .B(n714), .Z(n717) );
  NOR2_X1 U805 ( .A1(n715), .A2(G1961), .ZN(n716) );
  NOR2_X1 U806 ( .A1(n717), .A2(n716), .ZN(n720) );
  NOR2_X1 U807 ( .A1(G301), .A2(n720), .ZN(n718) );
  NOR2_X1 U808 ( .A1(n719), .A2(n718), .ZN(n729) );
  AND2_X1 U809 ( .A1(G301), .A2(n720), .ZN(n725) );
  NOR2_X1 U810 ( .A1(G2084), .A2(n739), .ZN(n731) );
  NOR2_X1 U811 ( .A1(n730), .A2(n731), .ZN(n721) );
  NAND2_X1 U812 ( .A1(G8), .A2(n721), .ZN(n722) );
  NOR2_X1 U813 ( .A1(n723), .A2(G168), .ZN(n724) );
  NOR2_X1 U814 ( .A1(n725), .A2(n724), .ZN(n727) );
  NOR2_X1 U815 ( .A1(n729), .A2(n728), .ZN(n735) );
  NOR2_X1 U816 ( .A1(n730), .A2(n735), .ZN(n733) );
  NAND2_X1 U817 ( .A1(G8), .A2(n731), .ZN(n732) );
  XNOR2_X1 U818 ( .A(KEYINPUT101), .B(n734), .ZN(n749) );
  INV_X1 U819 ( .A(n735), .ZN(n737) );
  AND2_X1 U820 ( .A1(G286), .A2(G8), .ZN(n736) );
  NAND2_X1 U821 ( .A1(n737), .A2(n736), .ZN(n746) );
  INV_X1 U822 ( .A(G8), .ZN(n744) );
  NOR2_X1 U823 ( .A1(G1971), .A2(n802), .ZN(n738) );
  XNOR2_X1 U824 ( .A(n738), .B(KEYINPUT102), .ZN(n741) );
  NOR2_X1 U825 ( .A1(n739), .A2(G2090), .ZN(n740) );
  NOR2_X1 U826 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U827 ( .A1(n742), .A2(G303), .ZN(n743) );
  OR2_X1 U828 ( .A1(n744), .A2(n743), .ZN(n745) );
  AND2_X1 U829 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U830 ( .A(n747), .B(KEYINPUT32), .ZN(n748) );
  NAND2_X1 U831 ( .A1(n749), .A2(n748), .ZN(n797) );
  NOR2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n946) );
  NOR2_X1 U833 ( .A1(G1971), .A2(G303), .ZN(n959) );
  NOR2_X1 U834 ( .A1(n946), .A2(n959), .ZN(n750) );
  NAND2_X1 U835 ( .A1(n797), .A2(n750), .ZN(n751) );
  XNOR2_X1 U836 ( .A(n751), .B(KEYINPUT103), .ZN(n754) );
  NAND2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n947) );
  INV_X1 U838 ( .A(n802), .ZN(n752) );
  NAND2_X1 U839 ( .A1(n947), .A2(n752), .ZN(n753) );
  NOR2_X1 U840 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U841 ( .A1(n755), .A2(KEYINPUT33), .ZN(n758) );
  NAND2_X1 U842 ( .A1(n946), .A2(KEYINPUT33), .ZN(n756) );
  NOR2_X1 U843 ( .A1(n756), .A2(n802), .ZN(n757) );
  NOR2_X1 U844 ( .A1(n758), .A2(n757), .ZN(n794) );
  XOR2_X1 U845 ( .A(G1981), .B(G305), .Z(n962) );
  NAND2_X1 U846 ( .A1(G131), .A2(n889), .ZN(n760) );
  NAND2_X1 U847 ( .A1(G107), .A2(n882), .ZN(n759) );
  NAND2_X1 U848 ( .A1(n760), .A2(n759), .ZN(n764) );
  NAND2_X1 U849 ( .A1(G95), .A2(n886), .ZN(n762) );
  NAND2_X1 U850 ( .A1(G119), .A2(n880), .ZN(n761) );
  NAND2_X1 U851 ( .A1(n762), .A2(n761), .ZN(n763) );
  OR2_X1 U852 ( .A1(n764), .A2(n763), .ZN(n863) );
  NAND2_X1 U853 ( .A1(G1991), .A2(n863), .ZN(n776) );
  XOR2_X1 U854 ( .A(KEYINPUT91), .B(KEYINPUT38), .Z(n766) );
  NAND2_X1 U855 ( .A1(G105), .A2(n886), .ZN(n765) );
  XNOR2_X1 U856 ( .A(n766), .B(n765), .ZN(n773) );
  NAND2_X1 U857 ( .A1(G117), .A2(n882), .ZN(n768) );
  NAND2_X1 U858 ( .A1(G129), .A2(n880), .ZN(n767) );
  NAND2_X1 U859 ( .A1(n768), .A2(n767), .ZN(n771) );
  NAND2_X1 U860 ( .A1(n889), .A2(G141), .ZN(n769) );
  XOR2_X1 U861 ( .A(KEYINPUT92), .B(n769), .Z(n770) );
  NOR2_X1 U862 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U863 ( .A1(n773), .A2(n772), .ZN(n862) );
  NAND2_X1 U864 ( .A1(G1996), .A2(n862), .ZN(n774) );
  XOR2_X1 U865 ( .A(KEYINPUT93), .B(n774), .Z(n775) );
  NAND2_X1 U866 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U867 ( .A(KEYINPUT94), .B(n777), .Z(n811) );
  XOR2_X1 U868 ( .A(G1986), .B(G290), .Z(n961) );
  NAND2_X1 U869 ( .A1(n811), .A2(n961), .ZN(n780) );
  NOR2_X1 U870 ( .A1(n779), .A2(n778), .ZN(n823) );
  NAND2_X1 U871 ( .A1(n780), .A2(n823), .ZN(n792) );
  NAND2_X1 U872 ( .A1(G140), .A2(n889), .ZN(n782) );
  NAND2_X1 U873 ( .A1(G104), .A2(n886), .ZN(n781) );
  NAND2_X1 U874 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U875 ( .A(KEYINPUT34), .B(n783), .ZN(n790) );
  XNOR2_X1 U876 ( .A(KEYINPUT90), .B(KEYINPUT35), .ZN(n788) );
  NAND2_X1 U877 ( .A1(n880), .A2(G128), .ZN(n786) );
  NAND2_X1 U878 ( .A1(n882), .A2(G116), .ZN(n784) );
  XOR2_X1 U879 ( .A(KEYINPUT89), .B(n784), .Z(n785) );
  NAND2_X1 U880 ( .A1(n786), .A2(n785), .ZN(n787) );
  XOR2_X1 U881 ( .A(n788), .B(n787), .Z(n789) );
  NOR2_X1 U882 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U883 ( .A(KEYINPUT36), .B(n791), .ZN(n868) );
  XNOR2_X1 U884 ( .A(G2067), .B(KEYINPUT37), .ZN(n820) );
  NOR2_X1 U885 ( .A1(n868), .A2(n820), .ZN(n1013) );
  NAND2_X1 U886 ( .A1(n823), .A2(n1013), .ZN(n818) );
  AND2_X1 U887 ( .A1(n792), .A2(n818), .ZN(n807) );
  AND2_X1 U888 ( .A1(n962), .A2(n807), .ZN(n793) );
  NAND2_X1 U889 ( .A1(n794), .A2(n793), .ZN(n809) );
  NOR2_X1 U890 ( .A1(G2090), .A2(G303), .ZN(n795) );
  XNOR2_X1 U891 ( .A(n795), .B(KEYINPUT104), .ZN(n796) );
  NAND2_X1 U892 ( .A1(n796), .A2(G8), .ZN(n798) );
  NAND2_X1 U893 ( .A1(n798), .A2(n797), .ZN(n799) );
  NAND2_X1 U894 ( .A1(n799), .A2(n802), .ZN(n805) );
  NOR2_X1 U895 ( .A1(G1981), .A2(G305), .ZN(n800) );
  XOR2_X1 U896 ( .A(n800), .B(KEYINPUT24), .Z(n801) );
  NOR2_X1 U897 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U898 ( .A(KEYINPUT95), .B(n803), .ZN(n804) );
  NAND2_X1 U899 ( .A1(n805), .A2(n804), .ZN(n806) );
  NAND2_X1 U900 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U901 ( .A1(n809), .A2(n808), .ZN(n810) );
  XNOR2_X1 U902 ( .A(n810), .B(KEYINPUT105), .ZN(n826) );
  INV_X1 U903 ( .A(n811), .ZN(n1025) );
  NOR2_X1 U904 ( .A1(G1991), .A2(n863), .ZN(n812) );
  XOR2_X1 U905 ( .A(KEYINPUT107), .B(n812), .Z(n1007) );
  NOR2_X1 U906 ( .A1(G1986), .A2(G290), .ZN(n813) );
  NOR2_X1 U907 ( .A1(n1007), .A2(n813), .ZN(n814) );
  NOR2_X1 U908 ( .A1(n1025), .A2(n814), .ZN(n816) );
  NOR2_X1 U909 ( .A1(n862), .A2(G1996), .ZN(n815) );
  XNOR2_X1 U910 ( .A(n815), .B(KEYINPUT106), .ZN(n1017) );
  NOR2_X1 U911 ( .A1(n816), .A2(n1017), .ZN(n817) );
  XNOR2_X1 U912 ( .A(n817), .B(KEYINPUT39), .ZN(n819) );
  NAND2_X1 U913 ( .A1(n819), .A2(n818), .ZN(n821) );
  NAND2_X1 U914 ( .A1(n868), .A2(n820), .ZN(n1011) );
  NAND2_X1 U915 ( .A1(n821), .A2(n1011), .ZN(n822) );
  XNOR2_X1 U916 ( .A(KEYINPUT108), .B(n822), .ZN(n824) );
  NAND2_X1 U917 ( .A1(n824), .A2(n823), .ZN(n825) );
  NAND2_X1 U918 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U919 ( .A(n827), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U920 ( .A(G301), .ZN(G171) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n828), .ZN(G217) );
  AND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n829) );
  NAND2_X1 U923 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G3), .A2(G1), .ZN(n830) );
  XOR2_X1 U925 ( .A(KEYINPUT113), .B(n830), .Z(n831) );
  NAND2_X1 U926 ( .A1(n832), .A2(n831), .ZN(G188) );
  XNOR2_X1 U927 ( .A(G108), .B(KEYINPUT119), .ZN(G238) );
  INV_X1 U929 ( .A(G120), .ZN(G236) );
  INV_X1 U930 ( .A(G96), .ZN(G221) );
  NOR2_X1 U931 ( .A1(n834), .A2(n833), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  INV_X1 U933 ( .A(n835), .ZN(G319) );
  XOR2_X1 U934 ( .A(G2100), .B(G2096), .Z(n837) );
  XNOR2_X1 U935 ( .A(KEYINPUT42), .B(G2678), .ZN(n836) );
  XNOR2_X1 U936 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U937 ( .A(KEYINPUT43), .B(G2090), .Z(n839) );
  XNOR2_X1 U938 ( .A(G2067), .B(G2072), .ZN(n838) );
  XNOR2_X1 U939 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U940 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U941 ( .A(G2084), .B(G2078), .ZN(n842) );
  XNOR2_X1 U942 ( .A(n843), .B(n842), .ZN(G227) );
  XOR2_X1 U943 ( .A(G1961), .B(G1966), .Z(n845) );
  XNOR2_X1 U944 ( .A(G1981), .B(G1971), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U946 ( .A(n846), .B(KEYINPUT41), .Z(n848) );
  XNOR2_X1 U947 ( .A(G1996), .B(G1991), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U949 ( .A(G2474), .B(G1956), .Z(n850) );
  XNOR2_X1 U950 ( .A(G1986), .B(G1976), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n852), .B(n851), .ZN(G229) );
  NAND2_X1 U953 ( .A1(n880), .A2(G124), .ZN(n853) );
  XNOR2_X1 U954 ( .A(n853), .B(KEYINPUT44), .ZN(n855) );
  NAND2_X1 U955 ( .A1(G136), .A2(n889), .ZN(n854) );
  NAND2_X1 U956 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U957 ( .A(KEYINPUT114), .B(n856), .ZN(n860) );
  NAND2_X1 U958 ( .A1(G100), .A2(n886), .ZN(n858) );
  NAND2_X1 U959 ( .A1(G112), .A2(n882), .ZN(n857) );
  NAND2_X1 U960 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U961 ( .A1(n860), .A2(n859), .ZN(G162) );
  XOR2_X1 U962 ( .A(G164), .B(G162), .Z(n861) );
  XNOR2_X1 U963 ( .A(n862), .B(n861), .ZN(n867) );
  XNOR2_X1 U964 ( .A(KEYINPUT48), .B(KEYINPUT118), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n863), .B(KEYINPUT46), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n865), .B(n864), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n867), .B(n866), .ZN(n870) );
  XNOR2_X1 U968 ( .A(n868), .B(n1008), .ZN(n869) );
  XNOR2_X1 U969 ( .A(n870), .B(n869), .ZN(n879) );
  NAND2_X1 U970 ( .A1(G118), .A2(n882), .ZN(n872) );
  NAND2_X1 U971 ( .A1(G130), .A2(n880), .ZN(n871) );
  NAND2_X1 U972 ( .A1(n872), .A2(n871), .ZN(n877) );
  NAND2_X1 U973 ( .A1(G142), .A2(n889), .ZN(n874) );
  NAND2_X1 U974 ( .A1(G106), .A2(n886), .ZN(n873) );
  NAND2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U976 ( .A(KEYINPUT45), .B(n875), .Z(n876) );
  NOR2_X1 U977 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U978 ( .A(n879), .B(n878), .Z(n895) );
  NAND2_X1 U979 ( .A1(n880), .A2(G127), .ZN(n881) );
  XNOR2_X1 U980 ( .A(n881), .B(KEYINPUT116), .ZN(n884) );
  NAND2_X1 U981 ( .A1(G115), .A2(n882), .ZN(n883) );
  NAND2_X1 U982 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U983 ( .A(n885), .B(KEYINPUT47), .ZN(n888) );
  NAND2_X1 U984 ( .A1(G103), .A2(n886), .ZN(n887) );
  NAND2_X1 U985 ( .A1(n888), .A2(n887), .ZN(n892) );
  NAND2_X1 U986 ( .A1(G139), .A2(n889), .ZN(n890) );
  XNOR2_X1 U987 ( .A(KEYINPUT115), .B(n890), .ZN(n891) );
  NOR2_X1 U988 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U989 ( .A(KEYINPUT117), .B(n893), .Z(n1003) );
  XNOR2_X1 U990 ( .A(G160), .B(n1003), .ZN(n894) );
  XNOR2_X1 U991 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U992 ( .A1(G37), .A2(n896), .ZN(G395) );
  XOR2_X1 U993 ( .A(n897), .B(G286), .Z(n900) );
  XNOR2_X1 U994 ( .A(G301), .B(n898), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U996 ( .A(n901), .B(n954), .ZN(n902) );
  NOR2_X1 U997 ( .A1(G37), .A2(n902), .ZN(G397) );
  XOR2_X1 U998 ( .A(G2427), .B(KEYINPUT112), .Z(n904) );
  XNOR2_X1 U999 ( .A(G1341), .B(G1348), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(n904), .B(n903), .ZN(n914) );
  XOR2_X1 U1001 ( .A(G2451), .B(KEYINPUT111), .Z(n906) );
  XNOR2_X1 U1002 ( .A(G2430), .B(G2435), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(n906), .B(n905), .ZN(n910) );
  XOR2_X1 U1004 ( .A(G2438), .B(KEYINPUT110), .Z(n908) );
  XNOR2_X1 U1005 ( .A(G2443), .B(G2454), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1007 ( .A(n910), .B(n909), .Z(n912) );
  XNOR2_X1 U1008 ( .A(G2446), .B(KEYINPUT109), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n912), .B(n911), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(n914), .B(n913), .ZN(n915) );
  NAND2_X1 U1011 ( .A1(n915), .A2(G14), .ZN(n921) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n921), .ZN(n918) );
  NOR2_X1 U1013 ( .A1(G227), .A2(G229), .ZN(n916) );
  XNOR2_X1 U1014 ( .A(KEYINPUT49), .B(n916), .ZN(n917) );
  NOR2_X1 U1015 ( .A1(n918), .A2(n917), .ZN(n920) );
  NOR2_X1 U1016 ( .A1(G395), .A2(G397), .ZN(n919) );
  NAND2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(G69), .ZN(G235) );
  INV_X1 U1020 ( .A(n921), .ZN(G401) );
  INV_X1 U1021 ( .A(KEYINPUT55), .ZN(n1027) );
  XNOR2_X1 U1022 ( .A(G2090), .B(G35), .ZN(n935) );
  XOR2_X1 U1023 ( .A(G1991), .B(G25), .Z(n922) );
  NAND2_X1 U1024 ( .A1(n922), .A2(G28), .ZN(n932) );
  XNOR2_X1 U1025 ( .A(G2067), .B(G26), .ZN(n924) );
  XNOR2_X1 U1026 ( .A(G33), .B(G2072), .ZN(n923) );
  NOR2_X1 U1027 ( .A1(n924), .A2(n923), .ZN(n930) );
  XOR2_X1 U1028 ( .A(n925), .B(G27), .Z(n928) );
  INV_X1 U1029 ( .A(G1996), .ZN(n926) );
  XOR2_X1 U1030 ( .A(n926), .B(G32), .Z(n927) );
  NOR2_X1 U1031 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1032 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1033 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1034 ( .A(KEYINPUT53), .B(n933), .ZN(n934) );
  NOR2_X1 U1035 ( .A1(n935), .A2(n934), .ZN(n938) );
  XOR2_X1 U1036 ( .A(G2084), .B(G34), .Z(n936) );
  XNOR2_X1 U1037 ( .A(KEYINPUT54), .B(n936), .ZN(n937) );
  NAND2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1039 ( .A(n1027), .B(n939), .ZN(n941) );
  INV_X1 U1040 ( .A(G29), .ZN(n940) );
  NAND2_X1 U1041 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1042 ( .A1(G11), .A2(n942), .ZN(n1001) );
  XNOR2_X1 U1043 ( .A(G16), .B(KEYINPUT56), .ZN(n970) );
  XNOR2_X1 U1044 ( .A(G1961), .B(G171), .ZN(n953) );
  XNOR2_X1 U1045 ( .A(G1956), .B(n943), .ZN(n945) );
  NAND2_X1 U1046 ( .A1(G1971), .A2(G303), .ZN(n944) );
  NAND2_X1 U1047 ( .A1(n945), .A2(n944), .ZN(n951) );
  INV_X1 U1048 ( .A(n946), .ZN(n948) );
  NAND2_X1 U1049 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1050 ( .A(KEYINPUT123), .B(n949), .Z(n950) );
  NOR2_X1 U1051 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1052 ( .A1(n953), .A2(n952), .ZN(n956) );
  XNOR2_X1 U1053 ( .A(G1341), .B(n954), .ZN(n955) );
  NOR2_X1 U1054 ( .A1(n956), .A2(n955), .ZN(n968) );
  XNOR2_X1 U1055 ( .A(G1348), .B(n957), .ZN(n958) );
  NOR2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(G1966), .B(G168), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1060 ( .A(KEYINPUT57), .B(n964), .Z(n965) );
  NOR2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n999) );
  INV_X1 U1064 ( .A(G16), .ZN(n997) );
  XNOR2_X1 U1065 ( .A(G1966), .B(G21), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(G1961), .B(G5), .ZN(n971) );
  NOR2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n985) );
  XOR2_X1 U1068 ( .A(G1341), .B(G19), .Z(n977) );
  XOR2_X1 U1069 ( .A(KEYINPUT125), .B(G4), .Z(n974) );
  XNOR2_X1 U1070 ( .A(G1348), .B(KEYINPUT59), .ZN(n973) );
  XNOR2_X1 U1071 ( .A(n974), .B(n973), .ZN(n975) );
  XNOR2_X1 U1072 ( .A(KEYINPUT124), .B(n975), .ZN(n976) );
  NAND2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n982) );
  XOR2_X1 U1074 ( .A(G1981), .B(G6), .Z(n980) );
  XNOR2_X1 U1075 ( .A(n978), .B(G20), .ZN(n979) );
  NAND2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1078 ( .A(n983), .B(KEYINPUT60), .ZN(n984) );
  NAND2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n993) );
  XNOR2_X1 U1080 ( .A(G1986), .B(G24), .ZN(n987) );
  XNOR2_X1 U1081 ( .A(G1971), .B(G22), .ZN(n986) );
  NOR2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n990) );
  XOR2_X1 U1083 ( .A(G1976), .B(KEYINPUT126), .Z(n988) );
  XNOR2_X1 U1084 ( .A(G23), .B(n988), .ZN(n989) );
  NAND2_X1 U1085 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1086 ( .A(KEYINPUT58), .B(n991), .ZN(n992) );
  NOR2_X1 U1087 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1088 ( .A(n994), .B(KEYINPUT61), .Z(n995) );
  XNOR2_X1 U1089 ( .A(KEYINPUT127), .B(n995), .ZN(n996) );
  NAND2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1031) );
  XOR2_X1 U1093 ( .A(G164), .B(G2078), .Z(n1002) );
  XNOR2_X1 U1094 ( .A(KEYINPUT122), .B(n1002), .ZN(n1005) );
  XOR2_X1 U1095 ( .A(G2072), .B(n1003), .Z(n1004) );
  NOR2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1097 ( .A(KEYINPUT50), .B(n1006), .ZN(n1023) );
  XNOR2_X1 U1098 ( .A(G160), .B(G2084), .ZN(n1015) );
  NOR2_X1 U1099 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1100 ( .A(n1009), .B(KEYINPUT120), .ZN(n1010) );
  NAND2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1021) );
  XNOR2_X1 U1104 ( .A(G2090), .B(G162), .ZN(n1016) );
  XNOR2_X1 U1105 ( .A(n1016), .B(KEYINPUT121), .ZN(n1018) );
  NOR2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(KEYINPUT51), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1111 ( .A(KEYINPUT52), .B(n1026), .ZN(n1028) );
  NAND2_X1 U1112 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1113 ( .A1(n1029), .A2(G29), .ZN(n1030) );
  NAND2_X1 U1114 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1032), .Z(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

