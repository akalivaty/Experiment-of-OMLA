

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758;

  XNOR2_X1 U366 ( .A(n393), .B(n539), .ZN(n676) );
  AND2_X1 U367 ( .A1(n400), .A2(n559), .ZN(n612) );
  XNOR2_X1 U368 ( .A(n418), .B(KEYINPUT31), .ZN(n680) );
  XNOR2_X1 U369 ( .A(n561), .B(KEYINPUT114), .ZN(n421) );
  NAND2_X1 U370 ( .A1(n557), .A2(n695), .ZN(n690) );
  XNOR2_X1 U371 ( .A(G902), .B(KEYINPUT15), .ZN(n626) );
  XNOR2_X1 U372 ( .A(n641), .B(KEYINPUT62), .ZN(n642) );
  NOR2_X2 U373 ( .A1(n623), .A2(n441), .ZN(n430) );
  XNOR2_X1 U374 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U375 ( .A(n504), .B(G134), .ZN(n533) );
  XNOR2_X1 U376 ( .A(n490), .B(n489), .ZN(n510) );
  XOR2_X1 U377 ( .A(KEYINPUT3), .B(G101), .Z(n489) );
  INV_X1 U378 ( .A(G119), .ZN(n487) );
  XNOR2_X1 U379 ( .A(n430), .B(KEYINPUT22), .ZN(n356) );
  XNOR2_X1 U380 ( .A(n392), .B(n584), .ZN(n585) );
  AND2_X1 U381 ( .A1(n390), .A2(n587), .ZN(n389) );
  NOR2_X1 U382 ( .A1(G902), .A2(G237), .ZN(n498) );
  INV_X1 U383 ( .A(KEYINPUT48), .ZN(n600) );
  NOR2_X1 U384 ( .A1(n597), .A2(n683), .ZN(n598) );
  INV_X1 U385 ( .A(n667), .ZN(n416) );
  AND2_X1 U386 ( .A1(n399), .A2(n395), .ZN(n614) );
  XNOR2_X1 U387 ( .A(n431), .B(n453), .ZN(n407) );
  OR2_X1 U388 ( .A1(n637), .A2(n452), .ZN(n431) );
  XNOR2_X1 U389 ( .A(n533), .B(n443), .ZN(n747) );
  XNOR2_X1 U390 ( .A(G131), .B(G137), .ZN(n442) );
  INV_X1 U391 ( .A(KEYINPUT115), .ZN(n563) );
  NAND2_X1 U392 ( .A1(n707), .A2(n351), .ZN(n379) );
  NAND2_X1 U393 ( .A1(G214), .A2(n512), .ZN(n704) );
  OR2_X1 U394 ( .A1(n655), .A2(G902), .ZN(n451) );
  NAND2_X1 U395 ( .A1(n362), .A2(n353), .ZN(n361) );
  NAND2_X1 U396 ( .A1(n438), .A2(n436), .ZN(n435) );
  NAND2_X1 U397 ( .A1(n629), .A2(n437), .ZN(n436) );
  NAND2_X1 U398 ( .A1(n439), .A2(KEYINPUT65), .ZN(n438) );
  NAND2_X1 U399 ( .A1(n626), .A2(KEYINPUT65), .ZN(n437) );
  OR2_X1 U400 ( .A1(n637), .A2(n444), .ZN(n446) );
  XNOR2_X1 U401 ( .A(n747), .B(G146), .ZN(n495) );
  XNOR2_X1 U402 ( .A(n511), .B(n733), .ZN(n647) );
  INV_X1 U403 ( .A(n609), .ZN(n355) );
  XNOR2_X1 U404 ( .A(n424), .B(n423), .ZN(n732) );
  INV_X1 U405 ( .A(G107), .ZN(n423) );
  XNOR2_X1 U406 ( .A(G104), .B(G110), .ZN(n424) );
  XNOR2_X1 U407 ( .A(n388), .B(n387), .ZN(n597) );
  INV_X1 U408 ( .A(KEYINPUT75), .ZN(n387) );
  INV_X1 U409 ( .A(n680), .ZN(n417) );
  XOR2_X1 U410 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n518) );
  NOR2_X1 U411 ( .A1(G237), .A2(G953), .ZN(n491) );
  XNOR2_X1 U412 ( .A(G116), .B(G113), .ZN(n488) );
  XOR2_X1 U413 ( .A(G104), .B(G122), .Z(n522) );
  XNOR2_X1 U414 ( .A(G113), .B(G143), .ZN(n521) );
  NAND2_X1 U415 ( .A1(G234), .A2(G237), .ZN(n477) );
  INV_X1 U416 ( .A(n705), .ZN(n434) );
  XNOR2_X1 U417 ( .A(n420), .B(KEYINPUT78), .ZN(n621) );
  NOR2_X1 U418 ( .A1(n691), .A2(n690), .ZN(n420) );
  AND2_X1 U419 ( .A1(n375), .A2(n374), .ZN(n373) );
  NOR2_X1 U420 ( .A1(n690), .A2(KEYINPUT111), .ZN(n372) );
  INV_X1 U421 ( .A(G902), .ZN(n535) );
  AND2_X1 U422 ( .A1(n758), .A2(n350), .ZN(n409) );
  XNOR2_X1 U423 ( .A(KEYINPUT24), .B(KEYINPUT71), .ZN(n462) );
  XNOR2_X1 U424 ( .A(KEYINPUT93), .B(KEYINPUT94), .ZN(n463) );
  XNOR2_X1 U425 ( .A(G140), .B(KEYINPUT10), .ZN(n461) );
  NAND2_X1 U426 ( .A1(n378), .A2(n377), .ZN(n376) );
  AND2_X1 U427 ( .A1(n380), .A2(n379), .ZN(n364) );
  XNOR2_X1 U428 ( .A(n541), .B(KEYINPUT19), .ZN(n542) );
  NAND2_X1 U429 ( .A1(n589), .A2(n704), .ZN(n405) );
  XNOR2_X1 U430 ( .A(n508), .B(G122), .ZN(n509) );
  XOR2_X1 U431 ( .A(KEYINPUT74), .B(KEYINPUT16), .Z(n508) );
  AND2_X1 U432 ( .A1(n361), .A2(n435), .ZN(n360) );
  XNOR2_X1 U433 ( .A(n385), .B(n384), .ZN(n727) );
  XNOR2_X1 U434 ( .A(n347), .B(n532), .ZN(n384) );
  XNOR2_X1 U435 ( .A(n386), .B(n534), .ZN(n385) );
  AND2_X1 U436 ( .A1(n637), .A2(n636), .ZN(n731) );
  XNOR2_X1 U437 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U438 ( .A(G101), .B(G140), .ZN(n445) );
  INV_X1 U439 ( .A(G953), .ZN(n736) );
  XNOR2_X1 U440 ( .A(n572), .B(n422), .ZN(n573) );
  INV_X1 U441 ( .A(KEYINPUT42), .ZN(n422) );
  NOR2_X1 U442 ( .A1(n719), .A2(n581), .ZN(n572) );
  XNOR2_X1 U443 ( .A(n413), .B(n352), .ZN(n574) );
  XNOR2_X1 U444 ( .A(n396), .B(KEYINPUT35), .ZN(n613) );
  NAND2_X1 U445 ( .A1(n397), .A2(n588), .ZN(n396) );
  XNOR2_X1 U446 ( .A(n404), .B(n398), .ZN(n397) );
  INV_X1 U447 ( .A(KEYINPUT34), .ZN(n398) );
  XNOR2_X1 U448 ( .A(n401), .B(n611), .ZN(n757) );
  NAND2_X1 U449 ( .A1(n619), .A2(n346), .ZN(n620) );
  XNOR2_X1 U450 ( .A(n573), .B(G137), .ZN(G39) );
  AND2_X1 U451 ( .A1(n371), .A2(n369), .ZN(n346) );
  XOR2_X1 U452 ( .A(n529), .B(n528), .Z(n347) );
  AND2_X1 U453 ( .A1(n685), .A2(KEYINPUT87), .ZN(n348) );
  XNOR2_X1 U454 ( .A(n527), .B(n526), .ZN(n555) );
  AND2_X2 U455 ( .A1(n686), .A2(n358), .ZN(n662) );
  XOR2_X1 U456 ( .A(n513), .B(KEYINPUT85), .Z(n349) );
  OR2_X1 U457 ( .A1(n685), .A2(KEYINPUT87), .ZN(n350) );
  INV_X1 U458 ( .A(n392), .ZN(n708) );
  OR2_X1 U459 ( .A1(n676), .A2(n679), .ZN(n392) );
  XOR2_X1 U460 ( .A(n563), .B(KEYINPUT41), .Z(n351) );
  XOR2_X1 U461 ( .A(KEYINPUT113), .B(KEYINPUT40), .Z(n352) );
  AND2_X1 U462 ( .A1(n629), .A2(KEYINPUT65), .ZN(n353) );
  AND2_X1 U463 ( .A1(n627), .A2(n630), .ZN(n354) );
  AND2_X2 U464 ( .A1(n356), .A2(n355), .ZN(n615) );
  AND2_X1 U465 ( .A1(n356), .A2(n691), .ZN(n556) );
  AND2_X2 U466 ( .A1(n414), .A2(KEYINPUT2), .ZN(n357) );
  NAND2_X1 U467 ( .A1(n748), .A2(n414), .ZN(n362) );
  INV_X1 U468 ( .A(n362), .ZN(n687) );
  NAND2_X1 U469 ( .A1(n357), .A2(n748), .ZN(n363) );
  NAND2_X1 U470 ( .A1(n360), .A2(n359), .ZN(n358) );
  NAND2_X1 U471 ( .A1(n687), .A2(n354), .ZN(n359) );
  XNOR2_X2 U472 ( .A(n363), .B(n631), .ZN(n686) );
  NAND2_X1 U473 ( .A1(n364), .A2(n376), .ZN(n719) );
  NAND2_X1 U474 ( .A1(n573), .A2(n574), .ZN(n576) );
  XNOR2_X1 U475 ( .A(n365), .B(n517), .ZN(n519) );
  XNOR2_X1 U476 ( .A(n518), .B(n516), .ZN(n365) );
  NAND2_X1 U477 ( .A1(n555), .A2(n394), .ZN(n393) );
  XNOR2_X2 U478 ( .A(G143), .B(G128), .ZN(n504) );
  NAND2_X1 U479 ( .A1(n501), .A2(n500), .ZN(n368) );
  AND2_X1 U480 ( .A1(n366), .A2(n501), .ZN(n433) );
  NOR2_X1 U481 ( .A1(n367), .A2(n434), .ZN(n366) );
  INV_X1 U482 ( .A(n500), .ZN(n367) );
  NOR2_X1 U483 ( .A1(n368), .A2(n590), .ZN(n673) );
  NAND2_X1 U484 ( .A1(n690), .A2(KEYINPUT111), .ZN(n374) );
  NAND2_X1 U485 ( .A1(n570), .A2(KEYINPUT111), .ZN(n375) );
  INV_X1 U486 ( .A(n690), .ZN(n369) );
  NAND2_X1 U487 ( .A1(n373), .A2(n370), .ZN(n484) );
  NAND2_X1 U488 ( .A1(n372), .A2(n371), .ZN(n370) );
  INV_X1 U489 ( .A(n570), .ZN(n371) );
  NOR2_X1 U490 ( .A1(n707), .A2(n351), .ZN(n377) );
  INV_X1 U491 ( .A(n421), .ZN(n378) );
  NAND2_X1 U492 ( .A1(n421), .A2(n351), .ZN(n380) );
  XNOR2_X1 U493 ( .A(n381), .B(KEYINPUT107), .ZN(n624) );
  NAND2_X1 U494 ( .A1(n402), .A2(n382), .ZN(n381) );
  NAND2_X1 U495 ( .A1(n415), .A2(n392), .ZN(n382) );
  XNOR2_X2 U496 ( .A(n383), .B(KEYINPUT106), .ZN(n402) );
  NAND2_X1 U497 ( .A1(n618), .A2(n617), .ZN(n383) );
  NAND2_X1 U498 ( .A1(n727), .A2(n535), .ZN(n538) );
  NAND2_X1 U499 ( .A1(n407), .A2(G217), .ZN(n386) );
  NAND2_X1 U500 ( .A1(n391), .A2(n389), .ZN(n388) );
  INV_X1 U501 ( .A(n673), .ZN(n390) );
  NAND2_X1 U502 ( .A1(n586), .A2(n674), .ZN(n391) );
  INV_X1 U503 ( .A(n577), .ZN(n394) );
  INV_X1 U504 ( .A(n613), .ZN(n395) );
  NOR2_X1 U505 ( .A1(n757), .A2(n612), .ZN(n399) );
  XNOR2_X1 U506 ( .A(n556), .B(KEYINPUT108), .ZN(n400) );
  NAND2_X1 U507 ( .A1(n615), .A2(n610), .ZN(n401) );
  XNOR2_X1 U508 ( .A(n402), .B(G101), .ZN(G3) );
  XNOR2_X2 U509 ( .A(n403), .B(KEYINPUT45), .ZN(n414) );
  NAND2_X1 U510 ( .A1(n624), .A2(n625), .ZN(n403) );
  NAND2_X1 U511 ( .A1(n711), .A2(n554), .ZN(n404) );
  XNOR2_X2 U512 ( .A(n405), .B(n542), .ZN(n579) );
  XNOR2_X2 U513 ( .A(n406), .B(KEYINPUT0), .ZN(n623) );
  NAND2_X1 U514 ( .A1(n579), .A2(n548), .ZN(n406) );
  NAND2_X1 U515 ( .A1(n407), .A2(G221), .ZN(n460) );
  XNOR2_X2 U516 ( .A(n440), .B(n472), .ZN(n557) );
  NOR2_X2 U517 ( .A1(n411), .A2(n408), .ZN(n748) );
  NAND2_X1 U518 ( .A1(n410), .A2(n409), .ZN(n408) );
  NAND2_X1 U519 ( .A1(n412), .A2(n348), .ZN(n410) );
  NOR2_X1 U520 ( .A1(n412), .A2(KEYINPUT87), .ZN(n411) );
  XNOR2_X1 U521 ( .A(n601), .B(n600), .ZN(n412) );
  INV_X1 U522 ( .A(n574), .ZN(n560) );
  NAND2_X1 U523 ( .A1(n607), .A2(n676), .ZN(n413) );
  XNOR2_X1 U524 ( .A(n433), .B(n432), .ZN(n607) );
  NAND2_X1 U525 ( .A1(n414), .A2(n736), .ZN(n741) );
  INV_X1 U526 ( .A(n637), .ZN(n749) );
  XNOR2_X2 U527 ( .A(G953), .B(KEYINPUT64), .ZN(n637) );
  NOR2_X1 U528 ( .A1(n637), .A2(n429), .ZN(n428) );
  NAND2_X1 U529 ( .A1(n417), .A2(n416), .ZN(n415) );
  NAND2_X1 U530 ( .A1(n419), .A2(n554), .ZN(n418) );
  INV_X1 U531 ( .A(n700), .ZN(n419) );
  NAND2_X1 U532 ( .A1(n621), .A2(n694), .ZN(n622) );
  XNOR2_X2 U533 ( .A(n570), .B(n549), .ZN(n691) );
  NOR2_X1 U534 ( .A1(n421), .A2(n708), .ZN(n709) );
  XNOR2_X1 U535 ( .A(n425), .B(n505), .ZN(n507) );
  XNOR2_X1 U536 ( .A(n428), .B(n426), .ZN(n425) );
  XNOR2_X1 U537 ( .A(n502), .B(n427), .ZN(n426) );
  XNOR2_X2 U538 ( .A(KEYINPUT4), .B(KEYINPUT18), .ZN(n427) );
  INV_X1 U539 ( .A(G224), .ZN(n429) );
  INV_X1 U540 ( .A(n540), .ZN(n589) );
  INV_X1 U541 ( .A(KEYINPUT39), .ZN(n432) );
  INV_X1 U542 ( .A(n629), .ZN(n439) );
  INV_X1 U543 ( .A(n557), .ZN(n564) );
  NAND2_X1 U544 ( .A1(n661), .A2(n535), .ZN(n440) );
  XNOR2_X1 U545 ( .A(n486), .B(n485), .ZN(n501) );
  NAND2_X1 U546 ( .A1(n562), .A2(n695), .ZN(n441) );
  INV_X1 U547 ( .A(KEYINPUT5), .ZN(n492) );
  XNOR2_X1 U548 ( .A(n493), .B(n492), .ZN(n494) );
  INV_X1 U549 ( .A(KEYINPUT83), .ZN(n541) );
  XNOR2_X1 U550 ( .A(n488), .B(n487), .ZN(n490) );
  INV_X1 U551 ( .A(KEYINPUT82), .ZN(n485) );
  XNOR2_X1 U552 ( .A(n442), .B(KEYINPUT4), .ZN(n443) );
  XNOR2_X1 U553 ( .A(n732), .B(KEYINPUT72), .ZN(n506) );
  INV_X1 U554 ( .A(G227), .ZN(n444) );
  XNOR2_X1 U555 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U556 ( .A(n506), .B(n447), .ZN(n448) );
  XNOR2_X1 U557 ( .A(n495), .B(n448), .ZN(n655) );
  INV_X1 U558 ( .A(KEYINPUT70), .ZN(n449) );
  XNOR2_X1 U559 ( .A(n449), .B(G469), .ZN(n450) );
  XNOR2_X2 U560 ( .A(n451), .B(n450), .ZN(n570) );
  INV_X1 U561 ( .A(G234), .ZN(n452) );
  XOR2_X1 U562 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n453) );
  XNOR2_X1 U563 ( .A(G110), .B(KEYINPUT95), .ZN(n455) );
  XNOR2_X1 U564 ( .A(KEYINPUT23), .B(G119), .ZN(n454) );
  XNOR2_X1 U565 ( .A(n455), .B(n454), .ZN(n458) );
  XNOR2_X1 U566 ( .A(G128), .B(G137), .ZN(n456) );
  XNOR2_X1 U567 ( .A(n456), .B(KEYINPUT86), .ZN(n457) );
  XNOR2_X1 U568 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U569 ( .A(n460), .B(n459), .ZN(n466) );
  XNOR2_X1 U570 ( .A(G146), .B(G125), .ZN(n503) );
  XNOR2_X1 U571 ( .A(n503), .B(n461), .ZN(n745) );
  XNOR2_X1 U572 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U573 ( .A(n745), .B(n464), .ZN(n465) );
  XNOR2_X1 U574 ( .A(n466), .B(n465), .ZN(n661) );
  NAND2_X1 U575 ( .A1(n626), .A2(G234), .ZN(n468) );
  INV_X1 U576 ( .A(KEYINPUT20), .ZN(n467) );
  XNOR2_X1 U577 ( .A(n468), .B(n467), .ZN(n474) );
  INV_X1 U578 ( .A(G217), .ZN(n469) );
  OR2_X1 U579 ( .A1(n474), .A2(n469), .ZN(n471) );
  INV_X1 U580 ( .A(KEYINPUT25), .ZN(n470) );
  XNOR2_X1 U581 ( .A(n471), .B(n470), .ZN(n472) );
  INV_X1 U582 ( .A(G221), .ZN(n473) );
  OR2_X1 U583 ( .A1(n474), .A2(n473), .ZN(n476) );
  INV_X1 U584 ( .A(KEYINPUT21), .ZN(n475) );
  XNOR2_X1 U585 ( .A(n476), .B(n475), .ZN(n695) );
  XOR2_X1 U586 ( .A(KEYINPUT77), .B(KEYINPUT14), .Z(n478) );
  XNOR2_X1 U587 ( .A(n478), .B(n477), .ZN(n481) );
  NAND2_X1 U588 ( .A1(n481), .A2(G952), .ZN(n479) );
  XNOR2_X1 U589 ( .A(n479), .B(KEYINPUT90), .ZN(n717) );
  NOR2_X1 U590 ( .A1(G953), .A2(n717), .ZN(n480) );
  XNOR2_X1 U591 ( .A(n480), .B(KEYINPUT91), .ZN(n547) );
  NAND2_X1 U592 ( .A1(G902), .A2(n481), .ZN(n543) );
  NOR2_X1 U593 ( .A1(G900), .A2(n543), .ZN(n482) );
  NAND2_X1 U594 ( .A1(n482), .A2(n637), .ZN(n483) );
  NAND2_X1 U595 ( .A1(n547), .A2(n483), .ZN(n565) );
  NAND2_X1 U596 ( .A1(n484), .A2(n565), .ZN(n486) );
  XNOR2_X1 U597 ( .A(n491), .B(KEYINPUT80), .ZN(n515) );
  NAND2_X1 U598 ( .A1(G210), .A2(n515), .ZN(n493) );
  XNOR2_X1 U599 ( .A(n510), .B(n494), .ZN(n496) );
  XNOR2_X1 U600 ( .A(n496), .B(n495), .ZN(n641) );
  NAND2_X1 U601 ( .A1(n641), .A2(n535), .ZN(n497) );
  XNOR2_X2 U602 ( .A(n497), .B(G472), .ZN(n694) );
  XNOR2_X1 U603 ( .A(n498), .B(KEYINPUT79), .ZN(n512) );
  NAND2_X1 U604 ( .A1(n694), .A2(n704), .ZN(n499) );
  XOR2_X1 U605 ( .A(KEYINPUT30), .B(n499), .Z(n500) );
  XNOR2_X2 U606 ( .A(KEYINPUT84), .B(KEYINPUT17), .ZN(n502) );
  XNOR2_X1 U607 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U608 ( .A(n507), .B(n506), .ZN(n511) );
  XNOR2_X1 U609 ( .A(n510), .B(n509), .ZN(n733) );
  NAND2_X1 U610 ( .A1(n647), .A2(n626), .ZN(n514) );
  NAND2_X1 U611 ( .A1(G210), .A2(n512), .ZN(n513) );
  XNOR2_X2 U612 ( .A(n514), .B(n349), .ZN(n540) );
  BUF_X2 U613 ( .A(n540), .Z(n605) );
  XNOR2_X2 U614 ( .A(n605), .B(KEYINPUT38), .ZN(n705) );
  AND2_X1 U615 ( .A1(n515), .A2(G214), .ZN(n520) );
  XOR2_X1 U616 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n517) );
  XNOR2_X1 U617 ( .A(G131), .B(KEYINPUT97), .ZN(n516) );
  XNOR2_X1 U618 ( .A(n520), .B(n519), .ZN(n525) );
  XNOR2_X1 U619 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U620 ( .A(n745), .B(n523), .ZN(n524) );
  XNOR2_X1 U621 ( .A(n525), .B(n524), .ZN(n633) );
  NAND2_X1 U622 ( .A1(n633), .A2(n535), .ZN(n527) );
  XOR2_X1 U623 ( .A(KEYINPUT13), .B(G475), .Z(n526) );
  INV_X1 U624 ( .A(n555), .ZN(n578) );
  XOR2_X1 U625 ( .A(KEYINPUT102), .B(G107), .Z(n529) );
  XNOR2_X1 U626 ( .A(G116), .B(G122), .ZN(n528) );
  XOR2_X1 U627 ( .A(KEYINPUT7), .B(KEYINPUT100), .Z(n531) );
  XNOR2_X1 U628 ( .A(KEYINPUT101), .B(KEYINPUT9), .ZN(n530) );
  XNOR2_X1 U629 ( .A(n531), .B(n530), .ZN(n532) );
  INV_X1 U630 ( .A(n533), .ZN(n534) );
  INV_X1 U631 ( .A(KEYINPUT103), .ZN(n536) );
  XNOR2_X1 U632 ( .A(n536), .B(G478), .ZN(n537) );
  XNOR2_X1 U633 ( .A(n538), .B(n537), .ZN(n577) );
  INV_X1 U634 ( .A(KEYINPUT104), .ZN(n539) );
  XOR2_X1 U635 ( .A(n560), .B(G131), .Z(G33) );
  INV_X1 U636 ( .A(n543), .ZN(n544) );
  NOR2_X1 U637 ( .A1(G898), .A2(n736), .ZN(n735) );
  NAND2_X1 U638 ( .A1(n544), .A2(n735), .ZN(n545) );
  XNOR2_X1 U639 ( .A(KEYINPUT92), .B(n545), .ZN(n546) );
  NAND2_X1 U640 ( .A1(n547), .A2(n546), .ZN(n548) );
  INV_X1 U641 ( .A(n623), .ZN(n554) );
  XNOR2_X1 U642 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n549) );
  XNOR2_X1 U643 ( .A(KEYINPUT105), .B(KEYINPUT6), .ZN(n550) );
  XNOR2_X1 U644 ( .A(n694), .B(n550), .ZN(n609) );
  NAND2_X1 U645 ( .A1(n621), .A2(n609), .ZN(n553) );
  XNOR2_X1 U646 ( .A(KEYINPUT109), .B(KEYINPUT33), .ZN(n551) );
  XNOR2_X1 U647 ( .A(n551), .B(KEYINPUT73), .ZN(n552) );
  XNOR2_X1 U648 ( .A(n553), .B(n552), .ZN(n711) );
  AND2_X1 U649 ( .A1(n577), .A2(n555), .ZN(n588) );
  XOR2_X1 U650 ( .A(G122), .B(n613), .Z(G24) );
  NOR2_X1 U651 ( .A1(n555), .A2(n577), .ZN(n562) );
  INV_X1 U652 ( .A(n691), .ZN(n616) );
  BUF_X1 U653 ( .A(n557), .Z(n558) );
  NOR2_X1 U654 ( .A1(n694), .A2(n558), .ZN(n559) );
  XOR2_X1 U655 ( .A(G110), .B(n612), .Z(G12) );
  NAND2_X1 U656 ( .A1(n705), .A2(n704), .ZN(n561) );
  INV_X1 U657 ( .A(n562), .ZN(n707) );
  NAND2_X1 U658 ( .A1(n565), .A2(n695), .ZN(n566) );
  XNOR2_X1 U659 ( .A(KEYINPUT69), .B(n566), .ZN(n567) );
  AND2_X1 U660 ( .A1(n564), .A2(n567), .ZN(n591) );
  NAND2_X1 U661 ( .A1(n694), .A2(n591), .ZN(n569) );
  XOR2_X1 U662 ( .A(KEYINPUT28), .B(KEYINPUT112), .Z(n568) );
  XNOR2_X1 U663 ( .A(n569), .B(n568), .ZN(n571) );
  NAND2_X1 U664 ( .A1(n571), .A2(n371), .ZN(n581) );
  INV_X1 U665 ( .A(KEYINPUT46), .ZN(n575) );
  XNOR2_X1 U666 ( .A(n576), .B(n575), .ZN(n599) );
  AND2_X1 U667 ( .A1(n578), .A2(n577), .ZN(n679) );
  INV_X1 U668 ( .A(KEYINPUT76), .ZN(n584) );
  NOR2_X1 U669 ( .A1(n708), .A2(n584), .ZN(n582) );
  INV_X1 U670 ( .A(n579), .ZN(n580) );
  NOR2_X1 U671 ( .A1(n581), .A2(n580), .ZN(n674) );
  NAND2_X1 U672 ( .A1(n582), .A2(n674), .ZN(n583) );
  NAND2_X1 U673 ( .A1(n583), .A2(KEYINPUT47), .ZN(n587) );
  NOR2_X1 U674 ( .A1(KEYINPUT47), .A2(n585), .ZN(n586) );
  NAND2_X1 U675 ( .A1(n589), .A2(n588), .ZN(n590) );
  INV_X1 U676 ( .A(n676), .ZN(n593) );
  NAND2_X1 U677 ( .A1(n591), .A2(n704), .ZN(n592) );
  NOR2_X1 U678 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U679 ( .A1(n594), .A2(n609), .ZN(n602) );
  NOR2_X1 U680 ( .A1(n605), .A2(n602), .ZN(n595) );
  XNOR2_X1 U681 ( .A(n595), .B(KEYINPUT36), .ZN(n596) );
  AND2_X1 U682 ( .A1(n596), .A2(n616), .ZN(n683) );
  NAND2_X1 U683 ( .A1(n599), .A2(n598), .ZN(n601) );
  NOR2_X1 U684 ( .A1(n602), .A2(n616), .ZN(n604) );
  XOR2_X1 U685 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n603) );
  XNOR2_X1 U686 ( .A(n604), .B(n603), .ZN(n606) );
  NAND2_X1 U687 ( .A1(n606), .A2(n605), .ZN(n685) );
  NAND2_X1 U688 ( .A1(n607), .A2(n679), .ZN(n608) );
  XNOR2_X1 U689 ( .A(n608), .B(KEYINPUT116), .ZN(n758) );
  NOR2_X1 U690 ( .A1(n691), .A2(n558), .ZN(n610) );
  INV_X1 U691 ( .A(KEYINPUT32), .ZN(n611) );
  XNOR2_X1 U692 ( .A(n614), .B(KEYINPUT44), .ZN(n625) );
  XNOR2_X1 U693 ( .A(n615), .B(KEYINPUT88), .ZN(n618) );
  NOR2_X1 U694 ( .A1(n616), .A2(n564), .ZN(n617) );
  INV_X1 U695 ( .A(n694), .ZN(n619) );
  NOR2_X1 U696 ( .A1(n623), .A2(n620), .ZN(n667) );
  XNOR2_X1 U697 ( .A(n622), .B(KEYINPUT96), .ZN(n700) );
  INV_X1 U698 ( .A(n626), .ZN(n627) );
  NAND2_X1 U699 ( .A1(n627), .A2(KEYINPUT2), .ZN(n628) );
  XOR2_X1 U700 ( .A(KEYINPUT67), .B(n628), .Z(n629) );
  INV_X1 U701 ( .A(KEYINPUT65), .ZN(n630) );
  INV_X1 U702 ( .A(KEYINPUT81), .ZN(n631) );
  NAND2_X1 U703 ( .A1(n662), .A2(G475), .ZN(n635) );
  XNOR2_X1 U704 ( .A(KEYINPUT89), .B(KEYINPUT59), .ZN(n632) );
  XNOR2_X1 U705 ( .A(n635), .B(n634), .ZN(n638) );
  INV_X1 U706 ( .A(G952), .ZN(n636) );
  INV_X1 U707 ( .A(n731), .ZN(n658) );
  NAND2_X1 U708 ( .A1(n638), .A2(n658), .ZN(n640) );
  INV_X1 U709 ( .A(KEYINPUT60), .ZN(n639) );
  XNOR2_X1 U710 ( .A(n640), .B(n639), .ZN(G60) );
  NAND2_X1 U711 ( .A1(n662), .A2(G472), .ZN(n643) );
  XNOR2_X1 U712 ( .A(n643), .B(n642), .ZN(n644) );
  NAND2_X1 U713 ( .A1(n644), .A2(n658), .ZN(n645) );
  XNOR2_X1 U714 ( .A(n645), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U715 ( .A1(n662), .A2(G210), .ZN(n649) );
  XOR2_X1 U716 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n646) );
  XNOR2_X1 U717 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U718 ( .A(n649), .B(n648), .ZN(n650) );
  NAND2_X1 U719 ( .A1(n650), .A2(n658), .ZN(n652) );
  INV_X1 U720 ( .A(KEYINPUT56), .ZN(n651) );
  XNOR2_X1 U721 ( .A(n652), .B(n651), .ZN(G51) );
  NAND2_X1 U722 ( .A1(n662), .A2(G469), .ZN(n657) );
  XNOR2_X1 U723 ( .A(KEYINPUT122), .B(KEYINPUT57), .ZN(n653) );
  XNOR2_X1 U724 ( .A(n653), .B(KEYINPUT58), .ZN(n654) );
  XNOR2_X1 U725 ( .A(n657), .B(n656), .ZN(n659) );
  NAND2_X1 U726 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U727 ( .A(n660), .B(KEYINPUT123), .ZN(G54) );
  AND2_X1 U728 ( .A1(n662), .A2(G217), .ZN(n663) );
  XNOR2_X1 U729 ( .A(n661), .B(n663), .ZN(n664) );
  NOR2_X1 U730 ( .A1(n664), .A2(n731), .ZN(G66) );
  XOR2_X1 U731 ( .A(G104), .B(KEYINPUT117), .Z(n666) );
  NAND2_X1 U732 ( .A1(n667), .A2(n676), .ZN(n665) );
  XNOR2_X1 U733 ( .A(n666), .B(n665), .ZN(G6) );
  XOR2_X1 U734 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n669) );
  NAND2_X1 U735 ( .A1(n667), .A2(n679), .ZN(n668) );
  XNOR2_X1 U736 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U737 ( .A(G107), .B(n670), .ZN(G9) );
  XOR2_X1 U738 ( .A(G128), .B(KEYINPUT29), .Z(n672) );
  NAND2_X1 U739 ( .A1(n674), .A2(n679), .ZN(n671) );
  XNOR2_X1 U740 ( .A(n672), .B(n671), .ZN(G30) );
  XOR2_X1 U741 ( .A(G143), .B(n673), .Z(G45) );
  NAND2_X1 U742 ( .A1(n676), .A2(n674), .ZN(n675) );
  XNOR2_X1 U743 ( .A(n675), .B(G146), .ZN(G48) );
  NAND2_X1 U744 ( .A1(n676), .A2(n680), .ZN(n677) );
  XNOR2_X1 U745 ( .A(n677), .B(KEYINPUT118), .ZN(n678) );
  XNOR2_X1 U746 ( .A(G113), .B(n678), .ZN(G15) );
  NAND2_X1 U747 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U748 ( .A(n681), .B(G116), .ZN(G18) );
  XNOR2_X1 U749 ( .A(KEYINPUT37), .B(KEYINPUT119), .ZN(n682) );
  XOR2_X1 U750 ( .A(n683), .B(n682), .Z(n684) );
  XNOR2_X1 U751 ( .A(G125), .B(n684), .ZN(G27) );
  XNOR2_X1 U752 ( .A(G140), .B(n685), .ZN(G42) );
  INV_X1 U753 ( .A(n686), .ZN(n689) );
  NOR2_X1 U754 ( .A1(n687), .A2(KEYINPUT2), .ZN(n688) );
  NOR2_X1 U755 ( .A1(n689), .A2(n688), .ZN(n725) );
  NAND2_X1 U756 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U757 ( .A(KEYINPUT50), .B(n692), .Z(n693) );
  NOR2_X1 U758 ( .A1(n694), .A2(n693), .ZN(n698) );
  NOR2_X1 U759 ( .A1(n558), .A2(n695), .ZN(n696) );
  XNOR2_X1 U760 ( .A(n696), .B(KEYINPUT49), .ZN(n697) );
  NAND2_X1 U761 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U762 ( .A(KEYINPUT120), .B(n699), .ZN(n701) );
  NAND2_X1 U763 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U764 ( .A(KEYINPUT51), .B(n702), .ZN(n703) );
  NOR2_X1 U765 ( .A1(n703), .A2(n719), .ZN(n714) );
  NOR2_X1 U766 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U767 ( .A1(n707), .A2(n706), .ZN(n710) );
  NOR2_X1 U768 ( .A1(n710), .A2(n709), .ZN(n712) );
  INV_X1 U769 ( .A(n711), .ZN(n718) );
  NOR2_X1 U770 ( .A1(n712), .A2(n718), .ZN(n713) );
  NOR2_X1 U771 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U772 ( .A(n715), .B(KEYINPUT52), .ZN(n716) );
  NOR2_X1 U773 ( .A1(n717), .A2(n716), .ZN(n721) );
  NOR2_X1 U774 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U775 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U776 ( .A(KEYINPUT121), .B(n722), .Z(n723) );
  NAND2_X1 U777 ( .A1(n723), .A2(n736), .ZN(n724) );
  NOR2_X1 U778 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U779 ( .A(KEYINPUT53), .B(n726), .ZN(G75) );
  NAND2_X1 U780 ( .A1(n662), .A2(G478), .ZN(n729) );
  XOR2_X1 U781 ( .A(KEYINPUT124), .B(n727), .Z(n728) );
  XNOR2_X1 U782 ( .A(n729), .B(n728), .ZN(n730) );
  NOR2_X1 U783 ( .A1(n731), .A2(n730), .ZN(G63) );
  XNOR2_X1 U784 ( .A(n733), .B(n732), .ZN(n734) );
  NOR2_X1 U785 ( .A1(n735), .A2(n734), .ZN(n743) );
  XOR2_X1 U786 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n738) );
  NAND2_X1 U787 ( .A1(G224), .A2(G953), .ZN(n737) );
  XNOR2_X1 U788 ( .A(n738), .B(n737), .ZN(n739) );
  NAND2_X1 U789 ( .A1(n739), .A2(G898), .ZN(n740) );
  NAND2_X1 U790 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U791 ( .A(n743), .B(n742), .ZN(G69) );
  INV_X1 U792 ( .A(KEYINPUT126), .ZN(n744) );
  XNOR2_X1 U793 ( .A(n745), .B(n744), .ZN(n746) );
  XNOR2_X1 U794 ( .A(n747), .B(n746), .ZN(n751) );
  XOR2_X1 U795 ( .A(n748), .B(n751), .Z(n750) );
  NAND2_X1 U796 ( .A1(n750), .A2(n749), .ZN(n756) );
  XNOR2_X1 U797 ( .A(G227), .B(n751), .ZN(n752) );
  NAND2_X1 U798 ( .A1(n752), .A2(G900), .ZN(n753) );
  NAND2_X1 U799 ( .A1(G953), .A2(n753), .ZN(n754) );
  XOR2_X1 U800 ( .A(KEYINPUT127), .B(n754), .Z(n755) );
  NAND2_X1 U801 ( .A1(n756), .A2(n755), .ZN(G72) );
  XOR2_X1 U802 ( .A(G119), .B(n757), .Z(G21) );
  XNOR2_X1 U803 ( .A(G134), .B(n758), .ZN(G36) );
endmodule

