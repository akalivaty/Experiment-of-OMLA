//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 0 0 0 0 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1295, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1302, new_n1303,
    new_n1304, new_n1305, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1357, new_n1358, new_n1359;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n206), .A2(new_n207), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n212), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(KEYINPUT65), .B(G77), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G58), .A2(G232), .ZN(new_n229));
  NAND4_X1  g0029(.A1(new_n226), .A2(new_n227), .A3(new_n228), .A4(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n214), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n217), .B(new_n221), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT66), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n232), .A2(new_n234), .ZN(G361));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(G226), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XOR2_X1   g0049(.A(G107), .B(G116), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  NAND2_X1  g0052(.A1(G33), .A2(G97), .ZN(new_n253));
  AND2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  OAI211_X1 g0055(.A(G232), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT69), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT69), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G1698), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n258), .B(new_n260), .C1(new_n254), .C2(new_n255), .ZN(new_n261));
  INV_X1    g0061(.A(G226), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n253), .B(new_n256), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT76), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT69), .B(G1698), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n269), .A2(new_n270), .A3(G226), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT76), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n271), .A2(new_n272), .A3(new_n253), .A4(new_n256), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n264), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT13), .ZN(new_n276));
  INV_X1    g0076(.A(G41), .ZN(new_n277));
  INV_X1    g0077(.A(G45), .ZN(new_n278));
  AOI21_X1  g0078(.A(G1), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G41), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(G1), .A3(G13), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(new_n281), .A3(G274), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n283), .B1(G238), .B2(new_n286), .ZN(new_n287));
  AND3_X1   g0087(.A1(new_n275), .A2(new_n276), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n276), .B1(new_n275), .B2(new_n287), .ZN(new_n289));
  OAI21_X1  g0089(.A(G200), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n275), .A2(new_n287), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT13), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n275), .A2(new_n276), .A3(new_n287), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n292), .A2(G190), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n219), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(new_n211), .B2(G20), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G68), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n298), .B(KEYINPUT77), .ZN(new_n299));
  INV_X1    g0099(.A(new_n296), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT72), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(new_n212), .A3(new_n266), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT72), .B1(G20), .B2(G33), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G50), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n212), .A2(G33), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n307), .A2(G77), .B1(G20), .B2(new_n202), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n300), .B1(new_n305), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n299), .B1(KEYINPUT11), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(KEYINPUT11), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n202), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n314), .B(KEYINPUT12), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n310), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n290), .A2(new_n294), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G169), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n319), .B1(new_n292), .B2(new_n293), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT78), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT14), .ZN(new_n322));
  NOR3_X1   g0122(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(G169), .B1(new_n288), .B2(new_n289), .ZN(new_n324));
  AOI21_X1  g0124(.A(KEYINPUT78), .B1(new_n324), .B2(KEYINPUT14), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n322), .B(G169), .C1(new_n288), .C2(new_n289), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n292), .A2(G179), .A3(new_n293), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NOR3_X1   g0128(.A1(new_n323), .A2(new_n325), .A3(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n318), .B1(new_n329), .B2(new_n317), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n208), .A2(G20), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n304), .A2(G150), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT8), .B(G58), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT71), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT8), .ZN(new_n335));
  OR3_X1    g0135(.A1(new_n335), .A2(KEYINPUT71), .A3(G58), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n331), .B(new_n332), .C1(new_n337), .C2(new_n306), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n296), .ZN(new_n339));
  INV_X1    g0139(.A(new_n297), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n340), .A2(new_n207), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n312), .A2(G50), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n269), .A2(new_n270), .A3(G222), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n269), .A2(G1698), .ZN(new_n346));
  XOR2_X1   g0146(.A(KEYINPUT70), .B(G223), .Z(new_n347));
  OAI221_X1 g0147(.A(new_n345), .B1(new_n223), .B2(new_n269), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n274), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n283), .B1(G226), .B2(new_n286), .ZN(new_n350));
  AOI21_X1  g0150(.A(G169), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(KEYINPUT73), .B1(new_n344), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT73), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n339), .A2(new_n343), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n349), .A2(new_n350), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n353), .B(new_n354), .C1(new_n355), .C2(G169), .ZN(new_n356));
  XNOR2_X1  g0156(.A(KEYINPUT74), .B(G179), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n352), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT75), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n352), .A2(new_n356), .A3(KEYINPUT75), .A4(new_n358), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G200), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(new_n349), .B2(new_n350), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n365), .B1(new_n355), .B2(G190), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT9), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n344), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n354), .A2(KEYINPUT9), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n366), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT10), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT10), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n366), .B(new_n372), .C1(new_n368), .C2(new_n369), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n254), .A2(new_n255), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G107), .ZN(new_n376));
  INV_X1    g0176(.A(G232), .ZN(new_n377));
  INV_X1    g0177(.A(G238), .ZN(new_n378));
  OAI221_X1 g0178(.A(new_n376), .B1(new_n261), .B2(new_n377), .C1(new_n346), .C2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n274), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n283), .B1(G244), .B2(new_n286), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  XNOR2_X1  g0183(.A(KEYINPUT15), .B(G87), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n385), .A2(new_n307), .B1(new_n222), .B2(G20), .ZN(new_n386));
  INV_X1    g0186(.A(new_n333), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n304), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n300), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G77), .ZN(new_n390));
  OAI22_X1  g0190(.A1(new_n340), .A2(new_n390), .B1(new_n222), .B2(new_n312), .ZN(new_n391));
  OAI22_X1  g0191(.A1(new_n383), .A2(G169), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n357), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n382), .A2(new_n393), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n382), .A2(G200), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n389), .A2(new_n391), .ZN(new_n397));
  INV_X1    g0197(.A(G190), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n396), .B(new_n397), .C1(new_n398), .C2(new_n382), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n363), .A2(new_n374), .A3(new_n400), .ZN(new_n401));
  OAI211_X1 g0201(.A(G226), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G33), .A2(G87), .ZN(new_n403));
  INV_X1    g0203(.A(G223), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n402), .B(new_n403), .C1(new_n261), .C2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n274), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n282), .B1(new_n377), .B2(new_n285), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(new_n398), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n407), .B1(new_n274), .B2(new_n405), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n409), .B1(G200), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT16), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n267), .A2(new_n212), .A3(new_n268), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT7), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n375), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n202), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G58), .A2(G68), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n203), .A2(new_n205), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G20), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n304), .A2(G159), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n412), .B1(new_n417), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT7), .B1(new_n375), .B2(new_n212), .ZN(new_n424));
  NOR4_X1   g0224(.A1(new_n254), .A2(new_n255), .A3(new_n414), .A4(G20), .ZN(new_n425));
  OAI21_X1  g0225(.A(G68), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n419), .A2(G20), .B1(new_n304), .B2(G159), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n426), .A2(KEYINPUT16), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n423), .A2(new_n428), .A3(new_n296), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n337), .A2(new_n312), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n297), .B2(new_n337), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n411), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT17), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n431), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n426), .A2(new_n427), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n300), .B1(new_n436), .B2(new_n412), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n435), .B1(new_n437), .B2(new_n428), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n438), .A2(KEYINPUT17), .A3(new_n411), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n429), .A2(new_n431), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n410), .A2(new_n393), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n319), .B2(new_n410), .ZN(new_n442));
  AOI21_X1  g0242(.A(KEYINPUT18), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT79), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n440), .A2(KEYINPUT18), .A3(new_n442), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n440), .A2(new_n442), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT18), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n447), .A2(new_n444), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n434), .B(new_n439), .C1(new_n446), .C2(new_n450), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n330), .A2(new_n401), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT84), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT19), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n212), .B1(new_n253), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(G97), .A2(G107), .ZN(new_n457));
  INV_X1    g0257(.A(G87), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n212), .B(G68), .C1(new_n254), .C2(new_n255), .ZN(new_n461));
  INV_X1    g0261(.A(G97), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n455), .B1(new_n306), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n460), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT83), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n300), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT83), .A4(new_n463), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n385), .A2(new_n312), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n211), .A2(G33), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n300), .A2(new_n312), .A3(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(new_n458), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n468), .A2(new_n470), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n211), .A2(G45), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n281), .A2(G250), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n281), .A2(G274), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n477), .B1(new_n478), .B2(new_n476), .ZN(new_n479));
  OAI211_X1 g0279(.A(G244), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G116), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n480), .B(new_n481), .C1(new_n261), .C2(new_n378), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n479), .B1(new_n482), .B2(new_n274), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(new_n364), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n454), .B1(new_n475), .B2(new_n484), .ZN(new_n485));
  AOI211_X1 g0285(.A(new_n469), .B(new_n473), .C1(new_n466), .C2(new_n467), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n482), .A2(new_n274), .ZN(new_n487));
  INV_X1    g0287(.A(new_n479), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G200), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n486), .A2(KEYINPUT84), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n483), .A2(G190), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n485), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n468), .B(new_n470), .C1(new_n384), .C2(new_n472), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n489), .A2(new_n319), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n483), .A2(new_n357), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT82), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n483), .A2(KEYINPUT82), .A3(new_n357), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n494), .A2(new_n495), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n493), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT4), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(new_n261), .B2(new_n224), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n269), .A2(new_n270), .A3(KEYINPUT4), .A4(G244), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G283), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(G250), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT81), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n269), .A2(KEYINPUT81), .A3(G250), .A4(G1698), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n274), .B1(new_n506), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT5), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n277), .ZN(new_n514));
  NAND2_X1  g0314(.A1(KEYINPUT5), .A2(G41), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n278), .A2(G1), .ZN(new_n517));
  INV_X1    g0317(.A(new_n219), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n516), .A2(new_n517), .B1(new_n518), .B2(new_n280), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G257), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n476), .B1(new_n514), .B2(new_n515), .ZN(new_n521));
  INV_X1    g0321(.A(G274), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n522), .B1(new_n518), .B2(new_n280), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n512), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G200), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n509), .A2(new_n510), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n529), .A2(new_n504), .A3(new_n505), .A4(new_n503), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n525), .B1(new_n530), .B2(new_n274), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(G190), .ZN(new_n532));
  OAI21_X1  g0332(.A(G107), .B1(new_n424), .B2(new_n425), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT6), .ZN(new_n534));
  AND2_X1   g0334(.A1(G97), .A2(G107), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n534), .B1(new_n535), .B2(new_n457), .ZN(new_n536));
  INV_X1    g0336(.A(G107), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n537), .A2(KEYINPUT6), .A3(G97), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n539), .A2(G20), .B1(G77), .B2(new_n304), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n300), .B1(new_n533), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n312), .A2(G97), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n472), .B2(new_n462), .ZN(new_n544));
  OAI21_X1  g0344(.A(KEYINPUT80), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n533), .A2(new_n540), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n296), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT80), .ZN(new_n548));
  INV_X1    g0348(.A(new_n544), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n528), .A2(new_n532), .A3(new_n545), .A4(new_n550), .ZN(new_n551));
  AOI211_X1 g0351(.A(new_n357), .B(new_n525), .C1(new_n530), .C2(new_n274), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n319), .B1(new_n512), .B2(new_n526), .ZN(new_n553));
  OAI22_X1  g0353(.A1(new_n552), .A2(new_n553), .B1(new_n541), .B2(new_n544), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(G257), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n556));
  NAND2_X1  g0356(.A1(G33), .A2(G294), .ZN(new_n557));
  OAI21_X1  g0357(.A(G250), .B1(new_n254), .B2(new_n255), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n258), .A2(new_n260), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n556), .B(new_n557), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n560), .A2(new_n274), .B1(G264), .B2(new_n519), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n319), .B1(new_n561), .B2(new_n524), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n274), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n519), .A2(G264), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n563), .A2(new_n524), .A3(new_n564), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n562), .A2(KEYINPUT87), .B1(new_n565), .B2(G179), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n563), .A2(new_n524), .A3(new_n564), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(G169), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT87), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n212), .B(G87), .C1(new_n254), .C2(new_n255), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT22), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT22), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n269), .A2(new_n573), .A3(new_n212), .A4(G87), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT24), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n481), .A2(G20), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT23), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n212), .B2(G107), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n537), .A2(KEYINPUT23), .A3(G20), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n577), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n575), .A2(new_n576), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n576), .B1(new_n575), .B2(new_n581), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n296), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n472), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT86), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(KEYINPUT25), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n537), .B1(new_n586), .B2(KEYINPUT25), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n587), .B1(new_n588), .B2(new_n312), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n313), .A2(new_n586), .A3(KEYINPUT25), .A4(new_n537), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n585), .A2(G107), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n566), .A2(new_n570), .B1(new_n584), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n561), .A2(G190), .A3(new_n524), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n567), .A2(G200), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n584), .A2(new_n591), .A3(new_n593), .A4(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(KEYINPUT88), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n267), .A2(G303), .A3(new_n268), .ZN(new_n598));
  OAI211_X1 g0398(.A(G264), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n599));
  INV_X1    g0399(.A(G257), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n598), .B(new_n599), .C1(new_n261), .C2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n274), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n519), .A2(G270), .B1(new_n523), .B2(new_n521), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n604), .A2(KEYINPUT21), .A3(G169), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n602), .A2(new_n603), .A3(G179), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(G116), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n313), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n300), .A2(G116), .A3(new_n312), .A4(new_n471), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n295), .A2(new_n219), .B1(G20), .B2(new_n608), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n505), .B(new_n212), .C1(G33), .C2(new_n462), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n611), .A2(KEYINPUT20), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(KEYINPUT20), .B1(new_n611), .B2(new_n612), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n609), .B(new_n610), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n607), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n615), .B1(new_n604), .B2(G200), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(new_n398), .B2(new_n604), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n604), .A2(G169), .A3(new_n615), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT21), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(KEYINPUT85), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT85), .B1(new_n619), .B2(new_n620), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n616), .B(new_n618), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n584), .A2(new_n591), .ZN(new_n626));
  INV_X1    g0426(.A(G179), .ZN(new_n627));
  OAI22_X1  g0427(.A1(new_n568), .A2(new_n569), .B1(new_n627), .B2(new_n567), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n562), .A2(KEYINPUT87), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n626), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT88), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(new_n631), .A3(new_n595), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n597), .A2(new_n625), .A3(new_n632), .ZN(new_n633));
  NOR4_X1   g0433(.A1(new_n453), .A2(new_n501), .A3(new_n555), .A4(new_n633), .ZN(G372));
  OAI21_X1  g0434(.A(new_n321), .B1(new_n320), .B2(new_n322), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n324), .A2(KEYINPUT78), .A3(KEYINPUT14), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n635), .A2(new_n636), .A3(new_n326), .A4(new_n327), .ZN(new_n637));
  INV_X1    g0437(.A(new_n317), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n392), .A2(new_n394), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n637), .A2(new_n638), .B1(new_n318), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n439), .A2(new_n434), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n440), .A2(KEYINPUT18), .A3(new_n442), .ZN(new_n642));
  OAI22_X1  g0442(.A1(new_n640), .A2(new_n641), .B1(new_n443), .B2(new_n642), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n643), .A2(new_n374), .B1(new_n361), .B2(new_n362), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT89), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n489), .A2(new_n647), .A3(G200), .ZN(new_n648));
  OAI21_X1  g0448(.A(KEYINPUT89), .B1(new_n483), .B2(new_n364), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n486), .A2(new_n648), .A3(new_n492), .A4(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n548), .B1(new_n547), .B2(new_n549), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n541), .A2(KEYINPUT80), .A3(new_n544), .ZN(new_n653));
  OAI22_X1  g0453(.A1(new_n552), .A2(new_n553), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n645), .B1(new_n651), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(KEYINPUT90), .ZN(new_n656));
  INV_X1    g0456(.A(new_n554), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n657), .A2(KEYINPUT26), .A3(new_n500), .A4(new_n493), .ZN(new_n658));
  INV_X1    g0458(.A(new_n553), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n531), .A2(new_n393), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n550), .A2(new_n545), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n661), .A2(new_n662), .A3(new_n646), .A4(new_n650), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT90), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(new_n664), .A3(new_n645), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n656), .A2(new_n658), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n646), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n646), .A2(new_n595), .A3(new_n650), .ZN(new_n668));
  INV_X1    g0468(.A(new_n615), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n669), .B1(new_n605), .B2(new_n606), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n619), .A2(new_n620), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT85), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n670), .B1(new_n673), .B2(new_n621), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n668), .B1(new_n674), .B2(new_n630), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n551), .A2(new_n554), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n667), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n666), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n644), .B1(new_n453), .B2(new_n679), .ZN(G369));
  NAND3_X1  g0480(.A1(new_n211), .A2(new_n212), .A3(G13), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G213), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G343), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n669), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n624), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n616), .B1(new_n622), .B2(new_n623), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n688), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G330), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT91), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n592), .A2(KEYINPUT88), .A3(new_n596), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n631), .B1(new_n630), .B2(new_n595), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n626), .A2(new_n686), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n592), .A2(new_n686), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n694), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n690), .A2(new_n687), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n697), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n592), .A2(new_n687), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n702), .A2(new_n708), .ZN(G399));
  INV_X1    g0509(.A(new_n215), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(G41), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n459), .A2(G116), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(G1), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n218), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n714), .B1(new_n715), .B2(new_n712), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT92), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT28), .ZN(new_n718));
  AOI211_X1 g0518(.A(KEYINPUT29), .B(new_n686), .C1(new_n666), .C2(new_n677), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT29), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT95), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n555), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n674), .A2(new_n630), .ZN(new_n723));
  INV_X1    g0523(.A(new_n668), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n551), .A2(new_n554), .A3(KEYINPUT95), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n722), .A2(new_n723), .A3(new_n724), .A4(new_n725), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n493), .A2(new_n500), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n727), .A2(new_n645), .A3(new_n657), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n667), .B1(new_n663), .B2(KEYINPUT26), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n726), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n720), .B1(new_n730), .B2(new_n687), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n719), .A2(new_n731), .ZN(new_n732));
  AND4_X1   g0532(.A1(new_n487), .A2(new_n563), .A3(new_n488), .A4(new_n564), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n602), .A2(new_n603), .A3(G179), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n531), .A2(new_n733), .A3(KEYINPUT30), .A4(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT93), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT30), .ZN(new_n738));
  INV_X1    g0538(.A(new_n515), .ZN(new_n739));
  NOR2_X1   g0539(.A1(KEYINPUT5), .A2(G41), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n517), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(G270), .A3(new_n281), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(new_n524), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n743), .B1(new_n274), .B2(new_n601), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n744), .A2(G179), .A3(new_n483), .A4(new_n561), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n738), .B1(new_n745), .B2(new_n527), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n744), .A2(new_n393), .A3(new_n483), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n747), .A2(new_n527), .A3(new_n567), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n483), .A2(new_n561), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n606), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n750), .A2(KEYINPUT93), .A3(KEYINPUT30), .A4(new_n531), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n737), .A2(new_n746), .A3(new_n748), .A4(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n752), .A2(KEYINPUT31), .A3(new_n686), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT94), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n752), .A2(KEYINPUT94), .A3(KEYINPUT31), .A4(new_n686), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n752), .A2(new_n686), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT31), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n755), .A2(new_n756), .A3(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n727), .A2(new_n676), .A3(new_n687), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n633), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(G330), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n732), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n718), .B1(new_n765), .B2(G1), .ZN(G364));
  INV_X1    g0566(.A(KEYINPUT91), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n693), .B(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G13), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n211), .B1(new_n770), .B2(G45), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n768), .B1(G330), .B2(new_n692), .C1(new_n711), .C2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n711), .A2(new_n772), .ZN(new_n774));
  XOR2_X1   g0574(.A(new_n774), .B(KEYINPUT96), .Z(new_n775));
  NOR2_X1   g0575(.A1(new_n710), .A2(new_n375), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G355), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(G116), .B2(new_n215), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n710), .A2(new_n269), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n779), .B(KEYINPUT97), .Z(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(new_n278), .B2(new_n218), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n248), .A2(G45), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n778), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G13), .A2(G33), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT98), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G20), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n219), .B1(G20), .B2(new_n319), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n775), .B1(new_n784), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n357), .A2(new_n212), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G200), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n398), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(G190), .ZN(new_n795));
  AOI22_X1  g0595(.A1(G50), .A2(new_n794), .B1(new_n795), .B2(G68), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n212), .A2(G179), .ZN(new_n797));
  NOR2_X1   g0597(.A1(G190), .A2(G200), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G159), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT32), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n398), .A2(G200), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n212), .B1(new_n803), .B2(new_n627), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n462), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n797), .A2(new_n398), .A3(G200), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(new_n537), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n797), .A2(G190), .A3(G200), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n458), .ZN(new_n809));
  NOR4_X1   g0609(.A1(new_n805), .A2(new_n807), .A3(new_n809), .A4(new_n375), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n796), .A2(new_n802), .A3(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT99), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n792), .A2(new_n812), .ZN(new_n813));
  NOR3_X1   g0613(.A1(new_n357), .A2(KEYINPUT99), .A3(new_n212), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n803), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n798), .B1(new_n813), .B2(new_n814), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n201), .A2(new_n815), .B1(new_n816), .B2(new_n223), .ZN(new_n817));
  INV_X1    g0617(.A(G283), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n806), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n799), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n269), .B(new_n819), .C1(G329), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n794), .A2(G326), .ZN(new_n822));
  XNOR2_X1  g0622(.A(KEYINPUT33), .B(G317), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n795), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n804), .ZN(new_n825));
  INV_X1    g0625(.A(new_n808), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n825), .A2(G294), .B1(new_n826), .B2(G303), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n821), .A2(new_n822), .A3(new_n824), .A4(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(G311), .ZN(new_n829));
  INV_X1    g0629(.A(G322), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n829), .A2(new_n816), .B1(new_n815), .B2(new_n830), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n811), .A2(new_n817), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n791), .B1(new_n788), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n787), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n833), .B1(new_n692), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n773), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(G396));
  OAI21_X1  g0637(.A(new_n399), .B1(new_n397), .B2(new_n687), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n395), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n639), .A2(new_n687), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n679), .B2(new_n686), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n400), .A2(new_n687), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(new_n666), .B2(new_n677), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n763), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n711), .B2(new_n772), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n846), .A2(new_n763), .ZN(new_n849));
  INV_X1    g0649(.A(new_n788), .ZN(new_n850));
  AOI22_X1  g0650(.A1(G137), .A2(new_n794), .B1(new_n795), .B2(G150), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n800), .B2(new_n816), .ZN(new_n852));
  INV_X1    g0652(.A(new_n815), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n852), .B1(G143), .B2(new_n853), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT100), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n855), .A2(KEYINPUT34), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n207), .A2(new_n808), .B1(new_n806), .B2(new_n202), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT101), .ZN(new_n858));
  INV_X1    g0658(.A(G132), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n269), .B1(new_n799), .B2(new_n859), .C1(new_n804), .C2(new_n201), .ZN(new_n860));
  NOR3_X1   g0660(.A1(new_n856), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(KEYINPUT34), .B2(new_n855), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n269), .B(new_n805), .C1(G311), .C2(new_n820), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n863), .B1(new_n458), .B2(new_n806), .C1(new_n537), .C2(new_n808), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(G283), .B2(new_n795), .ZN(new_n865));
  INV_X1    g0665(.A(new_n816), .ZN(new_n866));
  AOI22_X1  g0666(.A1(G116), .A2(new_n866), .B1(new_n853), .B2(G294), .ZN(new_n867));
  INV_X1    g0667(.A(G303), .ZN(new_n868));
  INV_X1    g0668(.A(new_n794), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n865), .B(new_n867), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n850), .B1(new_n862), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n785), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n850), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n841), .ZN(new_n874));
  OAI221_X1 g0674(.A(new_n775), .B1(G77), .B2(new_n873), .C1(new_n874), .C2(new_n786), .ZN(new_n875));
  OAI22_X1  g0675(.A1(new_n848), .A2(new_n849), .B1(new_n871), .B2(new_n875), .ZN(G384));
  OR2_X1    g0676(.A1(new_n539), .A2(KEYINPUT35), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n539), .A2(KEYINPUT35), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n877), .A2(G116), .A3(new_n220), .A4(new_n878), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n879), .B(KEYINPUT36), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n218), .A2(new_n222), .A3(new_n418), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(G50), .B2(new_n202), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n882), .A2(G1), .A3(new_n769), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n883), .B(KEYINPUT102), .Z(new_n884));
  INV_X1    g0684(.A(G330), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT40), .ZN(new_n886));
  INV_X1    g0686(.A(new_n432), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT104), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n440), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n429), .A2(new_n431), .A3(KEYINPUT104), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n887), .B1(new_n891), .B2(new_n442), .ZN(new_n892));
  INV_X1    g0692(.A(new_n684), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n429), .A2(new_n431), .A3(KEYINPUT104), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT104), .B1(new_n429), .B2(new_n431), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT105), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT105), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n891), .A2(new_n898), .A3(new_n893), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n892), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(KEYINPUT37), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n440), .A2(new_n893), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT37), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n447), .A2(new_n902), .A3(new_n903), .A4(new_n432), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n897), .A2(new_n899), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n451), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT38), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n909), .B1(new_n451), .B2(new_n906), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n908), .A2(new_n909), .B1(new_n905), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n638), .A2(new_n686), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n318), .B(new_n912), .C1(new_n329), .C2(new_n317), .ZN(new_n913));
  INV_X1    g0713(.A(new_n318), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n638), .B(new_n686), .C1(new_n637), .C2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n841), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n753), .B(new_n759), .C1(new_n633), .C2(new_n761), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n886), .B1(new_n911), .B2(new_n918), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n434), .B(new_n439), .C1(new_n642), .C2(new_n443), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n438), .A2(new_n684), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n410), .A2(new_n319), .ZN(new_n923));
  AND3_X1   g0723(.A1(new_n406), .A2(new_n408), .A3(new_n393), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n432), .B1(new_n438), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT37), .B1(new_n926), .B2(new_n921), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n904), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n922), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT106), .B1(new_n929), .B2(new_n909), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT106), .ZN(new_n931));
  AOI211_X1 g0731(.A(new_n931), .B(KEYINPUT38), .C1(new_n922), .C2(new_n928), .ZN(new_n932));
  INV_X1    g0732(.A(new_n904), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(new_n900), .B2(KEYINPUT37), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n897), .A2(new_n899), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n447), .A2(new_n448), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n642), .B2(KEYINPUT79), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n641), .B1(new_n937), .B2(new_n449), .ZN(new_n938));
  OAI21_X1  g0738(.A(KEYINPUT38), .B1(new_n935), .B2(new_n938), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n930), .A2(new_n932), .B1(new_n934), .B2(new_n939), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n940), .A2(KEYINPUT40), .A3(new_n917), .A4(new_n916), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n919), .A2(new_n941), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n452), .A2(new_n917), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n885), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n942), .B2(new_n943), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n913), .A2(new_n915), .ZN(new_n946));
  INV_X1    g0746(.A(new_n840), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n946), .B1(new_n844), .B2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT103), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n946), .B(KEYINPUT103), .C1(new_n844), .C2(new_n947), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n935), .A2(new_n938), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n909), .B1(new_n952), .B2(new_n934), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n905), .A2(new_n910), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n950), .A2(new_n951), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n953), .A2(new_n954), .A3(KEYINPUT39), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n637), .A2(new_n638), .A3(new_n687), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n921), .A2(new_n920), .B1(new_n927), .B2(new_n904), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n931), .B1(new_n960), .B2(KEYINPUT38), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n929), .A2(KEYINPUT106), .A3(new_n909), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n961), .A2(new_n962), .B1(new_n905), .B2(new_n910), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n957), .B(new_n959), .C1(KEYINPUT39), .C2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n936), .A2(new_n445), .A3(new_n684), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n956), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n452), .B1(new_n719), .B2(new_n731), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n644), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n966), .B(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n945), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n211), .B2(new_n770), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n945), .A2(new_n969), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n880), .B(new_n884), .C1(new_n971), .C2(new_n972), .ZN(G367));
  NOR2_X1   g0773(.A1(new_n654), .A2(new_n687), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n722), .A2(new_n725), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n662), .A2(new_n686), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n707), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT44), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n978), .B(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n977), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n708), .A2(new_n981), .A3(KEYINPUT45), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT45), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n707), .B2(new_n977), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n980), .A2(new_n702), .A3(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n702), .B1(new_n980), .B2(new_n985), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n705), .B1(new_n701), .B2(new_n704), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n768), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n694), .A2(new_n990), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n765), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n764), .B1(new_n989), .B2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n711), .B(KEYINPUT41), .Z(new_n998));
  OAI21_X1  g0798(.A(new_n771), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n977), .A2(new_n705), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT42), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n554), .B1(new_n977), .B2(new_n630), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n687), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n475), .A2(new_n686), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n651), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n667), .B2(new_n1005), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT107), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT43), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1004), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1001), .A2(new_n1009), .A3(new_n1008), .A4(new_n1003), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n702), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n981), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1014), .B(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1008), .A2(new_n787), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n780), .A2(new_n243), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1020), .B(new_n789), .C1(new_n215), .C2(new_n384), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n775), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT108), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G294), .A2(new_n795), .B1(new_n794), .B2(G311), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n806), .A2(new_n462), .ZN(new_n1025));
  INV_X1    g0825(.A(G317), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n375), .B1(new_n799), .B2(new_n1026), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1025), .B(new_n1027), .C1(G107), .C2(new_n825), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n826), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT46), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n808), .B2(new_n608), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1024), .A2(new_n1028), .A3(new_n1029), .A4(new_n1031), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n818), .A2(new_n816), .B1(new_n815), .B2(new_n868), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n795), .A2(G159), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n794), .A2(G143), .ZN(new_n1035));
  INV_X1    g0835(.A(G137), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n269), .B1(new_n799), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(G58), .B2(new_n826), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n804), .A2(new_n202), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n806), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1039), .B1(new_n222), .B2(new_n1040), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1034), .A2(new_n1035), .A3(new_n1038), .A4(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(G150), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n207), .A2(new_n816), .B1(new_n815), .B2(new_n1043), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n1032), .A2(new_n1033), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT47), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n850), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n1046), .B2(new_n1045), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n1023), .A2(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n999), .A2(new_n1018), .B1(new_n1019), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(G387));
  NOR2_X1   g0851(.A1(new_n701), .A2(new_n834), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n713), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n776), .A2(new_n1053), .B1(new_n537), .B2(new_n710), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n387), .A2(new_n207), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT50), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n713), .B(new_n278), .C1(new_n202), .C2(new_n390), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n780), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n240), .A2(new_n278), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1054), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n789), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n775), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n337), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n866), .A2(G68), .B1(new_n1063), .B2(new_n795), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT109), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n375), .B(new_n1025), .C1(G150), .C2(new_n820), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n825), .A2(new_n385), .B1(new_n826), .B2(new_n222), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1066), .B(new_n1067), .C1(new_n800), .C2(new_n869), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(G50), .B2(new_n853), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1065), .A2(new_n1069), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G311), .A2(new_n795), .B1(new_n794), .B2(G322), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1071), .B1(new_n868), .B2(new_n816), .C1(new_n1026), .C2(new_n815), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT48), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n825), .A2(G283), .B1(new_n826), .B2(G294), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1078), .A2(KEYINPUT110), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(KEYINPUT110), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1079), .A2(KEYINPUT49), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1040), .A2(G116), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n269), .B1(new_n820), .B2(G326), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(KEYINPUT49), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1070), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1052), .B(new_n1062), .C1(new_n1086), .C2(new_n788), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n772), .B2(new_n994), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n995), .A2(new_n711), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n994), .A2(new_n765), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1088), .B1(new_n1089), .B2(new_n1090), .ZN(G393));
  NAND2_X1  g0891(.A1(new_n988), .A2(KEYINPUT111), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n988), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n986), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1092), .B1(new_n1094), .B2(KEYINPUT111), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n977), .A2(new_n787), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n775), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n789), .B1(new_n462), .B2(new_n215), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n780), .B2(new_n251), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n869), .A2(new_n1026), .B1(new_n815), .B2(new_n829), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT52), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n269), .B(new_n807), .C1(G322), .C2(new_n820), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n825), .A2(G116), .B1(new_n826), .B2(G283), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n795), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1102), .B(new_n1103), .C1(new_n868), .C2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(G294), .B2(new_n866), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1101), .A2(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n853), .A2(G159), .B1(G150), .B2(new_n794), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT112), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(KEYINPUT51), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n806), .A2(new_n458), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n375), .B(new_n1111), .C1(G143), .C2(new_n820), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n825), .A2(G77), .B1(new_n826), .B2(G68), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1112), .B(new_n1113), .C1(new_n207), .C2(new_n1104), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n387), .B2(new_n866), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1110), .A2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1109), .A2(KEYINPUT51), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1107), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n1097), .B(new_n1099), .C1(new_n1118), .C2(new_n788), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1095), .A2(new_n772), .B1(new_n1096), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n712), .B1(new_n989), .B2(new_n996), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n1095), .B2(new_n996), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1122), .ZN(G390));
  NAND4_X1  g0923(.A1(new_n946), .A2(G330), .A3(new_n917), .A4(new_n874), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT39), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n940), .A2(new_n1126), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1127), .A2(new_n957), .B1(new_n948), .B2(new_n958), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n730), .A2(new_n687), .A3(new_n839), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n1129), .A2(new_n840), .B1(new_n913), .B2(new_n915), .ZN(new_n1130));
  NOR3_X1   g0930(.A1(new_n1130), .A2(new_n959), .A3(new_n963), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1125), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n948), .A2(new_n958), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n957), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n961), .A2(new_n962), .ZN(new_n1135));
  AOI21_X1  g0935(.A(KEYINPUT39), .B1(new_n1135), .B2(new_n954), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1133), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1129), .A2(new_n840), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n913), .A2(new_n915), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n958), .B(new_n940), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n916), .B(G330), .C1(new_n762), .C2(new_n760), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1137), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1132), .A2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g0944(.A(G330), .B(new_n874), .C1(new_n760), .C2(new_n762), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n1140), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n1124), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n845), .A2(new_n840), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n917), .A2(G330), .A3(new_n874), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1140), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1142), .A2(new_n1151), .A3(new_n1139), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n452), .A2(G330), .A3(new_n917), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n967), .A2(new_n644), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1144), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1155), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1132), .A2(new_n1143), .A3(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1158), .A2(new_n711), .A3(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1132), .A2(new_n772), .A3(new_n1143), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n775), .B1(new_n1063), .B2(new_n873), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n269), .B(new_n809), .C1(G294), .C2(new_n820), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n825), .A2(G77), .B1(new_n1040), .B2(G68), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n1166), .B1(new_n537), .B2(new_n1104), .C1(new_n818), .C2(new_n869), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n462), .A2(new_n816), .B1(new_n815), .B2(new_n608), .ZN(new_n1168));
  INV_X1    g0968(.A(G128), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n1169), .A2(new_n869), .B1(new_n1104), .B2(new_n1036), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n808), .A2(new_n1043), .ZN(new_n1171));
  XOR2_X1   g0971(.A(new_n1171), .B(KEYINPUT53), .Z(new_n1172));
  AOI21_X1  g0972(.A(new_n375), .B1(new_n820), .B2(G125), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1173), .B1(new_n207), .B2(new_n806), .C1(new_n800), .C2(new_n804), .ZN(new_n1174));
  OR3_X1    g0974(.A1(new_n1170), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(KEYINPUT54), .B(G143), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n859), .A2(new_n815), .B1(new_n816), .B2(new_n1176), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n1167), .A2(new_n1168), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1163), .B1(new_n1178), .B2(new_n788), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1127), .A2(new_n957), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1179), .B1(new_n1181), .B2(new_n786), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1161), .A2(new_n1162), .A3(new_n1182), .ZN(G378));
  AOI21_X1  g0983(.A(new_n886), .B1(new_n1135), .B2(new_n954), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n946), .A2(new_n874), .A3(new_n917), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n885), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n344), .A2(new_n684), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n374), .B2(new_n359), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n374), .A2(new_n359), .A3(new_n1188), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1192), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  AND3_X1   g0996(.A1(new_n1186), .A2(new_n919), .A3(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1196), .B1(new_n1186), .B2(new_n919), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n966), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n956), .A2(new_n965), .A3(new_n964), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n941), .A2(G330), .ZN(new_n1201));
  AOI21_X1  g1001(.A(KEYINPUT40), .B1(new_n1185), .B2(new_n955), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1195), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1186), .A2(new_n919), .A3(new_n1196), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1200), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1199), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1160), .A2(new_n1156), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1206), .A2(new_n1207), .A3(KEYINPUT57), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n711), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT57), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT116), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1206), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1199), .A2(new_n1205), .A3(KEYINPUT116), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1212), .A2(new_n1207), .A3(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1209), .B1(new_n1210), .B2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1212), .A2(new_n772), .A3(new_n1213), .ZN(new_n1216));
  OR2_X1    g1016(.A1(new_n1196), .A2(new_n786), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n774), .B1(G50), .B2(new_n873), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n794), .A2(G125), .B1(G150), .B2(new_n825), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(new_n859), .B2(new_n1104), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n808), .A2(new_n1176), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT114), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n815), .B2(new_n1169), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT115), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1220), .B(new_n1224), .C1(G137), .C2(new_n866), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1225), .B(KEYINPUT59), .ZN(new_n1226));
  AOI211_X1 g1026(.A(G33), .B(G41), .C1(new_n820), .C2(G124), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1226), .B(new_n1227), .C1(new_n800), .C2(new_n806), .ZN(new_n1228));
  XOR2_X1   g1028(.A(KEYINPUT113), .B(KEYINPUT58), .Z(new_n1229));
  NAND2_X1  g1029(.A1(new_n375), .A2(new_n277), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n1230), .B(new_n1039), .C1(G283), .C2(new_n820), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n806), .A2(new_n201), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n222), .B2(new_n826), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1234), .B1(new_n462), .B2(new_n1104), .C1(new_n608), .C2(new_n869), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n537), .A2(new_n815), .B1(new_n816), .B2(new_n384), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1229), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1230), .B(new_n207), .C1(G33), .C2(G41), .ZN(new_n1238));
  OR3_X1    g1038(.A1(new_n1235), .A2(new_n1229), .A3(new_n1236), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1228), .A2(new_n1237), .A3(new_n1238), .A4(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1218), .B1(new_n1240), .B2(new_n788), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1217), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1216), .A2(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(KEYINPUT117), .B1(new_n1215), .B2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT117), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1242), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1199), .A2(new_n1205), .A3(KEYINPUT116), .ZN(new_n1247));
  AOI21_X1  g1047(.A(KEYINPUT116), .B1(new_n1199), .B2(new_n1205), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1246), .B1(new_n1249), .B2(new_n772), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT57), .B1(new_n1249), .B2(new_n1207), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1245), .B(new_n1250), .C1(new_n1251), .C2(new_n1209), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1244), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(G375));
  NAND2_X1  g1054(.A1(new_n1153), .A2(new_n772), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n775), .B1(G68), .B2(new_n873), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n825), .A2(new_n385), .B1(new_n820), .B2(G303), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1257), .B1(new_n462), .B2(new_n808), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n269), .B1(new_n1040), .B2(G77), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1258), .B1(KEYINPUT118), .B2(new_n1259), .ZN(new_n1260));
  OAI221_X1 g1060(.A(new_n1260), .B1(new_n537), .B2(new_n816), .C1(new_n818), .C2(new_n815), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(G116), .A2(new_n795), .B1(new_n794), .B2(G294), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(KEYINPUT118), .B2(new_n1259), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n269), .B1(new_n799), .B2(new_n1169), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n804), .A2(new_n207), .B1(new_n808), .B2(new_n800), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n1264), .B(new_n1265), .C1(G58), .C2(new_n1040), .ZN(new_n1266));
  OAI221_X1 g1066(.A(new_n1266), .B1(new_n859), .B2(new_n869), .C1(new_n1104), .C2(new_n1176), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n1036), .A2(new_n815), .B1(new_n816), .B2(new_n1043), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n1261), .A2(new_n1263), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  OR2_X1    g1069(.A1(new_n1269), .A2(KEYINPUT119), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n850), .B1(new_n1269), .B2(KEYINPUT119), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1256), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n946), .B2(new_n872), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1255), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(KEYINPUT120), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT120), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1255), .A2(new_n1276), .A3(new_n1273), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n998), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1149), .A2(new_n1152), .A3(new_n1155), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1157), .A2(new_n1279), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1278), .A2(new_n1281), .ZN(G381));
  INV_X1    g1082(.A(KEYINPUT121), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1088), .B(new_n836), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1284), .A2(G384), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1120), .A2(new_n1122), .A3(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(G378), .ZN(new_n1287));
  INV_X1    g1087(.A(G381), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1286), .A2(new_n1287), .A3(new_n1050), .A4(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1283), .B1(new_n1253), .B2(new_n1290), .ZN(new_n1291));
  AOI211_X1 g1091(.A(KEYINPUT121), .B(new_n1289), .C1(new_n1244), .C2(new_n1252), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(G407));
  NAND2_X1  g1094(.A1(new_n1253), .A2(new_n1287), .ZN(new_n1295));
  INV_X1    g1095(.A(G213), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1296), .A2(G343), .ZN(new_n1297));
  XOR2_X1   g1097(.A(new_n1297), .B(KEYINPUT122), .Z(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(G213), .B1(new_n1295), .B2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(KEYINPUT123), .B1(new_n1293), .B2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(G378), .B1(new_n1244), .B2(new_n1252), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1296), .B1(new_n1302), .B2(new_n1298), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT123), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n1303), .B(new_n1304), .C1(new_n1292), .C2(new_n1291), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1301), .A2(new_n1305), .ZN(G409));
  OAI211_X1 g1106(.A(G378), .B(new_n1250), .C1(new_n1251), .C2(new_n1209), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n771), .B1(new_n1206), .B2(KEYINPUT124), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1308), .B1(KEYINPUT124), .B2(new_n1206), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1212), .A2(new_n1279), .A3(new_n1207), .A4(new_n1213), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1309), .A2(new_n1242), .A3(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n1287), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1297), .B1(new_n1307), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT125), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT60), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1280), .B1(new_n1159), .B2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n711), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1149), .A2(new_n1152), .A3(new_n1155), .A4(KEYINPUT60), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1314), .B1(new_n1317), .B2(new_n1319), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1316), .A2(KEYINPUT125), .A3(new_n711), .A4(new_n1318), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1320), .A2(new_n1278), .A3(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(G384), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1320), .A2(G384), .A3(new_n1278), .A4(new_n1321), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1313), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT63), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(G393), .A2(G396), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(new_n1284), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1332), .B1(new_n1122), .B2(new_n1120), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1333), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1332), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1334), .A2(new_n1050), .A3(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1335), .ZN(new_n1337));
  OAI21_X1  g1137(.A(G387), .B1(new_n1337), .B2(new_n1333), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT61), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1336), .A2(new_n1338), .A3(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1298), .B1(new_n1307), .B2(new_n1312), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1326), .A2(new_n1329), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1340), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1343));
  AND2_X1   g1143(.A1(new_n1297), .A2(G2897), .ZN(new_n1344));
  AND3_X1   g1144(.A1(new_n1324), .A2(new_n1325), .A3(new_n1344), .ZN(new_n1345));
  AOI22_X1  g1145(.A1(new_n1324), .A2(new_n1325), .B1(G2897), .B2(new_n1298), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1345), .A2(new_n1346), .ZN(new_n1347));
  OAI211_X1 g1147(.A(new_n1330), .B(new_n1343), .C1(new_n1313), .C2(new_n1347), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1339), .B1(new_n1341), .B2(new_n1347), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT62), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1328), .A2(new_n1350), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1341), .A2(KEYINPUT62), .A3(new_n1327), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1349), .B1(new_n1351), .B2(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1336), .A2(new_n1338), .ZN(new_n1354));
  XNOR2_X1  g1154(.A(new_n1354), .B(KEYINPUT126), .ZN(new_n1355));
  OAI21_X1  g1155(.A(new_n1348), .B1(new_n1353), .B2(new_n1355), .ZN(G405));
  XNOR2_X1  g1156(.A(new_n1354), .B(new_n1326), .ZN(new_n1357));
  OAI21_X1  g1157(.A(G378), .B1(new_n1215), .B2(new_n1243), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1295), .A2(new_n1358), .ZN(new_n1359));
  XNOR2_X1  g1159(.A(new_n1357), .B(new_n1359), .ZN(G402));
endmodule


