//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 1 0 0 0 0 1 1 0 0 0 1 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 0 1 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 1 0 0 0 0 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983;
  INV_X1    g000(.A(KEYINPUT12), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT1), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G128), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  AND3_X1   g007(.A1(new_n193), .A2(KEYINPUT64), .A3(G146), .ZN(new_n194));
  AOI21_X1  g008(.A(KEYINPUT64), .B1(new_n193), .B2(G146), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n189), .B(new_n192), .C1(new_n194), .C2(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n193), .A2(G146), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n198), .B1(new_n188), .B2(G143), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n193), .A2(KEYINPUT64), .A3(G146), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n197), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n190), .B1(G143), .B2(new_n188), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n196), .B1(new_n201), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(G104), .B(G107), .ZN(new_n207));
  INV_X1    g021(.A(G101), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT76), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G104), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT3), .B1(new_n210), .B2(G107), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n213), .A3(G104), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n210), .A2(G107), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n211), .A2(new_n214), .A3(new_n208), .A4(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT76), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n213), .A2(G104), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n210), .A2(G107), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n217), .B(G101), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n209), .A2(new_n216), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT77), .B1(new_n206), .B2(new_n221), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n209), .A2(new_n216), .A3(new_n220), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT77), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n224), .A3(new_n205), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n193), .A2(G146), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n189), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n227), .B1(new_n202), .B2(new_n203), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n196), .A2(new_n228), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n222), .A2(new_n225), .B1(new_n221), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT11), .ZN(new_n231));
  INV_X1    g045(.A(G134), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(G137), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(G137), .ZN(new_n234));
  INV_X1    g048(.A(G137), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(KEYINPUT11), .A3(G134), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n233), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G131), .ZN(new_n238));
  INV_X1    g052(.A(G131), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n233), .A2(new_n236), .A3(new_n239), .A4(new_n234), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n187), .B1(new_n230), .B2(new_n242), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n223), .A2(new_n224), .A3(new_n205), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n224), .B1(new_n223), .B2(new_n205), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n196), .A2(new_n228), .ZN(new_n246));
  OAI22_X1  g060(.A1(new_n244), .A2(new_n245), .B1(new_n223), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(KEYINPUT12), .A3(new_n241), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n243), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT10), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n250), .B1(new_n244), .B2(new_n245), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT78), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n254));
  AND3_X1   g068(.A1(new_n196), .A2(new_n228), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n254), .B1(new_n196), .B2(new_n228), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n221), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n211), .A2(new_n214), .A3(new_n215), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G101), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(KEYINPUT4), .A3(new_n216), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n260), .A2(new_n263), .A3(G101), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT0), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n267), .A2(new_n203), .ZN(new_n268));
  AOI22_X1  g082(.A1(new_n189), .A2(new_n226), .B1(KEYINPUT0), .B2(G128), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n267), .A2(new_n203), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n201), .A2(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n259), .A2(KEYINPUT10), .B1(new_n266), .B2(new_n271), .ZN(new_n272));
  OAI211_X1 g086(.A(KEYINPUT78), .B(new_n250), .C1(new_n244), .C2(new_n245), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n253), .A2(new_n242), .A3(new_n272), .A4(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n249), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT68), .B(G953), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G227), .ZN(new_n277));
  XNOR2_X1  g091(.A(G110), .B(G140), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n277), .B(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n275), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n253), .A2(new_n272), .A3(new_n273), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n241), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(new_n274), .A3(new_n279), .ZN(new_n284));
  AOI21_X1  g098(.A(G902), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G469), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT79), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G902), .ZN(new_n288));
  XNOR2_X1  g102(.A(KEYINPUT80), .B(G469), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n279), .B1(new_n283), .B2(new_n274), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n249), .A2(new_n274), .A3(new_n279), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n288), .B(new_n289), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT79), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n274), .A2(new_n279), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n294), .A2(new_n283), .B1(new_n275), .B2(new_n280), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n293), .B(G469), .C1(new_n295), .C2(G902), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n287), .A2(new_n292), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G221), .ZN(new_n298));
  XOR2_X1   g112(.A(KEYINPUT9), .B(G234), .Z(new_n299));
  AOI21_X1  g113(.A(new_n298), .B1(new_n299), .B2(new_n288), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n235), .A2(G134), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n232), .A2(G137), .ZN(new_n305));
  OAI21_X1  g119(.A(G131), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n240), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n307), .B1(new_n255), .B2(new_n257), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n271), .A2(new_n241), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(KEYINPUT30), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT66), .ZN(new_n311));
  INV_X1    g125(.A(G116), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n311), .B1(new_n312), .B2(G119), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(G119), .ZN(new_n314));
  INV_X1    g128(.A(G119), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(KEYINPUT66), .A3(G116), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n313), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT65), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT2), .B(G113), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n319), .B1(new_n317), .B2(new_n318), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n307), .A2(new_n246), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n309), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT30), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n310), .A2(new_n323), .A3(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n329), .B(G101), .ZN(new_n330));
  INV_X1    g144(.A(G237), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n276), .A2(G210), .A3(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n330), .B(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n308), .A2(new_n322), .A3(new_n309), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n328), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT31), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT28), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n325), .A2(new_n323), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n308), .A2(KEYINPUT28), .A3(new_n322), .A4(new_n309), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n333), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT69), .B(KEYINPUT31), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n328), .A2(new_n333), .A3(new_n334), .A4(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n336), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT70), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(G472), .A2(G902), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n336), .A2(new_n343), .A3(KEYINPUT70), .A4(new_n345), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(KEYINPUT32), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT32), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n348), .A2(new_n353), .A3(new_n349), .A4(new_n350), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n338), .A2(new_n340), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n322), .B1(new_n308), .B2(new_n309), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT71), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT71), .ZN(new_n358));
  INV_X1    g172(.A(new_n334), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(new_n356), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n358), .B1(new_n360), .B2(new_n337), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n357), .A2(new_n361), .A3(KEYINPUT29), .A4(new_n333), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n328), .A2(new_n334), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n342), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT29), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n364), .B(new_n365), .C1(new_n342), .C2(new_n341), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n362), .A2(new_n366), .A3(new_n288), .ZN(new_n367));
  AOI22_X1  g181(.A1(new_n352), .A2(new_n354), .B1(G472), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G125), .ZN(new_n369));
  OR3_X1    g183(.A1(new_n369), .A2(KEYINPUT16), .A3(G140), .ZN(new_n370));
  XOR2_X1   g184(.A(G125), .B(G140), .Z(new_n371));
  INV_X1    g185(.A(KEYINPUT16), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(new_n188), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n203), .A2(G119), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT73), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n375), .B(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n315), .A2(G128), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  XOR2_X1   g193(.A(KEYINPUT24), .B(G110), .Z(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G110), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT23), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n375), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n203), .A2(KEYINPUT23), .A3(G119), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n384), .A2(new_n378), .A3(new_n385), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n374), .B(new_n381), .C1(new_n382), .C2(new_n386), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n384), .A2(new_n385), .A3(new_n382), .A4(new_n378), .ZN(new_n388));
  OR2_X1    g202(.A1(new_n388), .A2(KEYINPUT74), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(KEYINPUT74), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n389), .B(new_n390), .C1(new_n379), .C2(new_n380), .ZN(new_n391));
  OR2_X1    g205(.A1(new_n371), .A2(G146), .ZN(new_n392));
  OR2_X1    g206(.A1(new_n373), .A2(new_n188), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n387), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n276), .A2(G221), .A3(G234), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT22), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n396), .B(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n398), .B(new_n235), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n387), .A3(new_n394), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n288), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT25), .ZN(new_n404));
  INV_X1    g218(.A(G217), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n405), .B1(G234), .B2(new_n288), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n406), .B(KEYINPUT72), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT25), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n401), .A2(new_n408), .A3(new_n288), .A4(new_n402), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n404), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  OR2_X1    g224(.A1(new_n403), .A2(new_n406), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT75), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n412), .B(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n368), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(G214), .B1(G237), .B2(G902), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n262), .B(new_n264), .C1(new_n320), .C2(new_n321), .ZN(new_n417));
  INV_X1    g231(.A(new_n317), .ZN(new_n418));
  INV_X1    g232(.A(new_n319), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n313), .A2(new_n316), .A3(KEYINPUT5), .A4(new_n314), .ZN(new_n420));
  NOR3_X1   g234(.A1(new_n312), .A2(KEYINPUT5), .A3(G119), .ZN(new_n421));
  INV_X1    g235(.A(G113), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n418), .A2(new_n419), .B1(new_n420), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n223), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n417), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(G110), .B(G122), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(KEYINPUT81), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n429), .A2(KEYINPUT6), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n229), .A2(new_n369), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT84), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n431), .B(new_n432), .C1(new_n369), .C2(new_n271), .ZN(new_n433));
  INV_X1    g247(.A(G224), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(G953), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n271), .A2(new_n369), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n246), .A2(G125), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT84), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n433), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n435), .B1(new_n433), .B2(new_n438), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT83), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT82), .ZN(new_n443));
  OAI21_X1  g257(.A(KEYINPUT6), .B1(new_n429), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n417), .A2(new_n425), .A3(new_n427), .ZN(new_n445));
  INV_X1    g259(.A(new_n428), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n446), .B1(new_n417), .B2(new_n425), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n445), .B1(new_n447), .B2(KEYINPUT82), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n442), .B1(new_n444), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n429), .A2(new_n443), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT6), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n451), .B1(new_n447), .B2(KEYINPUT82), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n450), .A2(new_n452), .A3(KEYINPUT83), .A4(new_n445), .ZN(new_n453));
  AOI211_X1 g267(.A(new_n430), .B(new_n441), .C1(new_n449), .C2(new_n453), .ZN(new_n454));
  XOR2_X1   g268(.A(new_n427), .B(KEYINPUT8), .Z(new_n455));
  INV_X1    g269(.A(KEYINPUT85), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n420), .B(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n423), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n418), .A2(new_n419), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n455), .B1(new_n460), .B2(new_n223), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n424), .A2(new_n221), .ZN(new_n462));
  OAI22_X1  g276(.A1(new_n436), .A2(new_n437), .B1(KEYINPUT86), .B2(new_n435), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT7), .B1(new_n434), .B2(G953), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n464), .ZN(new_n466));
  OAI221_X1 g280(.A(new_n466), .B1(KEYINPUT86), .B2(new_n435), .C1(new_n436), .C2(new_n437), .ZN(new_n467));
  AOI22_X1  g281(.A1(new_n461), .A2(new_n462), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n445), .B1(new_n468), .B2(KEYINPUT87), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n465), .A2(new_n467), .ZN(new_n470));
  INV_X1    g284(.A(new_n455), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n457), .A2(new_n423), .B1(new_n419), .B2(new_n418), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n471), .B(new_n462), .C1(new_n472), .C2(new_n221), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT87), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n288), .B1(new_n469), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(G210), .B1(G237), .B2(G902), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NOR3_X1   g293(.A1(new_n454), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n449), .A2(new_n453), .ZN(new_n481));
  INV_X1    g295(.A(new_n430), .ZN(new_n482));
  INV_X1    g296(.A(new_n441), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n445), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n485), .B1(new_n474), .B2(new_n475), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n468), .A2(KEYINPUT87), .ZN(new_n487));
  AOI21_X1  g301(.A(G902), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n478), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n416), .B1(new_n480), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  AND2_X1   g305(.A1(KEYINPUT68), .A2(G953), .ZN(new_n492));
  NOR2_X1   g306(.A1(KEYINPUT68), .A2(G953), .ZN(new_n493));
  OAI211_X1 g307(.A(G214), .B(new_n331), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n193), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n276), .A2(G143), .A3(G214), .A4(new_n331), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(G131), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT17), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n495), .A2(new_n496), .A3(new_n239), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n373), .B(G146), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n497), .A2(KEYINPUT17), .A3(G131), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n371), .A2(G146), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n392), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT18), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n507), .A2(new_n239), .ZN(new_n508));
  OAI221_X1 g322(.A(new_n506), .B1(new_n497), .B2(new_n508), .C1(new_n498), .C2(new_n507), .ZN(new_n509));
  XNOR2_X1  g323(.A(G113), .B(G122), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(new_n210), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n504), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT88), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n504), .A2(new_n509), .A3(KEYINPUT88), .A4(new_n511), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n498), .A2(new_n500), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n371), .B(KEYINPUT19), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n517), .B(new_n393), .C1(G146), .C2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n509), .ZN(new_n520));
  INV_X1    g334(.A(new_n511), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n516), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(G475), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT20), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n525), .A2(KEYINPUT89), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n523), .A2(new_n524), .A3(new_n288), .A4(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n511), .B1(new_n504), .B2(new_n509), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n528), .B1(new_n514), .B2(new_n515), .ZN(new_n529));
  OAI21_X1  g343(.A(G475), .B1(new_n529), .B2(G902), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n514), .A2(new_n515), .B1(new_n521), .B2(new_n520), .ZN(new_n531));
  NOR3_X1   g345(.A1(new_n531), .A2(G475), .A3(G902), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT89), .B(KEYINPUT20), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n527), .B(new_n530), .C1(new_n532), .C2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(G952), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(G953), .ZN(new_n538));
  INV_X1    g352(.A(G234), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n538), .B1(new_n539), .B2(new_n331), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  AOI211_X1 g355(.A(new_n288), .B(new_n276), .C1(G234), .C2(G237), .ZN(new_n542));
  XOR2_X1   g356(.A(KEYINPUT21), .B(G898), .Z(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n541), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(G128), .B(G143), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n547), .B(new_n232), .ZN(new_n548));
  INV_X1    g362(.A(G122), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(G116), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n312), .A2(G122), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n213), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(KEYINPUT14), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT92), .ZN(new_n555));
  OR2_X1    g369(.A1(new_n551), .A2(KEYINPUT14), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT92), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n551), .A2(new_n557), .A3(KEYINPUT14), .ZN(new_n558));
  AND4_X1   g372(.A1(new_n550), .A2(new_n555), .A3(new_n556), .A4(new_n558), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n548), .B(new_n553), .C1(new_n559), .C2(new_n213), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n547), .A2(new_n232), .ZN(new_n561));
  OR2_X1    g375(.A1(new_n561), .A2(KEYINPUT91), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n552), .B(new_n213), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT90), .B(KEYINPUT13), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n547), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n193), .A2(G128), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n565), .B(G134), .C1(new_n566), .C2(new_n564), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n561), .A2(KEYINPUT91), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n562), .A2(new_n563), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n560), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G953), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n299), .A2(G217), .A3(new_n571), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n572), .B(KEYINPUT93), .Z(new_n573));
  NAND2_X1  g387(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n573), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n575), .A2(new_n560), .A3(new_n569), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n574), .A2(new_n576), .A3(KEYINPUT94), .ZN(new_n577));
  OR3_X1    g391(.A1(new_n570), .A2(KEYINPUT94), .A3(new_n573), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n578), .A3(new_n288), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT95), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(G478), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n582), .A2(KEYINPUT15), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n577), .A2(new_n578), .A3(KEYINPUT95), .A4(new_n288), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n581), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  OR2_X1    g399(.A1(new_n579), .A2(new_n583), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n536), .A2(new_n546), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n303), .A2(new_n415), .A3(new_n491), .A4(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(G101), .ZN(G3));
  AND2_X1   g406(.A1(new_n348), .A2(new_n350), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n348), .A2(new_n288), .A3(new_n350), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n593), .A2(new_n349), .B1(new_n594), .B2(G472), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n297), .A2(new_n301), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n414), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n416), .B(new_n546), .C1(new_n480), .C2(new_n489), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n574), .A2(KEYINPUT96), .A3(new_n576), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n570), .A2(KEYINPUT96), .A3(new_n573), .ZN(new_n602));
  OAI21_X1  g416(.A(KEYINPUT33), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT33), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n577), .A2(new_n578), .A3(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n603), .A2(G478), .A3(new_n288), .A4(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n581), .A2(new_n582), .A3(new_n584), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n535), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n600), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n599), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT34), .B(G104), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  AOI21_X1  g427(.A(G475), .B1(new_n516), .B2(new_n522), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n534), .B1(new_n614), .B2(new_n288), .ZN(new_n615));
  INV_X1    g429(.A(new_n526), .ZN(new_n616));
  NOR4_X1   g430(.A1(new_n531), .A2(G475), .A3(G902), .A4(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT97), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n530), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g434(.A(KEYINPUT97), .B(G475), .C1(new_n529), .C2(G902), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n618), .A2(new_n622), .A3(new_n587), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n600), .A2(new_n623), .A3(KEYINPUT98), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT98), .ZN(new_n625));
  INV_X1    g439(.A(new_n416), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n479), .B1(new_n454), .B2(new_n477), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n484), .A2(new_n478), .A3(new_n488), .ZN(new_n628));
  AOI211_X1 g442(.A(new_n626), .B(new_n545), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n623), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n625), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n599), .B1(new_n624), .B2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G107), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  NOR2_X1   g448(.A1(new_n400), .A2(KEYINPUT36), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(new_n395), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n406), .A2(G902), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n410), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n416), .B(new_n639), .C1(new_n480), .C2(new_n489), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n596), .A2(new_n590), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT37), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(new_n382), .ZN(G12));
  NAND2_X1  g458(.A1(new_n352), .A2(new_n354), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n367), .A2(G472), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n641), .A2(new_n647), .A3(new_n301), .A4(new_n297), .ZN(new_n648));
  INV_X1    g462(.A(G900), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n541), .B1(new_n542), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n623), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(new_n203), .ZN(G30));
  XNOR2_X1  g468(.A(new_n650), .B(KEYINPUT39), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n302), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT40), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n535), .A2(new_n587), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n627), .A2(new_n628), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT38), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(G472), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n335), .B1(new_n360), .B2(new_n333), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n663), .B1(new_n664), .B2(new_n288), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n665), .B1(new_n352), .B2(new_n354), .ZN(new_n666));
  NOR4_X1   g480(.A1(new_n662), .A2(new_n626), .A3(new_n639), .A4(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n657), .A2(new_n659), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G143), .ZN(G45));
  INV_X1    g483(.A(KEYINPUT99), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n302), .A2(new_n368), .A3(new_n640), .ZN(new_n671));
  INV_X1    g485(.A(new_n650), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n535), .A2(new_n608), .A3(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n670), .B1(new_n671), .B2(new_n674), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n648), .A2(KEYINPUT99), .A3(new_n673), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT100), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(new_n188), .ZN(G48));
  NAND2_X1  g493(.A1(new_n283), .A2(new_n274), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n280), .ZN(new_n681));
  INV_X1    g495(.A(new_n291), .ZN(new_n682));
  AOI21_X1  g496(.A(G902), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n301), .B(new_n292), .C1(new_n683), .C2(new_n286), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n368), .A2(new_n414), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n610), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT41), .B(G113), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G15));
  OAI21_X1  g502(.A(new_n685), .B1(new_n631), .B2(new_n624), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G116), .ZN(G18));
  NOR2_X1   g504(.A1(new_n368), .A2(new_n589), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n640), .A2(new_n684), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G119), .ZN(G21));
  NOR2_X1   g508(.A1(new_n658), .A2(KEYINPUT101), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT101), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n696), .B1(new_n535), .B2(new_n587), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n695), .A2(new_n490), .A3(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n684), .A2(new_n545), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n594), .A2(G472), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n357), .A2(new_n361), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n336), .B(new_n345), .C1(new_n701), .C2(new_n333), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n349), .ZN(new_n703));
  INV_X1    g517(.A(new_n412), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n700), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n698), .A2(new_n699), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G122), .ZN(G24));
  AND2_X1   g521(.A1(new_n700), .A2(new_n703), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n708), .A2(new_n674), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n692), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G125), .ZN(G27));
  NAND3_X1  g525(.A1(new_n627), .A2(new_n416), .A3(new_n628), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n673), .A2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT102), .ZN(new_n714));
  OAI21_X1  g528(.A(G469), .B1(new_n295), .B2(G902), .ZN(new_n715));
  AOI211_X1 g529(.A(new_n714), .B(new_n300), .C1(new_n715), .C2(new_n292), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n292), .B1(new_n285), .B2(new_n286), .ZN(new_n717));
  AOI21_X1  g531(.A(KEYINPUT102), .B1(new_n717), .B2(new_n301), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n713), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n647), .A2(new_n704), .ZN(new_n720));
  OAI21_X1  g534(.A(KEYINPUT42), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n717), .A2(new_n301), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n714), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n300), .B1(new_n715), .B2(new_n292), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(KEYINPUT102), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT42), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n726), .A2(new_n727), .A3(new_n415), .A4(new_n713), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n721), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(new_n239), .ZN(G33));
  INV_X1    g544(.A(new_n712), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n726), .A2(new_n415), .A3(new_n651), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(KEYINPUT103), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G134), .ZN(G36));
  INV_X1    g548(.A(new_n639), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n595), .A2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT106), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(KEYINPUT43), .B1(new_n536), .B2(KEYINPUT105), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n536), .A2(new_n608), .ZN(new_n740));
  OR2_X1    g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n740), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n738), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT44), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n738), .A2(KEYINPUT44), .A3(new_n743), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n731), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(KEYINPUT107), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n295), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(G469), .ZN(new_n752));
  NAND2_X1  g566(.A1(G469), .A2(G902), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(KEYINPUT46), .A3(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT46), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n755), .B(G469), .C1(new_n751), .C2(G902), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n754), .A2(new_n292), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n301), .ZN(new_n758));
  OR2_X1    g572(.A1(new_n758), .A2(new_n655), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n759), .A2(KEYINPUT104), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(KEYINPUT104), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n749), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G137), .ZN(G39));
  AND3_X1   g578(.A1(new_n757), .A2(KEYINPUT47), .A3(new_n301), .ZN(new_n765));
  AOI21_X1  g579(.A(KEYINPUT47), .B1(new_n757), .B2(new_n301), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n368), .B(new_n414), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n713), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XOR2_X1   g583(.A(new_n769), .B(G140), .Z(G42));
  INV_X1    g584(.A(new_n662), .ZN(new_n771));
  NOR4_X1   g585(.A1(new_n740), .A2(new_n626), .A3(new_n300), .A4(new_n412), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT108), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n772), .A2(new_n773), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n292), .B1(new_n683), .B2(new_n286), .ZN(new_n776));
  XOR2_X1   g590(.A(new_n776), .B(KEYINPUT49), .Z(new_n777));
  NAND4_X1  g591(.A1(new_n774), .A2(new_n666), .A3(new_n775), .A4(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n540), .B1(new_n741), .B2(new_n742), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n779), .A2(new_n705), .ZN(new_n780));
  INV_X1    g594(.A(new_n684), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(new_n491), .A3(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n783));
  INV_X1    g597(.A(new_n779), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n684), .A2(new_n712), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n783), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n779), .A2(KEYINPUT113), .A3(new_n785), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n720), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n791), .A2(KEYINPUT48), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(KEYINPUT48), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n538), .B(new_n782), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  AND4_X1   g608(.A1(new_n541), .A2(new_n785), .A3(new_n597), .A4(new_n666), .ZN(new_n795));
  INV_X1    g609(.A(new_n609), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n765), .A2(new_n766), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n800), .B1(new_n301), .B2(new_n776), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n801), .A2(new_n731), .A3(new_n780), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n779), .A2(new_n662), .A3(new_n781), .A4(new_n705), .ZN(new_n803));
  OAI21_X1  g617(.A(KEYINPUT112), .B1(new_n803), .B2(new_n416), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT50), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT50), .ZN(new_n806));
  OAI211_X1 g620(.A(KEYINPUT112), .B(new_n806), .C1(new_n803), .C2(new_n416), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n789), .A2(new_n639), .A3(new_n708), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n795), .A2(new_n536), .A3(new_n607), .A4(new_n606), .ZN(new_n810));
  XOR2_X1   g624(.A(new_n810), .B(KEYINPUT114), .Z(new_n811));
  NAND4_X1  g625(.A1(new_n802), .A2(new_n808), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT51), .B1(new_n802), .B2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n812), .B(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT116), .B1(new_n799), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n818));
  INV_X1    g632(.A(new_n653), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n819), .B(new_n710), .C1(new_n675), .C2(new_n676), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n717), .A2(new_n301), .A3(new_n735), .A4(new_n672), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT110), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n666), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n724), .A2(KEYINPUT110), .A3(new_n735), .A4(new_n672), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n698), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(KEYINPUT111), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n818), .B1(new_n820), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n710), .B1(new_n652), .B2(new_n648), .ZN(new_n828));
  INV_X1    g642(.A(new_n676), .ZN(new_n829));
  OAI21_X1  g643(.A(KEYINPUT99), .B1(new_n648), .B2(new_n673), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT111), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n825), .B(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n831), .A2(new_n833), .A3(KEYINPUT52), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n827), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n721), .A2(new_n728), .A3(new_n732), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n685), .A2(new_n610), .B1(new_n691), .B2(new_n692), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n689), .A3(new_n706), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n536), .A2(new_n587), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n600), .B1(new_n609), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n596), .A2(new_n840), .A3(new_n597), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n591), .A2(new_n841), .A3(new_n642), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n836), .A2(new_n838), .A3(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n647), .A2(new_n301), .A3(new_n297), .A4(new_n672), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n618), .A2(new_n622), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n844), .A2(new_n587), .A3(new_n845), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n726), .A2(new_n709), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n639), .B(new_n731), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT109), .B1(new_n843), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n838), .A2(new_n842), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n721), .A2(new_n728), .A3(new_n732), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n850), .A2(KEYINPUT109), .A3(new_n851), .A4(new_n848), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n835), .B1(new_n849), .B2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n837), .A2(new_n689), .A3(new_n706), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n591), .A2(new_n841), .A3(new_n642), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n848), .A2(new_n851), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT109), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n861), .A2(new_n852), .B1(new_n827), .B2(new_n834), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT53), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n817), .B1(new_n856), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n859), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n820), .A2(new_n826), .A3(new_n818), .ZN(new_n866));
  AOI21_X1  g680(.A(KEYINPUT52), .B1(new_n831), .B2(new_n833), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n865), .B(KEYINPUT53), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n817), .B(new_n868), .C1(new_n862), .C2(KEYINPUT53), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n794), .A2(new_n798), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT116), .ZN(new_n873));
  INV_X1    g687(.A(new_n814), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n874), .A2(new_n812), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n812), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n872), .B(new_n873), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n816), .A2(new_n871), .A3(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(G952), .A2(G953), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n778), .B1(new_n878), .B2(new_n879), .ZN(G75));
  OAI21_X1  g694(.A(new_n868), .B1(new_n862), .B2(KEYINPUT53), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n882), .A2(new_n288), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(G210), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT56), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n481), .A2(new_n482), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(new_n483), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT55), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n884), .A2(new_n885), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n888), .B1(new_n884), .B2(new_n885), .ZN(new_n890));
  INV_X1    g704(.A(new_n276), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n537), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT117), .Z(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n889), .A2(new_n890), .A3(new_n894), .ZN(G51));
  NOR3_X1   g709(.A1(new_n882), .A2(new_n288), .A3(new_n752), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n753), .B(KEYINPUT118), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT57), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n817), .B1(new_n856), .B2(new_n868), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n898), .B1(new_n899), .B2(new_n870), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n290), .A2(new_n291), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT119), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n896), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT120), .B1(new_n903), .B2(new_n894), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT120), .ZN(new_n905));
  INV_X1    g719(.A(new_n902), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n881), .A2(KEYINPUT54), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n869), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n906), .B1(new_n908), .B2(new_n898), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n905), .B(new_n893), .C1(new_n909), .C2(new_n896), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n904), .A2(new_n910), .ZN(G54));
  NAND3_X1  g725(.A1(new_n883), .A2(KEYINPUT58), .A3(G475), .ZN(new_n912));
  OR2_X1    g726(.A1(new_n912), .A2(new_n523), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n523), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n894), .B1(new_n913), .B2(new_n914), .ZN(G60));
  NAND2_X1  g729(.A1(new_n603), .A2(new_n605), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(G478), .A2(G902), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT59), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n908), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT121), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n919), .B1(new_n864), .B2(new_n870), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n894), .B1(new_n923), .B2(new_n916), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n908), .A2(KEYINPUT121), .A3(new_n917), .A4(new_n919), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n922), .A2(new_n924), .A3(new_n925), .ZN(G63));
  NAND2_X1  g740(.A1(G217), .A2(G902), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT60), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n882), .A2(new_n928), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n401), .A2(new_n402), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n928), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n881), .A2(new_n636), .A3(new_n933), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n934), .A2(new_n893), .ZN(new_n935));
  NAND2_X1  g749(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT123), .Z(new_n937));
  OR2_X1    g751(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n932), .A2(new_n935), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n937), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n935), .A2(new_n938), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n940), .B1(new_n941), .B2(new_n931), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n939), .A2(new_n942), .ZN(G66));
  OAI21_X1  g757(.A(G953), .B1(new_n544), .B2(new_n434), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n850), .B2(new_n891), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n886), .B1(G898), .B2(new_n276), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(G69));
  NAND2_X1  g761(.A1(new_n891), .A2(new_n649), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT126), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n769), .B1(new_n749), .B2(new_n762), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n762), .A2(new_n698), .A3(new_n790), .ZN(new_n951));
  AND4_X1   g765(.A1(new_n831), .A2(new_n950), .A3(new_n851), .A4(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n949), .B1(new_n952), .B2(new_n891), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n310), .A2(new_n327), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(new_n518), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(G227), .A2(G900), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n891), .A2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n955), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT124), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(KEYINPUT62), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n839), .A2(new_n609), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n656), .A2(new_n415), .A3(new_n731), .A4(new_n962), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT125), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n831), .A2(new_n668), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n960), .A2(KEYINPUT62), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n950), .A2(new_n961), .A3(new_n964), .A4(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n959), .B1(new_n969), .B2(new_n891), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n956), .A2(new_n958), .A3(new_n970), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n891), .B(new_n957), .C1(new_n953), .C2(new_n959), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(G72));
  NAND2_X1  g787(.A1(new_n968), .A2(new_n363), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n974), .B(new_n850), .C1(new_n952), .C2(new_n363), .ZN(new_n975));
  NAND2_X1  g789(.A1(G472), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT63), .Z(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT127), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n975), .A2(new_n335), .A3(new_n364), .A4(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n364), .A2(new_n335), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n856), .A2(new_n863), .ZN(new_n981));
  INV_X1    g795(.A(new_n977), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n894), .B1(new_n979), .B2(new_n983), .ZN(G57));
endmodule


