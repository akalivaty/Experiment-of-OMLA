//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0 0 1 0 0 0 1 1 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079;
  INV_X1    g000(.A(KEYINPUT67), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT2), .ZN(new_n188));
  INV_X1    g002(.A(G113), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n187), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  NAND3_X1  g004(.A1(KEYINPUT67), .A2(KEYINPUT2), .A3(G113), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n188), .A2(new_n189), .A3(KEYINPUT66), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT66), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n193), .B1(KEYINPUT2), .B2(G113), .ZN(new_n194));
  AOI22_X1  g008(.A1(new_n190), .A2(new_n191), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(G116), .B(G119), .ZN(new_n196));
  XNOR2_X1  g010(.A(new_n195), .B(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G143), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G146), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n199), .A2(new_n201), .A3(KEYINPUT0), .A4(G128), .ZN(new_n202));
  XNOR2_X1  g016(.A(G143), .B(G146), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT0), .B(G128), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT11), .ZN(new_n206));
  INV_X1    g020(.A(G134), .ZN(new_n207));
  OAI211_X1 g021(.A(KEYINPUT64), .B(new_n206), .C1(new_n207), .C2(G137), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G137), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G134), .ZN(new_n211));
  AOI21_X1  g025(.A(KEYINPUT64), .B1(new_n211), .B2(new_n206), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT65), .B(G137), .ZN(new_n214));
  NAND2_X1  g028(.A1(KEYINPUT11), .A2(G134), .ZN(new_n215));
  OAI22_X1  g029(.A1(new_n214), .A2(new_n215), .B1(G134), .B2(new_n210), .ZN(new_n216));
  OAI21_X1  g030(.A(G131), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n210), .A2(G134), .ZN(new_n218));
  AND2_X1   g032(.A1(KEYINPUT65), .A2(G137), .ZN(new_n219));
  NOR2_X1   g033(.A1(KEYINPUT65), .A2(G137), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n215), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n218), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n206), .B1(new_n207), .B2(G137), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT64), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n208), .ZN(new_n227));
  INV_X1    g041(.A(G131), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n223), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n205), .B1(new_n217), .B2(new_n229), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n223), .A2(new_n227), .A3(new_n228), .ZN(new_n231));
  INV_X1    g045(.A(G128), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n199), .B(new_n201), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n199), .A2(new_n201), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n199), .A2(KEYINPUT1), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n235), .A3(G128), .ZN(new_n236));
  INV_X1    g050(.A(new_n211), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n237), .B1(new_n214), .B2(new_n207), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n233), .B(new_n236), .C1(new_n238), .C2(new_n228), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n231), .A2(new_n239), .ZN(new_n240));
  NOR3_X1   g054(.A1(new_n230), .A2(new_n240), .A3(KEYINPUT30), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT30), .ZN(new_n242));
  INV_X1    g056(.A(new_n205), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n228), .B1(new_n223), .B2(new_n227), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n243), .B1(new_n231), .B2(new_n244), .ZN(new_n245));
  OR2_X1    g059(.A1(new_n238), .A2(new_n228), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n236), .A2(new_n233), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n246), .A2(new_n248), .A3(new_n229), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n242), .B1(new_n245), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n197), .B1(new_n241), .B2(new_n250), .ZN(new_n251));
  XOR2_X1   g065(.A(new_n195), .B(new_n196), .Z(new_n252));
  NAND3_X1  g066(.A1(new_n245), .A2(new_n252), .A3(new_n249), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT69), .B(G953), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT68), .B(G237), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G210), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n257), .B(KEYINPUT27), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT26), .B(G101), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n258), .B(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n251), .A2(new_n253), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT31), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT30), .B1(new_n230), .B2(new_n240), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n245), .A2(new_n242), .A3(new_n249), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n252), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n253), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n268), .A2(KEYINPUT31), .A3(new_n260), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n252), .B1(new_n245), .B2(new_n249), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT28), .B1(new_n267), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT28), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n253), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n253), .A2(KEYINPUT70), .A3(new_n272), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n271), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n259), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n258), .B(new_n278), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n263), .A2(new_n269), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(G472), .A2(G902), .ZN(new_n281));
  XOR2_X1   g095(.A(new_n281), .B(KEYINPUT71), .Z(new_n282));
  OAI21_X1  g096(.A(KEYINPUT32), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n277), .A2(new_n279), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT31), .B1(new_n268), .B2(new_n260), .ZN(new_n285));
  NOR4_X1   g099(.A1(new_n266), .A2(new_n279), .A3(new_n262), .A4(new_n267), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT32), .ZN(new_n288));
  INV_X1    g102(.A(new_n282), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n283), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(KEYINPUT74), .B(G902), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n251), .A2(new_n253), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT29), .B1(new_n294), .B2(new_n279), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n253), .A2(KEYINPUT70), .A3(new_n272), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT70), .B1(new_n253), .B2(new_n272), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n298), .A2(new_n271), .A3(new_n260), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n293), .B1(new_n295), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n270), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n272), .B1(new_n301), .B2(new_n253), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n302), .B1(new_n298), .B2(KEYINPUT72), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT73), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT72), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n305), .B1(new_n296), .B2(new_n297), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n260), .A2(KEYINPUT29), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n303), .A2(new_n304), .A3(new_n306), .A4(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n275), .A2(KEYINPUT72), .A3(new_n276), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n306), .A2(new_n309), .A3(new_n271), .A4(new_n307), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT73), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n300), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G472), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n291), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT79), .ZN(new_n315));
  INV_X1    g129(.A(G217), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n316), .B1(new_n292), .B2(G234), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  AND2_X1   g132(.A1(KEYINPUT69), .A2(G953), .ZN(new_n319));
  NOR2_X1   g133(.A1(KEYINPUT69), .A2(G953), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(G221), .A3(G234), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT22), .B(G137), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n322), .B(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n232), .A2(G119), .ZN(new_n325));
  INV_X1    g139(.A(G119), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G128), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT24), .B(G110), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT23), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n331), .B1(new_n326), .B2(G128), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n232), .A2(KEYINPUT23), .A3(G119), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(new_n327), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n330), .B1(G110), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT16), .ZN(new_n337));
  INV_X1    g151(.A(G140), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n338), .A2(G125), .ZN(new_n339));
  INV_X1    g153(.A(G125), .ZN(new_n340));
  OR2_X1    g154(.A1(KEYINPUT75), .A2(G140), .ZN(new_n341));
  NAND2_X1  g155(.A1(KEYINPUT75), .A2(G140), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n339), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AND2_X1   g159(.A1(KEYINPUT75), .A2(G140), .ZN(new_n346));
  NOR2_X1   g160(.A1(KEYINPUT75), .A2(G140), .ZN(new_n347));
  OAI21_X1  g161(.A(G125), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT76), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n337), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n338), .A2(G125), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n352), .A2(KEYINPUT16), .ZN(new_n353));
  OAI21_X1  g167(.A(G146), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n344), .B(G125), .C1(new_n346), .C2(new_n347), .ZN(new_n355));
  INV_X1    g169(.A(new_n339), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(KEYINPUT75), .B(G140), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n344), .B1(new_n358), .B2(G125), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT16), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n353), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(new_n198), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n336), .B1(new_n354), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT78), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n198), .B1(new_n360), .B2(new_n361), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n356), .A2(new_n351), .A3(new_n198), .ZN(new_n366));
  INV_X1    g180(.A(G110), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n332), .A2(new_n333), .A3(new_n367), .A4(new_n327), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n368), .A2(KEYINPUT77), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n328), .A2(new_n329), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n370), .B1(new_n368), .B2(KEYINPUT77), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n366), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n365), .A2(new_n372), .ZN(new_n373));
  NOR3_X1   g187(.A1(new_n363), .A2(new_n364), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n349), .A2(new_n356), .A3(new_n355), .ZN(new_n375));
  AOI211_X1 g189(.A(G146), .B(new_n353), .C1(new_n375), .C2(KEYINPUT16), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n335), .B1(new_n376), .B2(new_n365), .ZN(new_n377));
  OR2_X1    g191(.A1(new_n369), .A2(new_n371), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n354), .A2(new_n366), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(KEYINPUT78), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n324), .B1(new_n374), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n377), .A2(new_n379), .A3(KEYINPUT78), .ZN(new_n382));
  INV_X1    g196(.A(new_n324), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n381), .A2(new_n292), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT25), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n381), .A2(KEYINPUT25), .A3(new_n292), .A4(new_n384), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n318), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n364), .B1(new_n363), .B2(new_n373), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n383), .B1(new_n390), .B2(new_n382), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n382), .A2(new_n383), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n317), .A2(G902), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n315), .B1(new_n389), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(KEYINPUT25), .B1(new_n393), .B2(new_n292), .ZN(new_n398));
  INV_X1    g212(.A(new_n388), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n317), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(KEYINPUT79), .A3(new_n395), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n314), .A2(new_n397), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G224), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(G953), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n205), .A2(G125), .ZN(new_n405));
  AOI21_X1  g219(.A(G125), .B1(new_n236), .B2(new_n233), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n205), .A2(G125), .ZN(new_n408));
  INV_X1    g222(.A(new_n404), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n408), .B(new_n409), .C1(new_n248), .C2(G125), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n326), .A2(G116), .ZN(new_n412));
  OAI21_X1  g226(.A(G113), .B1(new_n412), .B2(KEYINPUT5), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n196), .A2(KEYINPUT5), .ZN(new_n415));
  AOI22_X1  g229(.A1(new_n195), .A2(new_n196), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT81), .ZN(new_n417));
  INV_X1    g231(.A(G107), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(new_n418), .A3(G104), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT3), .ZN(new_n420));
  INV_X1    g234(.A(G101), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT3), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n417), .A2(new_n422), .A3(new_n418), .A4(G104), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n418), .A2(G104), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n420), .A2(new_n421), .A3(new_n423), .A4(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G104), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n427), .A2(G107), .ZN(new_n428));
  OAI21_X1  g242(.A(G101), .B1(new_n428), .B2(new_n424), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n416), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(G110), .B(G122), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n420), .A2(new_n423), .A3(new_n425), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT82), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT4), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n420), .A2(KEYINPUT82), .A3(new_n423), .A4(new_n425), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n434), .A2(new_n435), .A3(G101), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n197), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n426), .A2(KEYINPUT4), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n421), .B1(new_n432), .B2(new_n433), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n439), .B1(new_n440), .B2(new_n436), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n430), .B(new_n431), .C1(new_n438), .C2(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n430), .B1(new_n438), .B2(new_n441), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT84), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n431), .A2(new_n444), .ZN(new_n445));
  AOI22_X1  g259(.A1(new_n442), .A2(KEYINPUT6), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n443), .A2(KEYINPUT6), .A3(new_n445), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n411), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n426), .A2(new_n429), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n416), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n431), .B(KEYINPUT8), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n413), .B1(new_n415), .B2(KEYINPUT85), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT85), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n196), .A2(new_n453), .A3(KEYINPUT5), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n452), .A2(new_n454), .B1(new_n196), .B2(new_n195), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n450), .B(new_n451), .C1(new_n455), .C2(new_n449), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n404), .A2(KEYINPUT7), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n458), .B1(new_n407), .B2(new_n410), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n405), .A2(new_n406), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n460), .A2(KEYINPUT7), .A3(new_n404), .ZN(new_n461));
  NOR3_X1   g275(.A1(new_n457), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(G902), .B1(new_n462), .B2(new_n442), .ZN(new_n463));
  OAI21_X1  g277(.A(G210), .B1(G237), .B2(G902), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n448), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n464), .B1(new_n448), .B2(new_n463), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(G214), .B1(G237), .B2(G902), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n217), .A2(new_n229), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n426), .A2(new_n233), .A3(new_n236), .A4(new_n429), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n426), .A2(new_n429), .B1(new_n236), .B2(new_n233), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT12), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n472), .B(KEYINPUT12), .C1(new_n474), .C2(new_n475), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n473), .B(KEYINPUT10), .ZN(new_n481));
  INV_X1    g295(.A(new_n472), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n437), .A2(new_n243), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n481), .B(new_n482), .C1(new_n441), .C2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n321), .A2(G227), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(KEYINPUT80), .ZN(new_n487));
  XNOR2_X1  g301(.A(G110), .B(G140), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n487), .B(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT83), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT10), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n473), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n474), .A2(KEYINPUT10), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n494), .B(new_n495), .C1(new_n483), .C2(new_n441), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n492), .B(new_n489), .C1(new_n496), .C2(new_n472), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n483), .A2(new_n441), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n495), .A2(new_n494), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n472), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n492), .B1(new_n484), .B2(new_n489), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n491), .B(G469), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(G469), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n480), .A2(new_n484), .A3(new_n489), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n489), .B1(new_n500), .B2(new_n484), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n504), .B(new_n292), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(G469), .A2(G902), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n503), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT9), .B(G234), .ZN(new_n510));
  OAI21_X1  g324(.A(G221), .B1(new_n510), .B2(G902), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(G237), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT68), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT68), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(G237), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n517), .A2(new_n321), .A3(G214), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n200), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT86), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n517), .A2(new_n321), .A3(G143), .A4(G214), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(KEYINPUT18), .A2(G131), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n523), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n519), .A2(new_n520), .A3(new_n525), .A4(new_n521), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n375), .A2(G146), .ZN(new_n527));
  AOI22_X1  g341(.A1(new_n524), .A2(new_n526), .B1(new_n366), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(G113), .B(G122), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(new_n427), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(G143), .B1(new_n256), .B2(G214), .ZN(new_n532));
  INV_X1    g346(.A(new_n521), .ZN(new_n533));
  OAI21_X1  g347(.A(G131), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n519), .A2(new_n228), .A3(new_n521), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n375), .A2(KEYINPUT19), .ZN(new_n537));
  OR3_X1    g351(.A1(new_n352), .A2(KEYINPUT19), .A3(new_n339), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(new_n198), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n536), .A2(new_n354), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n531), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT20), .ZN(new_n542));
  NOR2_X1   g356(.A1(G475), .A2(G902), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT87), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n542), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(new_n545), .B2(new_n544), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT17), .ZN(new_n548));
  AOI211_X1 g362(.A(new_n548), .B(new_n228), .C1(new_n519), .C2(new_n521), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n519), .A2(new_n228), .A3(new_n521), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n228), .B1(new_n519), .B2(new_n521), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n549), .B1(new_n552), .B2(new_n548), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n376), .A2(new_n365), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n528), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n530), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n541), .B(new_n547), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT88), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n541), .B(new_n543), .C1(new_n555), .C2(new_n556), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(KEYINPUT20), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n534), .A2(new_n548), .A3(new_n535), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n551), .A2(KEYINPUT17), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n561), .A2(new_n362), .A3(new_n354), .A4(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n524), .A2(new_n526), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n527), .A2(new_n366), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n567), .A2(new_n530), .B1(new_n531), .B2(new_n540), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT88), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n569), .A3(new_n547), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n558), .A2(new_n560), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT94), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n200), .A2(KEYINPUT13), .A3(G128), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(KEYINPUT93), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n574), .A2(new_n207), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n200), .A2(G128), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT13), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n232), .A2(G143), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n578), .A2(KEYINPUT93), .A3(new_n573), .A4(new_n579), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n576), .A2(new_n579), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n575), .A2(new_n580), .B1(new_n207), .B2(new_n581), .ZN(new_n582));
  AND2_X1   g396(.A1(KEYINPUT91), .A2(G122), .ZN(new_n583));
  NOR2_X1   g397(.A1(KEYINPUT91), .A2(G122), .ZN(new_n584));
  OAI21_X1  g398(.A(G116), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT92), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g401(.A(KEYINPUT92), .B(G116), .C1(new_n583), .C2(new_n584), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(G116), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(G122), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n418), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n591), .ZN(new_n593));
  AOI211_X1 g407(.A(G107), .B(new_n593), .C1(new_n587), .C2(new_n588), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n582), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n589), .A2(new_n418), .A3(new_n591), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n581), .B(new_n207), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n591), .B(KEYINPUT14), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n598), .B1(new_n587), .B2(new_n588), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n596), .B(new_n597), .C1(new_n599), .C2(new_n418), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n510), .A2(new_n316), .A3(G953), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n595), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n601), .B1(new_n595), .B2(new_n600), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n572), .B(new_n292), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(G478), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n605), .A2(KEYINPUT15), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n604), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(G234), .A2(G237), .ZN(new_n609));
  INV_X1    g423(.A(G953), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(G952), .A3(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(new_n611), .B(KEYINPUT95), .Z(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n293), .A2(new_n254), .A3(new_n609), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT21), .B(G898), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n613), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT89), .B(G475), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n530), .A2(KEYINPUT90), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n563), .A2(new_n566), .A3(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(G902), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n620), .B1(new_n563), .B2(new_n566), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n619), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n608), .A2(new_n618), .A3(new_n625), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n571), .A2(new_n626), .A3(KEYINPUT96), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT96), .ZN(new_n628));
  OR2_X1    g442(.A1(new_n604), .A2(new_n606), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n604), .A2(new_n606), .ZN(new_n630));
  AND4_X1   g444(.A1(new_n618), .A2(new_n625), .A3(new_n629), .A4(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n558), .A2(new_n560), .A3(new_n570), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n628), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n471), .B(new_n512), .C1(new_n627), .C2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n402), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT97), .B(G101), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G3));
  AND2_X1   g451(.A1(new_n401), .A2(new_n397), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n287), .A2(new_n289), .ZN(new_n639));
  OAI21_X1  g453(.A(G472), .B1(new_n280), .B2(new_n293), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n512), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT98), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n448), .A2(new_n463), .A3(new_n643), .A4(new_n464), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n644), .A2(new_n469), .ZN(new_n645));
  INV_X1    g459(.A(new_n464), .ZN(new_n646));
  INV_X1    g460(.A(new_n411), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n442), .A2(KEYINPUT6), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n443), .A2(new_n445), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n443), .A2(KEYINPUT6), .A3(new_n445), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n647), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n459), .A2(new_n461), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n653), .A2(new_n442), .A3(new_n456), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n622), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n646), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n656), .A2(KEYINPUT98), .A3(new_n465), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n645), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n602), .A2(new_n603), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n605), .B1(new_n660), .B2(new_n293), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT33), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n595), .A2(new_n600), .A3(new_n601), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT100), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n595), .A2(new_n600), .A3(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n601), .A2(KEYINPUT99), .ZN(new_n666));
  AOI22_X1  g480(.A1(KEYINPUT100), .A2(new_n663), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n662), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n602), .A2(new_n603), .A3(KEYINPUT33), .ZN(new_n670));
  OAI211_X1 g484(.A(G478), .B(new_n292), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  AOI22_X1  g485(.A1(new_n632), .A2(new_n625), .B1(new_n661), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n659), .A2(new_n618), .A3(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n642), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT34), .B(G104), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G6));
  INV_X1    g490(.A(KEYINPUT101), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n568), .A2(new_n542), .A3(new_n543), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n560), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n624), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n680), .A2(new_n622), .A3(new_n621), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n617), .B1(new_n681), .B2(new_n619), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n629), .A2(new_n630), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n679), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n677), .B1(new_n658), .B2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n684), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n686), .A2(KEYINPUT101), .A3(new_n657), .A4(new_n645), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n642), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT35), .B(G107), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G9));
  OAI21_X1  g505(.A(KEYINPUT96), .B1(new_n571), .B2(new_n626), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n631), .A2(new_n628), .A3(new_n632), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n509), .A2(new_n511), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n377), .A2(new_n379), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT102), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n383), .A2(KEYINPUT36), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n394), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n695), .B1(new_n400), .B2(new_n700), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n640), .A2(new_n639), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n694), .A2(new_n701), .A3(new_n471), .A4(new_n702), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT37), .B(G110), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G12));
  NAND2_X1  g519(.A1(new_n679), .A2(new_n683), .ZN(new_n706));
  INV_X1    g520(.A(G900), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n613), .B1(new_n615), .B2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n625), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n314), .A2(new_n701), .A3(new_n659), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G128), .ZN(G30));
  XOR2_X1   g527(.A(new_n708), .B(KEYINPUT39), .Z(new_n714));
  NAND2_X1  g528(.A1(new_n512), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT40), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n717));
  OR2_X1    g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n268), .A2(new_n279), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n301), .A2(new_n253), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n622), .B1(new_n721), .B2(new_n260), .ZN(new_n722));
  OAI21_X1  g536(.A(G472), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n291), .A2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n400), .A2(new_n700), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n468), .B(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n632), .A2(new_n625), .ZN(new_n730));
  AND4_X1   g544(.A1(new_n683), .A2(new_n729), .A3(new_n469), .A4(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n718), .A2(new_n719), .A3(new_n727), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G143), .ZN(G45));
  NAND2_X1  g547(.A1(new_n671), .A2(new_n661), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n730), .A2(new_n734), .A3(new_n709), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n314), .A2(new_n701), .A3(new_n735), .A4(new_n659), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G146), .ZN(G48));
  OAI21_X1  g551(.A(new_n292), .B1(new_n505), .B2(new_n506), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(G469), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n511), .A3(new_n507), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n314), .A2(new_n397), .A3(new_n401), .A4(new_n741), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n673), .ZN(new_n743));
  XOR2_X1   g557(.A(KEYINPUT41), .B(G113), .Z(new_n744));
  XNOR2_X1  g558(.A(new_n743), .B(new_n744), .ZN(G15));
  INV_X1    g559(.A(KEYINPUT105), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n746), .B1(new_n688), .B2(new_n742), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n401), .A2(new_n397), .ZN(new_n748));
  AOI22_X1  g562(.A1(new_n283), .A2(new_n290), .B1(new_n312), .B2(G472), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n685), .A2(new_n687), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n750), .A2(KEYINPUT105), .A3(new_n751), .A4(new_n741), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n747), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G116), .ZN(G18));
  NOR2_X1   g568(.A1(new_n658), .A2(new_n740), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n314), .A2(new_n694), .A3(new_n755), .A4(new_n726), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G119), .ZN(G21));
  AOI21_X1  g571(.A(new_n260), .B1(new_n303), .B2(new_n306), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n285), .A2(new_n286), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n289), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AND4_X1   g574(.A1(new_n395), .A2(new_n400), .A3(new_n640), .A4(new_n760), .ZN(new_n761));
  AND4_X1   g575(.A1(new_n683), .A2(new_n730), .A3(new_n657), .A4(new_n645), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n740), .A2(new_n617), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G122), .ZN(G24));
  INV_X1    g579(.A(new_n697), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n698), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n697), .B1(KEYINPUT36), .B2(new_n383), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n767), .A2(new_n768), .A3(new_n394), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n640), .B(new_n760), .C1(new_n769), .C2(new_n389), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n735), .A3(new_n755), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G125), .ZN(G27));
  NOR3_X1   g587(.A1(new_n466), .A2(new_n470), .A3(new_n467), .ZN(new_n774));
  AND4_X1   g588(.A1(new_n512), .A2(new_n672), .A3(new_n774), .A4(new_n709), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT42), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n389), .A2(new_n396), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n314), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT42), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n512), .A2(new_n672), .A3(new_n774), .A4(new_n709), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n780), .B1(new_n402), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT106), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT106), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n784), .B(new_n780), .C1(new_n402), .C2(new_n781), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n779), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  XOR2_X1   g600(.A(KEYINPUT107), .B(G131), .Z(new_n787));
  XNOR2_X1  g601(.A(new_n786), .B(new_n787), .ZN(G33));
  INV_X1    g602(.A(KEYINPUT108), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n789), .B1(new_n706), .B2(new_n710), .ZN(new_n790));
  INV_X1    g604(.A(new_n710), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n791), .A2(new_n679), .A3(KEYINPUT108), .A4(new_n683), .ZN(new_n792));
  AND4_X1   g606(.A1(new_n512), .A2(new_n790), .A3(new_n774), .A4(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(new_n314), .A3(new_n638), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G134), .ZN(G36));
  OAI21_X1  g609(.A(new_n491), .B1(new_n501), .B2(new_n502), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n504), .B1(new_n796), .B2(new_n797), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n508), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT46), .ZN(new_n802));
  OR3_X1    g616(.A1(new_n801), .A2(KEYINPUT109), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(KEYINPUT109), .B1(new_n801), .B2(new_n802), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n803), .A2(new_n507), .A3(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT110), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n801), .A2(new_n802), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n803), .A2(KEYINPUT110), .A3(new_n507), .A4(new_n804), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n810), .A2(new_n511), .A3(new_n714), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n769), .A2(new_n389), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n702), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n730), .B1(new_n661), .B2(new_n671), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT43), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n632), .A2(new_n625), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n734), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT43), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(KEYINPUT111), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT111), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n817), .B2(new_n820), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n814), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT44), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n825), .A2(KEYINPUT113), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT113), .B1(new_n825), .B2(new_n826), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT112), .ZN(new_n829));
  OAI211_X1 g643(.A(KEYINPUT44), .B(new_n814), .C1(new_n822), .C2(new_n824), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n829), .B1(new_n830), .B2(new_n774), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n830), .A2(new_n829), .A3(new_n774), .ZN(new_n832));
  OAI221_X1 g646(.A(new_n812), .B1(new_n827), .B2(new_n828), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(G137), .ZN(G39));
  NAND2_X1  g648(.A1(new_n810), .A2(new_n511), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT47), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n810), .A2(KEYINPUT47), .A3(new_n511), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n749), .A2(new_n748), .A3(new_n735), .A4(new_n774), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(G140), .ZN(G42));
  NAND3_X1  g656(.A1(new_n777), .A2(new_n511), .A3(new_n469), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n843), .B(KEYINPUT114), .Z(new_n844));
  INV_X1    g658(.A(new_n739), .ZN(new_n845));
  INV_X1    g659(.A(new_n507), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT49), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OR3_X1    g661(.A1(new_n845), .A2(new_n846), .A3(KEYINPUT49), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n815), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  OR4_X1    g663(.A1(new_n724), .A2(new_n844), .A3(new_n729), .A4(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n821), .A2(new_n612), .ZN(new_n851));
  INV_X1    g665(.A(new_n774), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n852), .A2(new_n740), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n638), .A2(new_n725), .A3(new_n613), .A4(new_n853), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n730), .A2(new_n734), .ZN(new_n856));
  OAI22_X1  g670(.A1(new_n854), .A2(new_n770), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n851), .A2(new_n761), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n729), .A2(new_n469), .A3(new_n740), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT50), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n859), .A2(KEYINPUT50), .A3(new_n860), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n857), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n511), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n739), .A2(new_n866), .A3(new_n507), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n837), .A2(new_n838), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT122), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n858), .A2(new_n852), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n868), .A2(KEYINPUT122), .ZN(new_n872));
  OAI211_X1 g686(.A(KEYINPUT51), .B(new_n865), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n868), .A2(new_n870), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT51), .B1(new_n874), .B2(new_n865), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n854), .A2(new_n778), .ZN(new_n876));
  XOR2_X1   g690(.A(new_n876), .B(KEYINPUT48), .Z(new_n877));
  NAND2_X1  g691(.A1(new_n610), .A2(G952), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n878), .B1(new_n859), .B2(new_n755), .ZN(new_n879));
  INV_X1    g693(.A(new_n672), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n877), .B(new_n879), .C1(new_n880), .C2(new_n855), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n875), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n873), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n756), .B(new_n764), .C1(new_n742), .C2(new_n673), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n753), .A2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n885), .B1(new_n747), .B2(new_n752), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(KEYINPUT121), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n703), .B1(new_n402), .B2(new_n634), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT115), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n542), .B1(new_n568), .B2(new_n543), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n556), .B1(new_n563), .B2(new_n566), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n566), .A2(new_n540), .A3(new_n556), .ZN(new_n898));
  NOR4_X1   g712(.A1(new_n897), .A2(new_n898), .A3(KEYINPUT20), .A4(new_n544), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n608), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n895), .B1(new_n900), .B2(new_n710), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n791), .A2(new_n679), .A3(KEYINPUT115), .A4(new_n608), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n901), .A2(new_n774), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n903), .A2(new_n749), .ZN(new_n904));
  AOI22_X1  g718(.A1(new_n750), .A2(new_n793), .B1(new_n904), .B2(new_n701), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n618), .B(new_n469), .C1(new_n466), .C2(new_n467), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n632), .A2(new_n625), .A3(new_n683), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n906), .B1(new_n880), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n638), .A2(new_n908), .A3(new_n641), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n775), .A2(KEYINPUT116), .A3(new_n771), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT116), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n911), .B1(new_n781), .B2(new_n770), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n894), .A2(new_n905), .A3(new_n909), .A4(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT53), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n786), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n749), .A2(new_n658), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n917), .B(new_n701), .C1(new_n711), .C2(new_n735), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT52), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n695), .A2(new_n708), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n762), .A2(new_n724), .A3(new_n813), .A4(new_n920), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n918), .A2(new_n919), .A3(new_n772), .A4(new_n921), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n772), .A2(new_n921), .A3(new_n736), .A4(new_n712), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(KEYINPUT52), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT118), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n918), .A2(new_n925), .A3(new_n772), .A4(new_n921), .ZN(new_n926));
  XNOR2_X1  g740(.A(KEYINPUT118), .B(KEYINPUT119), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n922), .A2(new_n924), .A3(new_n926), .A4(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n924), .A2(new_n922), .A3(new_n926), .ZN(new_n929));
  INV_X1    g743(.A(new_n927), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n892), .A2(new_n916), .A3(new_n928), .A4(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT54), .ZN(new_n933));
  INV_X1    g747(.A(new_n785), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n638), .A2(new_n775), .A3(new_n314), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n784), .B1(new_n935), .B2(new_n780), .ZN(new_n936));
  OAI22_X1  g750(.A1(new_n934), .A2(new_n936), .B1(new_n778), .B2(new_n776), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n904), .A2(new_n701), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT116), .B1(new_n775), .B2(new_n771), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n781), .A2(new_n770), .A3(new_n911), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n794), .B(new_n938), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n909), .B(new_n703), .C1(new_n402), .C2(new_n634), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n937), .A2(new_n943), .A3(new_n890), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n924), .A2(new_n922), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n915), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n932), .A2(new_n933), .A3(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n786), .A2(new_n914), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n948), .A2(new_n890), .A3(new_n922), .A4(new_n924), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(KEYINPUT53), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT117), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n944), .B(new_n951), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n931), .A2(new_n928), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n915), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n950), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n884), .B(new_n947), .C1(new_n955), .C2(new_n933), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n952), .A2(new_n954), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n957), .A2(KEYINPUT120), .A3(KEYINPUT54), .A4(new_n950), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n883), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(G952), .A2(G953), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n850), .B1(new_n959), .B2(new_n960), .ZN(G75));
  INV_X1    g775(.A(KEYINPUT56), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n932), .A2(new_n946), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n293), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n962), .B1(new_n964), .B2(new_n464), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n446), .A2(new_n447), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n647), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n448), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT55), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n965), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n965), .A2(new_n969), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n321), .A2(G952), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(G51));
  NOR2_X1   g787(.A1(new_n964), .A2(new_n800), .ZN(new_n974));
  INV_X1    g788(.A(new_n505), .ZN(new_n975));
  INV_X1    g789(.A(new_n506), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n508), .B(KEYINPUT57), .Z(new_n978));
  AND3_X1   g792(.A1(new_n932), .A2(new_n933), .A3(new_n946), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n933), .B1(new_n932), .B2(new_n946), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n974), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(KEYINPUT123), .B1(new_n982), .B2(new_n972), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT123), .ZN(new_n984));
  INV_X1    g798(.A(new_n972), .ZN(new_n985));
  INV_X1    g799(.A(new_n977), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n963), .A2(KEYINPUT54), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n947), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n986), .B1(new_n988), .B2(new_n978), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n984), .B(new_n985), .C1(new_n989), .C2(new_n974), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n983), .A2(new_n990), .ZN(G54));
  NAND4_X1  g805(.A1(new_n963), .A2(KEYINPUT58), .A3(G475), .A4(new_n293), .ZN(new_n992));
  INV_X1    g806(.A(new_n568), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n992), .A2(new_n993), .ZN(new_n995));
  NOR3_X1   g809(.A1(new_n994), .A2(new_n995), .A3(new_n972), .ZN(G60));
  INV_X1    g810(.A(new_n988), .ZN(new_n997));
  NAND2_X1  g811(.A1(G478), .A2(G902), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT59), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n999), .B1(new_n669), .B2(new_n670), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n985), .B1(new_n997), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n956), .A2(new_n958), .A3(new_n999), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n669), .A2(new_n670), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1001), .B1(new_n1002), .B2(new_n1003), .ZN(G63));
  INV_X1    g818(.A(KEYINPUT124), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n937), .A2(new_n943), .A3(KEYINPUT53), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1006), .B1(new_n889), .B2(new_n891), .ZN(new_n1007));
  AOI22_X1  g821(.A1(new_n1007), .A2(new_n953), .B1(new_n915), .B2(new_n949), .ZN(new_n1008));
  NAND2_X1  g822(.A1(G217), .A2(G902), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1009), .B(KEYINPUT60), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1005), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(new_n393), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1010), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n963), .A2(KEYINPUT124), .A3(new_n1013), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1011), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(KEYINPUT124), .B1(new_n963), .B2(new_n1013), .ZN(new_n1016));
  AOI211_X1 g830(.A(new_n1005), .B(new_n1010), .C1(new_n932), .C2(new_n946), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n699), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1015), .A2(new_n1018), .A3(new_n985), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT61), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n1015), .A2(new_n1018), .A3(KEYINPUT61), .A4(new_n985), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1021), .A2(new_n1022), .ZN(G66));
  OAI21_X1  g837(.A(G953), .B1(new_n616), .B2(new_n403), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n887), .A2(new_n942), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1024), .B1(new_n1025), .B2(new_n254), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n966), .B1(G898), .B2(new_n321), .ZN(new_n1027));
  XNOR2_X1  g841(.A(new_n1027), .B(KEYINPUT125), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1026), .B(new_n1028), .ZN(G69));
  AOI21_X1  g843(.A(new_n321), .B1(G227), .B2(G900), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n264), .A2(new_n265), .ZN(new_n1031));
  AND2_X1   g845(.A1(new_n537), .A2(new_n538), .ZN(new_n1032));
  XNOR2_X1  g846(.A(new_n1031), .B(new_n1032), .ZN(new_n1033));
  INV_X1    g847(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n1034), .B1(G900), .B2(new_n254), .ZN(new_n1035));
  INV_X1    g849(.A(new_n1035), .ZN(new_n1036));
  NAND4_X1  g850(.A1(new_n812), .A2(new_n314), .A3(new_n777), .A4(new_n762), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n786), .B1(new_n750), .B2(new_n793), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n841), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  AND2_X1   g853(.A1(new_n918), .A2(new_n772), .ZN(new_n1040));
  OAI22_X1  g854(.A1(new_n832), .A2(new_n831), .B1(new_n827), .B2(new_n828), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n1040), .B1(new_n1041), .B2(new_n811), .ZN(new_n1042));
  INV_X1    g856(.A(KEYINPUT126), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n833), .A2(KEYINPUT126), .A3(new_n1040), .ZN(new_n1045));
  AOI21_X1  g859(.A(new_n1039), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g860(.A(new_n1036), .B1(new_n1046), .B2(new_n321), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n672), .B1(new_n683), .B2(new_n818), .ZN(new_n1048));
  NOR4_X1   g862(.A1(new_n402), .A2(new_n715), .A3(new_n1048), .A4(new_n852), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n732), .A2(new_n1040), .ZN(new_n1050));
  INV_X1    g864(.A(KEYINPUT62), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g866(.A1(new_n732), .A2(KEYINPUT62), .A3(new_n1040), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n1049), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g868(.A1(new_n833), .A2(new_n1054), .A3(new_n841), .ZN(new_n1055));
  AOI21_X1  g869(.A(new_n1033), .B1(new_n1055), .B2(new_n321), .ZN(new_n1056));
  OAI21_X1  g870(.A(new_n1030), .B1(new_n1047), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g871(.A(new_n1039), .ZN(new_n1058));
  NOR2_X1   g872(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1059));
  AOI21_X1  g873(.A(KEYINPUT126), .B1(new_n833), .B2(new_n1040), .ZN(new_n1060));
  OAI211_X1 g874(.A(new_n321), .B(new_n1058), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g875(.A1(new_n1061), .A2(new_n1035), .ZN(new_n1062));
  INV_X1    g876(.A(new_n1030), .ZN(new_n1063));
  INV_X1    g877(.A(new_n1056), .ZN(new_n1064));
  NAND3_X1  g878(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g879(.A1(new_n1057), .A2(new_n1065), .ZN(G72));
  NAND2_X1  g880(.A1(new_n268), .A2(new_n279), .ZN(new_n1067));
  NAND2_X1  g881(.A1(new_n1046), .A2(new_n1025), .ZN(new_n1068));
  NAND2_X1  g882(.A1(G472), .A2(G902), .ZN(new_n1069));
  XOR2_X1   g883(.A(new_n1069), .B(KEYINPUT63), .Z(new_n1070));
  AOI21_X1  g884(.A(new_n1067), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g885(.A1(new_n294), .A2(new_n279), .ZN(new_n1072));
  NAND2_X1  g886(.A1(new_n1072), .A2(new_n261), .ZN(new_n1073));
  NAND4_X1  g887(.A1(new_n957), .A2(new_n950), .A3(new_n1070), .A4(new_n1073), .ZN(new_n1074));
  NAND4_X1  g888(.A1(new_n833), .A2(new_n1054), .A3(new_n841), .A4(new_n1025), .ZN(new_n1075));
  NAND3_X1  g889(.A1(new_n1075), .A2(KEYINPUT127), .A3(new_n1070), .ZN(new_n1076));
  NAND2_X1  g890(.A1(new_n1076), .A2(new_n720), .ZN(new_n1077));
  AOI21_X1  g891(.A(KEYINPUT127), .B1(new_n1075), .B2(new_n1070), .ZN(new_n1078));
  OAI211_X1 g892(.A(new_n1074), .B(new_n985), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g893(.A1(new_n1071), .A2(new_n1079), .ZN(G57));
endmodule


