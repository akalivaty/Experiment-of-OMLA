//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0 1 0 1 1 0 1 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  XNOR2_X1  g001(.A(G143), .B(G146), .ZN(new_n188));
  AND2_X1   g002(.A1(KEYINPUT0), .A2(G128), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT65), .B1(new_n193), .B2(G143), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(new_n191), .A3(G146), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n192), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT0), .B(G128), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n190), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  AND2_X1   g015(.A1(KEYINPUT66), .A2(G134), .ZN(new_n202));
  NOR2_X1   g016(.A1(KEYINPUT66), .A2(G134), .ZN(new_n203));
  INV_X1    g017(.A(G137), .ZN(new_n204));
  NOR3_X1   g018(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(G134), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT11), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT11), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n202), .A2(new_n203), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(G137), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n201), .B1(new_n208), .B2(new_n211), .ZN(new_n212));
  OR2_X1    g026(.A1(KEYINPUT66), .A2(G134), .ZN(new_n213));
  NAND2_X1  g027(.A1(KEYINPUT66), .A2(G134), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(G137), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n209), .B1(new_n215), .B2(new_n206), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT66), .B(G134), .ZN(new_n217));
  AOI21_X1  g031(.A(KEYINPUT11), .B1(new_n217), .B2(new_n204), .ZN(new_n218));
  NOR3_X1   g032(.A1(new_n216), .A2(new_n218), .A3(G131), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n200), .B1(new_n212), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G128), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n191), .A2(G146), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n193), .A2(G143), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n221), .B1(new_n224), .B2(KEYINPUT1), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n225), .B1(new_n197), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT69), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n208), .A2(new_n201), .A3(new_n211), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n210), .A2(G137), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n204), .A2(G134), .ZN(new_n231));
  OAI21_X1  g045(.A(G131), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT69), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n233), .B(new_n225), .C1(new_n197), .C2(new_n226), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n228), .A2(new_n229), .A3(new_n232), .A4(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G119), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G116), .ZN(new_n237));
  INV_X1    g051(.A(G116), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G119), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT68), .ZN(new_n241));
  XNOR2_X1  g055(.A(G116), .B(G119), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(KEYINPUT2), .A2(G113), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT67), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(KEYINPUT2), .A3(G113), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(KEYINPUT2), .A2(G113), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n241), .B(new_n244), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n250), .B1(new_n246), .B2(new_n248), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n242), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT70), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n251), .A2(new_n256), .A3(new_n253), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n220), .A2(new_n235), .A3(new_n255), .A4(new_n257), .ZN(new_n258));
  XOR2_X1   g072(.A(KEYINPUT26), .B(G101), .Z(new_n259));
  NOR2_X1   g073(.A1(G237), .A2(G953), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G210), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n259), .B(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n262), .B(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n258), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n229), .A2(new_n232), .A3(new_n227), .ZN(new_n268));
  OAI21_X1  g082(.A(G131), .B1(new_n216), .B2(new_n218), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n199), .B1(new_n229), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n267), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n220), .A2(new_n235), .A3(KEYINPUT30), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n272), .A3(new_n254), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n266), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT31), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n266), .A2(KEYINPUT31), .A3(new_n273), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n254), .B1(new_n268), .B2(new_n270), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n258), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT28), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT28), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n258), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n276), .A2(new_n277), .B1(new_n283), .B2(new_n264), .ZN(new_n284));
  INV_X1    g098(.A(G472), .ZN(new_n285));
  INV_X1    g099(.A(G902), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n187), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n266), .A2(KEYINPUT31), .A3(new_n273), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT31), .B1(new_n266), .B2(new_n273), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n281), .B1(new_n258), .B2(new_n278), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n258), .A2(new_n281), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI22_X1  g107(.A1(new_n289), .A2(new_n290), .B1(new_n293), .B2(new_n265), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n294), .A2(KEYINPUT32), .A3(new_n285), .A4(new_n286), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n288), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n280), .A2(new_n265), .A3(new_n282), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT72), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT29), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT72), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n280), .A2(new_n300), .A3(new_n265), .A4(new_n282), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n273), .A2(new_n258), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n264), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n298), .A2(new_n299), .A3(new_n301), .A4(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n220), .A2(new_n235), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n255), .A2(new_n257), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n281), .B1(new_n307), .B2(new_n258), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n308), .A2(new_n292), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n264), .A2(new_n299), .ZN(new_n310));
  AOI21_X1  g124(.A(G902), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n285), .B1(new_n304), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT73), .B1(new_n296), .B2(new_n312), .ZN(new_n313));
  XOR2_X1   g127(.A(KEYINPUT74), .B(G217), .Z(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n315), .B1(G234), .B2(new_n286), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(KEYINPUT75), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT77), .ZN(new_n318));
  INV_X1    g132(.A(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G125), .ZN(new_n320));
  INV_X1    g134(.A(G125), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G140), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n320), .A2(new_n322), .A3(KEYINPUT16), .ZN(new_n323));
  OR3_X1    g137(.A1(new_n321), .A2(KEYINPUT16), .A3(G140), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n318), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NOR3_X1   g139(.A1(new_n321), .A2(KEYINPUT16), .A3(G140), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n326), .A2(KEYINPUT77), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n193), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n327), .ZN(new_n329));
  XNOR2_X1  g143(.A(G125), .B(G140), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n326), .B1(new_n330), .B2(KEYINPUT16), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n329), .B(G146), .C1(new_n331), .C2(new_n318), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n236), .A2(G128), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n221), .A2(KEYINPUT23), .A3(G119), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n236), .A2(G128), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n334), .B(new_n335), .C1(new_n336), .C2(KEYINPUT23), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G110), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT24), .B(G110), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT76), .B1(new_n236), .B2(G128), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(new_n221), .A3(G119), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(new_n342), .A3(new_n334), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n333), .B(new_n338), .C1(new_n339), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n330), .A2(new_n193), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n339), .ZN(new_n346));
  OAI22_X1  g160(.A1(new_n346), .A2(KEYINPUT78), .B1(G110), .B2(new_n337), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n346), .A2(KEYINPUT78), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n332), .B(new_n345), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(KEYINPUT22), .B(G137), .ZN(new_n351));
  INV_X1    g165(.A(G221), .ZN(new_n352));
  INV_X1    g166(.A(G234), .ZN(new_n353));
  NOR3_X1   g167(.A1(new_n352), .A2(new_n353), .A3(G953), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n351), .B(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n350), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n355), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n344), .A2(new_n349), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(new_n286), .A3(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n359), .A2(new_n360), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n317), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n356), .A2(new_n358), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n286), .B1(new_n315), .B2(G234), .ZN(new_n365));
  XOR2_X1   g179(.A(new_n365), .B(KEYINPUT80), .Z(new_n366));
  OR2_X1    g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n301), .A2(new_n299), .A3(new_n303), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n300), .B1(new_n293), .B2(new_n265), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n311), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G472), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT73), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n373), .A2(new_n374), .A3(new_n288), .A4(new_n295), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n313), .A2(new_n369), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G478), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n377), .A2(KEYINPUT15), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n221), .A2(G143), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT96), .B1(new_n221), .B2(G143), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT96), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(new_n191), .A3(G128), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n380), .A2(new_n382), .A3(KEYINPUT13), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT13), .B1(new_n380), .B2(new_n382), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n379), .B(new_n383), .C1(new_n384), .C2(KEYINPUT97), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n384), .A2(KEYINPUT97), .ZN(new_n386));
  OAI21_X1  g200(.A(G134), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n380), .A2(new_n382), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(new_n210), .A3(new_n379), .ZN(new_n389));
  INV_X1    g203(.A(G122), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G116), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n238), .A2(G122), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n391), .A2(new_n392), .A3(KEYINPUT95), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(KEYINPUT95), .B1(new_n391), .B2(new_n392), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n394), .A2(G107), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G107), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n398), .B1(new_n393), .B2(new_n395), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n387), .A2(new_n389), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT14), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n391), .A2(new_n392), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(G107), .B1(new_n392), .B2(new_n402), .ZN(new_n404));
  INV_X1    g218(.A(new_n389), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n210), .B1(new_n388), .B2(new_n379), .ZN(new_n406));
  OAI221_X1 g220(.A(new_n399), .B1(new_n403), .B2(new_n404), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n401), .A2(new_n407), .ZN(new_n408));
  XOR2_X1   g222(.A(KEYINPUT9), .B(G234), .Z(new_n409));
  INV_X1    g223(.A(G953), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n314), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n411), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n401), .A2(new_n407), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT98), .B1(new_n415), .B2(new_n286), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n401), .A2(new_n407), .A3(new_n413), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n413), .B1(new_n401), .B2(new_n407), .ZN(new_n418));
  OAI211_X1 g232(.A(KEYINPUT98), .B(new_n286), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n378), .B1(new_n416), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT99), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n286), .B1(new_n417), .B2(new_n418), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT98), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n378), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n421), .A2(new_n422), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n378), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n423), .A2(new_n424), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n428), .B1(new_n429), .B2(new_n419), .ZN(new_n430));
  OAI21_X1  g244(.A(KEYINPUT99), .B1(new_n430), .B2(new_n425), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n320), .A2(new_n322), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G146), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n345), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT18), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n437), .A2(new_n201), .ZN(new_n438));
  INV_X1    g252(.A(G237), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(new_n410), .A3(G214), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n440), .A2(new_n191), .ZN(new_n441));
  AOI21_X1  g255(.A(G143), .B1(new_n260), .B2(G214), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n438), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n440), .A2(new_n191), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n260), .A2(G143), .A3(G214), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n444), .B(new_n445), .C1(new_n437), .C2(new_n201), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n436), .A2(new_n443), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT91), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT91), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n443), .A2(new_n436), .A3(new_n446), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G113), .B(G122), .ZN(new_n452));
  INV_X1    g266(.A(G104), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n452), .B(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(G131), .B1(new_n441), .B2(new_n442), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT17), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n444), .A2(new_n201), .A3(new_n445), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT92), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n455), .A2(KEYINPUT92), .A3(new_n456), .A4(new_n457), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g276(.A(KEYINPUT17), .B(G131), .C1(new_n441), .C2(new_n442), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n328), .A2(new_n332), .A3(new_n463), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n451), .B(new_n454), .C1(new_n462), .C2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT93), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n333), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n468), .A2(new_n463), .A3(new_n461), .A4(new_n460), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n469), .A2(KEYINPUT93), .A3(new_n454), .A4(new_n451), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n455), .A2(new_n457), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n434), .B(KEYINPUT19), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n332), .B(new_n472), .C1(G146), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n451), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n454), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(G475), .A2(G902), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n433), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n467), .A2(new_n470), .B1(new_n476), .B2(new_n475), .ZN(new_n481));
  INV_X1    g295(.A(new_n479), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n481), .A2(KEYINPUT20), .A3(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n451), .B1(new_n462), .B2(new_n464), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT94), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n484), .A2(new_n485), .A3(new_n476), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n485), .B1(new_n484), .B2(new_n476), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(G902), .B1(new_n488), .B2(new_n471), .ZN(new_n489));
  INV_X1    g303(.A(G475), .ZN(new_n490));
  OAI22_X1  g304(.A1(new_n480), .A2(new_n483), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n410), .A2(G952), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n492), .B1(new_n353), .B2(new_n439), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT21), .B(G898), .ZN(new_n495));
  AOI211_X1 g309(.A(new_n286), .B(new_n410), .C1(G234), .C2(G237), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NOR3_X1   g311(.A1(new_n432), .A2(new_n491), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G224), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n499), .A2(G953), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n500), .A2(KEYINPUT7), .ZN(new_n501));
  INV_X1    g315(.A(new_n227), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n321), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n199), .A2(G125), .ZN(new_n504));
  AOI211_X1 g318(.A(new_n499), .B(G953), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n504), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n506), .A2(new_n500), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n501), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n501), .B1(new_n503), .B2(new_n504), .ZN(new_n509));
  OAI21_X1  g323(.A(KEYINPUT3), .B1(new_n453), .B2(G107), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT3), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(new_n398), .A3(G104), .ZN(new_n512));
  INV_X1    g326(.A(G101), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n453), .A2(G107), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n510), .A2(new_n512), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT82), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n398), .A2(G104), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n514), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n516), .B1(new_n518), .B2(G101), .ZN(new_n519));
  AOI211_X1 g333(.A(KEYINPUT82), .B(new_n513), .C1(new_n517), .C2(new_n514), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n515), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT83), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT83), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n523), .B(new_n515), .C1(new_n519), .C2(new_n520), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n253), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n240), .A2(KEYINPUT68), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n243), .B1(new_n237), .B2(new_n239), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT5), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(G113), .B1(new_n237), .B2(KEYINPUT5), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n526), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n510), .A2(new_n512), .A3(new_n514), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(G101), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT81), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n515), .A2(KEYINPUT4), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT81), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n533), .A2(new_n537), .A3(G101), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n535), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT4), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n533), .A2(new_n540), .A3(G101), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n541), .B1(new_n251), .B2(new_n253), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n525), .A2(new_n532), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(G110), .B(G122), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n509), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT89), .ZN(new_n546));
  AOI21_X1  g360(.A(KEYINPUT88), .B1(new_n242), .B2(KEYINPUT5), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n547), .A2(new_n530), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n242), .A2(KEYINPUT88), .A3(KEYINPUT5), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n526), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n524), .ZN(new_n551));
  XNOR2_X1  g365(.A(G104), .B(G107), .ZN(new_n552));
  OAI21_X1  g366(.A(KEYINPUT82), .B1(new_n552), .B2(new_n513), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n518), .A2(new_n516), .A3(G101), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n523), .B1(new_n555), .B2(new_n515), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n550), .B1(new_n551), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT5), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n558), .B1(new_n241), .B2(new_n244), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n253), .B1(new_n559), .B2(new_n530), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n521), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  XOR2_X1   g376(.A(new_n544), .B(KEYINPUT8), .Z(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n546), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  AOI211_X1 g379(.A(KEYINPUT89), .B(new_n563), .C1(new_n557), .C2(new_n561), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n508), .B(new_n545), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n544), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n560), .B1(new_n522), .B2(new_n524), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n533), .A2(new_n540), .A3(G101), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n527), .A2(new_n252), .A3(new_n528), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n570), .B1(new_n571), .B2(new_n526), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n533), .A2(new_n537), .A3(G101), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n537), .B1(new_n533), .B2(G101), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n515), .A2(KEYINPUT4), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n568), .B1(new_n569), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n532), .B1(new_n551), .B2(new_n556), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n542), .A2(new_n539), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n544), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n578), .A2(KEYINPUT6), .A3(new_n581), .ZN(new_n582));
  OR2_X1    g396(.A1(new_n505), .A2(new_n507), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT6), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n584), .B(new_n568), .C1(new_n569), .C2(new_n577), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n582), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n567), .A2(new_n586), .A3(new_n286), .ZN(new_n587));
  OAI21_X1  g401(.A(G210), .B1(G237), .B2(G902), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n567), .A2(new_n586), .A3(new_n286), .A4(new_n588), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(KEYINPUT90), .A3(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT90), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n587), .A2(new_n593), .A3(new_n589), .ZN(new_n594));
  OAI21_X1  g408(.A(G214), .B1(G237), .B2(G902), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n592), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n352), .B1(new_n409), .B2(new_n286), .ZN(new_n597));
  XOR2_X1   g411(.A(KEYINPUT86), .B(G469), .Z(new_n598));
  NOR2_X1   g412(.A1(new_n541), .A2(new_n199), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n225), .B1(new_n226), .B2(new_n188), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n600), .B(new_n515), .C1(new_n519), .C2(new_n520), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT10), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n539), .A2(new_n599), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n212), .A2(new_n219), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n551), .A2(new_n556), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n228), .A2(KEYINPUT10), .A3(new_n234), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n603), .B(new_n604), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(G110), .B(G140), .ZN(new_n608));
  INV_X1    g422(.A(G227), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(G953), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n608), .B(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n522), .A2(new_n502), .A3(new_n524), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n601), .ZN(new_n615));
  INV_X1    g429(.A(new_n604), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(KEYINPUT84), .B1(new_n212), .B2(new_n219), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT12), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n615), .A2(new_n616), .A3(new_n620), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n613), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n228), .A2(KEYINPUT10), .A3(new_n234), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n525), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n603), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n616), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n612), .B1(new_n628), .B2(new_n607), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n286), .B(new_n598), .C1(new_n624), .C2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(KEYINPUT87), .ZN(new_n631));
  INV_X1    g445(.A(new_n607), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n604), .B1(new_n626), .B2(new_n603), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n611), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT84), .ZN(new_n635));
  AOI221_X4 g449(.A(new_n604), .B1(new_n635), .B2(new_n619), .C1(new_n614), .C2(new_n601), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n620), .B1(new_n615), .B2(new_n616), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n634), .B1(new_n638), .B2(new_n613), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT87), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n639), .A2(new_n640), .A3(new_n286), .A4(new_n598), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n631), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n632), .B1(new_n622), .B2(new_n623), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n607), .A2(KEYINPUT85), .A3(new_n612), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n628), .ZN(new_n645));
  AOI21_X1  g459(.A(KEYINPUT85), .B1(new_n607), .B2(new_n612), .ZN(new_n646));
  OAI22_X1  g460(.A1(new_n643), .A2(new_n612), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n286), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(G469), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n597), .B1(new_n642), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n498), .A2(new_n596), .A3(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n376), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(new_n513), .ZN(G3));
  OR2_X1    g467(.A1(new_n285), .A2(KEYINPUT100), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n294), .A2(new_n286), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n654), .B1(new_n294), .B2(new_n286), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n655), .A2(new_n368), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n650), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n377), .A2(new_n286), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n660), .B1(new_n423), .B2(G478), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT33), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n662), .B1(new_n414), .B2(KEYINPUT101), .ZN(new_n663));
  XOR2_X1   g477(.A(new_n415), .B(new_n663), .Z(new_n664));
  AOI21_X1  g478(.A(new_n661), .B1(new_n664), .B2(G478), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n491), .A2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n595), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n667), .B1(new_n590), .B2(new_n591), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR4_X1   g483(.A1(new_n658), .A2(new_n497), .A3(new_n666), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT34), .B(G104), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G6));
  OAI21_X1  g486(.A(KEYINPUT103), .B1(new_n489), .B2(new_n490), .ZN(new_n673));
  INV_X1    g487(.A(new_n471), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n484), .A2(new_n476), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(KEYINPUT94), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n484), .A2(new_n485), .A3(new_n476), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n286), .B1(new_n674), .B2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT103), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n679), .A2(new_n680), .A3(G475), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n673), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n682), .B1(new_n431), .B2(new_n427), .ZN(new_n683));
  AOI211_X1 g497(.A(new_n497), .B(new_n667), .C1(new_n590), .C2(new_n591), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n478), .A2(new_n433), .A3(new_n479), .ZN(new_n685));
  OAI21_X1  g499(.A(KEYINPUT20), .B1(new_n481), .B2(new_n482), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT102), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n685), .A2(new_n686), .A3(KEYINPUT102), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n683), .A2(new_n684), .A3(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n692), .A2(new_n658), .ZN(new_n693));
  XNOR2_X1  g507(.A(KEYINPUT35), .B(G107), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G9));
  NOR2_X1   g509(.A1(new_n355), .A2(KEYINPUT36), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n350), .B(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n698), .A2(new_n366), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n359), .B(new_n360), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n699), .B1(new_n700), .B2(new_n317), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n655), .A2(new_n701), .A3(new_n656), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n498), .A2(new_n596), .A3(new_n702), .A4(new_n650), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT37), .B(G110), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G12));
  INV_X1    g519(.A(new_n701), .ZN(new_n706));
  AND4_X1   g520(.A1(new_n313), .A2(new_n375), .A3(new_n650), .A4(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n682), .ZN(new_n708));
  INV_X1    g522(.A(G900), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n496), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n493), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n708), .A2(new_n691), .A3(new_n432), .A4(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT104), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n683), .A2(KEYINPUT104), .A3(new_n691), .A4(new_n711), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n707), .A2(new_n668), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G128), .ZN(G30));
  INV_X1    g531(.A(new_n296), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n307), .A2(new_n264), .A3(new_n258), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n286), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n264), .B1(new_n273), .B2(new_n258), .ZN(new_n721));
  OAI21_X1  g535(.A(G472), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n679), .A2(G475), .ZN(new_n725));
  AOI22_X1  g539(.A1(new_n427), .A2(new_n431), .B1(new_n725), .B2(new_n687), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NOR4_X1   g541(.A1(new_n724), .A2(new_n667), .A3(new_n706), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n711), .B(KEYINPUT39), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n650), .A2(new_n729), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n730), .A2(KEYINPUT40), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(KEYINPUT40), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n592), .A2(new_n594), .ZN(new_n733));
  XOR2_X1   g547(.A(new_n733), .B(KEYINPUT38), .Z(new_n734));
  NAND4_X1  g548(.A1(new_n728), .A2(new_n731), .A3(new_n732), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G143), .ZN(G45));
  NAND3_X1  g550(.A1(new_n491), .A2(new_n665), .A3(new_n711), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n707), .A2(new_n668), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G146), .ZN(G48));
  INV_X1    g554(.A(G469), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n741), .B1(new_n639), .B2(new_n286), .ZN(new_n742));
  AOI211_X1 g556(.A(new_n597), .B(new_n742), .C1(new_n631), .C2(new_n641), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n743), .A2(new_n491), .A3(new_n665), .A4(new_n684), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n376), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g559(.A(KEYINPUT41), .B(G113), .Z(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(G15));
  NAND4_X1  g561(.A1(new_n683), .A2(new_n743), .A3(new_n684), .A4(new_n691), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n376), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n238), .ZN(G18));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n751));
  AOI21_X1  g565(.A(KEYINPUT105), .B1(new_n743), .B2(new_n668), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n742), .B1(new_n631), .B2(new_n641), .ZN(new_n753));
  INV_X1    g567(.A(new_n597), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n753), .A2(KEYINPUT105), .A3(new_n754), .A4(new_n668), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n313), .A2(new_n498), .A3(new_n375), .A4(new_n706), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n751), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  AND4_X1   g573(.A1(new_n313), .A2(new_n375), .A3(new_n498), .A4(new_n706), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT105), .ZN(new_n761));
  INV_X1    g575(.A(new_n742), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n642), .A2(new_n754), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n761), .B1(new_n763), .B2(new_n669), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n755), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n760), .A2(KEYINPUT106), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n759), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G119), .ZN(G21));
  INV_X1    g582(.A(new_n497), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n743), .A2(new_n769), .A3(new_n668), .A4(new_n726), .ZN(new_n770));
  OAI21_X1  g584(.A(G472), .B1(new_n284), .B2(G902), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT107), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT107), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n773), .B(G472), .C1(new_n284), .C2(G902), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n276), .A2(new_n277), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n775), .B1(new_n265), .B2(new_n309), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n776), .A2(new_n285), .A3(new_n286), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n772), .A2(new_n369), .A3(new_n774), .A4(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n770), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(new_n390), .ZN(G24));
  NAND4_X1  g594(.A1(new_n772), .A2(new_n706), .A3(new_n774), .A4(new_n777), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(new_n737), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n782), .B1(new_n752), .B2(new_n756), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT108), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n765), .A2(KEYINPUT108), .A3(new_n782), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G125), .ZN(G27));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n789));
  AOI22_X1  g603(.A1(new_n631), .A2(new_n641), .B1(new_n648), .B2(G469), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT109), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n754), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n642), .A2(new_n791), .A3(new_n649), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n733), .A2(new_n595), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n792), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n313), .A2(new_n369), .A3(new_n375), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n797), .A3(new_n738), .ZN(new_n798));
  XNOR2_X1  g612(.A(KEYINPUT110), .B(KEYINPUT42), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n642), .A2(new_n649), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT109), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n667), .B1(new_n592), .B2(new_n594), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n802), .A2(new_n754), .A3(new_n803), .A4(new_n793), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n373), .A2(new_n288), .A3(new_n295), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n738), .A2(new_n805), .A3(KEYINPUT42), .A4(new_n369), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n789), .B1(new_n800), .B2(new_n808), .ZN(new_n809));
  AOI211_X1 g623(.A(KEYINPUT111), .B(new_n807), .C1(new_n798), .C2(new_n799), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G131), .ZN(G33));
  NAND4_X1  g626(.A1(new_n796), .A2(new_n797), .A3(new_n714), .A4(new_n715), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G134), .ZN(G36));
  INV_X1    g628(.A(KEYINPUT45), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n741), .B1(new_n647), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n816), .B1(new_n815), .B2(new_n647), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT112), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n817), .B(new_n818), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n819), .B(KEYINPUT46), .C1(new_n741), .C2(new_n286), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT113), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n817), .B(KEYINPUT112), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n741), .A2(new_n286), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(KEYINPUT113), .A3(KEYINPUT46), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n642), .B1(new_n825), .B2(KEYINPUT46), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n491), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n665), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT43), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n832), .B(new_n833), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n655), .A2(new_n656), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n835), .A2(new_n706), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n834), .A2(KEYINPUT44), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT44), .B1(new_n834), .B2(new_n836), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n837), .A2(new_n838), .A3(new_n795), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n830), .A2(new_n839), .A3(new_n754), .A4(new_n729), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(G137), .ZN(G39));
  NAND3_X1  g655(.A1(new_n738), .A2(new_n368), .A3(new_n803), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n842), .B1(new_n313), .B2(new_n375), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n828), .B1(new_n822), .B2(new_n826), .ZN(new_n844));
  XNOR2_X1  g658(.A(KEYINPUT114), .B(KEYINPUT47), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n844), .A2(new_n597), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n845), .B1(new_n830), .B2(new_n754), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n843), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT115), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI211_X1 g665(.A(KEYINPUT115), .B(new_n843), .C1(new_n847), .C2(new_n848), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(G140), .ZN(G42));
  NAND2_X1  g668(.A1(new_n724), .A2(new_n369), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n753), .B(KEYINPUT49), .Z(new_n856));
  NAND4_X1  g670(.A1(new_n831), .A2(new_n754), .A3(new_n595), .A4(new_n665), .ZN(new_n857));
  NOR4_X1   g671(.A1(new_n855), .A2(new_n734), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n858), .B(KEYINPUT116), .Z(new_n859));
  INV_X1    g673(.A(KEYINPUT53), .ZN(new_n860));
  AND4_X1   g674(.A1(new_n769), .A2(new_n592), .A3(new_n594), .A4(new_n595), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n421), .A2(new_n426), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n862), .A2(new_n725), .A3(new_n687), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n666), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n861), .A2(new_n650), .A3(new_n657), .A4(new_n864), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n865), .B(new_n703), .C1(new_n376), .C2(new_n651), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT117), .ZN(new_n867));
  OAI22_X1  g681(.A1(new_n376), .A2(new_n744), .B1(new_n770), .B2(new_n778), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(new_n749), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n757), .A2(new_n751), .A3(new_n758), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT106), .B1(new_n760), .B2(new_n765), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n867), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n711), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n682), .A2(new_n862), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n875), .A2(new_n691), .A3(new_n803), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT118), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n875), .A2(KEYINPUT118), .A3(new_n691), .A4(new_n803), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n707), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n796), .A2(new_n782), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n813), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n813), .A2(new_n880), .A3(KEYINPUT119), .A4(new_n881), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n811), .A2(new_n873), .A3(new_n886), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n765), .A2(KEYINPUT108), .A3(new_n782), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT108), .B1(new_n765), .B2(new_n782), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n716), .B(new_n739), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n727), .A2(new_n669), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n891), .A2(new_n723), .A3(new_n701), .A4(new_n711), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n802), .A2(new_n754), .A3(new_n793), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(KEYINPUT52), .B1(new_n890), .B2(new_n894), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n714), .A2(new_n715), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n313), .A2(new_n375), .A3(new_n650), .A4(new_n706), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n897), .A2(new_n669), .ZN(new_n898));
  AOI22_X1  g712(.A1(new_n785), .A2(new_n786), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT52), .ZN(new_n900));
  INV_X1    g714(.A(new_n894), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n899), .A2(new_n900), .A3(new_n739), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n895), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n860), .B1(new_n887), .B2(new_n903), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n895), .A2(new_n902), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT117), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n866), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n866), .A2(new_n906), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n767), .B(new_n869), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n909), .B1(new_n884), .B2(new_n885), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n905), .A2(new_n910), .A3(new_n811), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n899), .A2(new_n900), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n912), .A2(KEYINPUT53), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n904), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT120), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n914), .A2(new_n915), .A3(KEYINPUT54), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n807), .B1(new_n798), .B2(new_n799), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n912), .A2(new_n860), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n905), .A2(new_n910), .A3(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT54), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n904), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n916), .A2(new_n921), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n834), .A2(new_n494), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n795), .A2(new_n763), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OR2_X1    g739(.A1(new_n925), .A2(new_n781), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n855), .A2(new_n493), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n927), .A2(new_n924), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n491), .A2(new_n665), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n931), .A2(KEYINPUT121), .ZN(new_n932));
  OAI21_X1  g746(.A(KEYINPUT51), .B1(new_n931), .B2(KEYINPUT121), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n778), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n923), .A2(new_n935), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n734), .A2(new_n595), .A3(new_n763), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT50), .Z(new_n939));
  OAI21_X1  g753(.A(new_n846), .B1(new_n844), .B2(new_n597), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n830), .A2(new_n754), .A3(new_n845), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n753), .A2(new_n597), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n943), .A2(new_n803), .A3(new_n936), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n934), .A2(new_n939), .A3(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n928), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n492), .B1(new_n946), .B2(new_n666), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n368), .B1(new_n718), .B2(new_n373), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n923), .A2(new_n948), .A3(new_n924), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT48), .Z(new_n950));
  AOI211_X1 g764(.A(new_n947), .B(new_n950), .C1(new_n765), .C2(new_n936), .ZN(new_n951));
  INV_X1    g765(.A(new_n931), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n944), .A2(new_n952), .A3(new_n939), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n945), .B(new_n951), .C1(new_n953), .C2(KEYINPUT51), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n915), .B1(new_n914), .B2(KEYINPUT54), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n922), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(G952), .A2(G953), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n859), .B1(new_n956), .B2(new_n957), .ZN(G75));
  NOR2_X1   g772(.A1(new_n410), .A2(G952), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n904), .A2(new_n919), .ZN(new_n961));
  NAND2_X1  g775(.A1(G210), .A2(G902), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n582), .A2(new_n585), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(new_n583), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT55), .Z(new_n967));
  NOR2_X1   g781(.A1(new_n967), .A2(KEYINPUT56), .ZN(new_n968));
  AOI21_X1  g782(.A(KEYINPUT124), .B1(new_n964), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n962), .B1(new_n904), .B2(new_n919), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT124), .ZN(new_n971));
  INV_X1    g785(.A(new_n968), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n960), .B1(new_n969), .B2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT56), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT122), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n975), .B1(new_n970), .B2(new_n976), .ZN(new_n977));
  AOI211_X1 g791(.A(KEYINPUT122), .B(new_n962), .C1(new_n904), .C2(new_n919), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n967), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(KEYINPUT123), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT123), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n981), .B(new_n967), .C1(new_n977), .C2(new_n978), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n974), .B1(new_n980), .B2(new_n982), .ZN(G51));
  XNOR2_X1  g797(.A(new_n961), .B(new_n920), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n824), .B(KEYINPUT57), .Z(new_n985));
  OAI21_X1  g799(.A(new_n639), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n286), .B1(new_n904), .B2(new_n919), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n823), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n959), .B1(new_n986), .B2(new_n988), .ZN(G54));
  NAND3_X1  g803(.A1(new_n987), .A2(KEYINPUT58), .A3(G475), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n990), .A2(new_n481), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n990), .A2(new_n481), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n991), .A2(new_n992), .A3(new_n959), .ZN(G60));
  XNOR2_X1  g807(.A(new_n659), .B(KEYINPUT59), .ZN(new_n994));
  OR2_X1    g808(.A1(new_n664), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n960), .B1(new_n984), .B2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(new_n994), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n997), .B1(new_n922), .B2(new_n955), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n996), .B1(new_n664), .B2(new_n998), .ZN(G63));
  NAND2_X1  g813(.A1(G217), .A2(G902), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(KEYINPUT60), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n1001), .B1(new_n904), .B2(new_n919), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n1002), .A2(new_n697), .ZN(new_n1003));
  INV_X1    g817(.A(new_n358), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n357), .B1(new_n344), .B2(new_n349), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n960), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  OAI211_X1 g822(.A(KEYINPUT125), .B(new_n960), .C1(new_n1002), .C2(new_n1006), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1008), .B1(KEYINPUT61), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT61), .ZN(new_n1012));
  OAI211_X1 g826(.A(new_n1012), .B(new_n1009), .C1(new_n1003), .C2(new_n1007), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1011), .A2(new_n1013), .ZN(G66));
  OAI21_X1  g828(.A(G953), .B1(new_n495), .B2(new_n499), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1015), .B1(new_n873), .B2(G953), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n965), .B1(G898), .B2(new_n410), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT126), .Z(new_n1018));
  XNOR2_X1  g832(.A(new_n1016), .B(new_n1018), .ZN(G69));
  NAND2_X1  g833(.A1(new_n271), .A2(new_n272), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1020), .B(new_n473), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1022), .B1(new_n609), .B2(G953), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n830), .A2(new_n754), .A3(new_n729), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n891), .A2(new_n948), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n840), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g840(.A1(new_n811), .A2(new_n739), .A3(new_n813), .A4(new_n899), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AND2_X1   g842(.A1(new_n853), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1023), .B1(new_n1029), .B2(G953), .ZN(new_n1030));
  INV_X1    g844(.A(new_n730), .ZN(new_n1031));
  NAND4_X1  g845(.A1(new_n797), .A2(new_n1031), .A3(new_n803), .A4(new_n864), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n840), .A2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g847(.A(new_n1033), .B(KEYINPUT127), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n899), .A2(new_n735), .A3(new_n739), .ZN(new_n1035));
  XOR2_X1   g849(.A(new_n1035), .B(KEYINPUT62), .Z(new_n1036));
  NAND3_X1  g850(.A1(new_n853), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1037), .A2(new_n410), .A3(new_n1022), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n709), .B1(new_n1022), .B2(new_n609), .ZN(new_n1039));
  OAI211_X1 g853(.A(new_n1030), .B(new_n1038), .C1(new_n410), .C2(new_n1039), .ZN(G72));
  NAND2_X1  g854(.A1(G472), .A2(G902), .ZN(new_n1041));
  XOR2_X1   g855(.A(new_n1041), .B(KEYINPUT63), .Z(new_n1042));
  OAI21_X1  g856(.A(new_n1042), .B1(new_n1037), .B2(new_n909), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1043), .A2(new_n721), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n853), .A2(new_n873), .A3(new_n1028), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1045), .A2(new_n1042), .ZN(new_n1046));
  NAND4_X1  g860(.A1(new_n1046), .A2(new_n264), .A3(new_n258), .A4(new_n273), .ZN(new_n1047));
  INV_X1    g861(.A(new_n1042), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n1048), .B1(new_n303), .B2(new_n274), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n959), .B1(new_n914), .B2(new_n1049), .ZN(new_n1050));
  AND3_X1   g864(.A1(new_n1044), .A2(new_n1047), .A3(new_n1050), .ZN(G57));
endmodule


