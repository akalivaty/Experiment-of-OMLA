//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 0 0 0 1 1 0 1 0 1 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n851, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974;
  XOR2_X1   g000(.A(KEYINPUT31), .B(G50gat), .Z(new_n202));
  INV_X1    g001(.A(G228gat), .ZN(new_n203));
  INV_X1    g002(.A(G233gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n207));
  NAND2_X1  g006(.A1(G211gat), .A2(G218gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT22), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G204gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G197gat), .ZN(new_n212));
  INV_X1    g011(.A(G197gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G204gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n210), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G211gat), .ZN(new_n216));
  INV_X1    g015(.A(G218gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT70), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(new_n219), .A3(new_n208), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n215), .B(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n207), .B1(new_n221), .B2(KEYINPUT29), .ZN(new_n222));
  AND2_X1   g021(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT75), .B(G155gat), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT2), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G141gat), .ZN(new_n228));
  INV_X1    g027(.A(G148gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G141gat), .A2(G148gat), .ZN(new_n231));
  AND2_X1   g030(.A1(G155gat), .A2(G162gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(G155gat), .A2(G162gat), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n230), .B(new_n231), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n227), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT73), .ZN(new_n237));
  INV_X1    g036(.A(new_n233), .ZN(new_n238));
  NAND2_X1  g037(.A1(G155gat), .A2(G162gat), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NOR3_X1   g039(.A1(new_n232), .A2(new_n233), .A3(KEYINPUT73), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT2), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT74), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT74), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT2), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n232), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n247));
  OAI22_X1  g046(.A1(new_n240), .A2(new_n241), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n236), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n206), .B1(new_n222), .B2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT78), .B(KEYINPUT3), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n236), .A2(new_n248), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT29), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(new_n221), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT80), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n250), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n208), .ZN(new_n258));
  NOR2_X1   g057(.A1(G211gat), .A2(G218gat), .ZN(new_n259));
  NOR3_X1   g058(.A1(new_n258), .A2(new_n259), .A3(KEYINPUT70), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(new_n215), .ZN(new_n261));
  XNOR2_X1  g060(.A(G197gat), .B(G204gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n220), .A2(new_n210), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT3), .B1(new_n264), .B2(new_n253), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n243), .A2(new_n245), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(new_n239), .ZN(new_n267));
  INV_X1    g066(.A(new_n247), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n238), .A2(new_n237), .A3(new_n239), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT73), .B1(new_n232), .B2(new_n233), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n269), .A2(new_n272), .B1(new_n227), .B2(new_n235), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n205), .B1(new_n265), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n264), .B1(new_n252), .B2(new_n253), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT80), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n218), .A2(new_n208), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n277), .A2(new_n262), .A3(new_n210), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n277), .B1(new_n210), .B2(new_n262), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n253), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI22_X1  g079(.A1(new_n280), .A2(new_n251), .B1(new_n248), .B2(new_n236), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n206), .B1(new_n275), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n257), .A2(new_n276), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(G22gat), .ZN(new_n284));
  INV_X1    g083(.A(G22gat), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n257), .A2(new_n276), .A3(new_n282), .A4(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G78gat), .B(G106gat), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n284), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n287), .B1(new_n284), .B2(new_n286), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n202), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n284), .A2(new_n286), .ZN(new_n291));
  INV_X1    g090(.A(new_n287), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n284), .A2(new_n286), .A3(new_n287), .ZN(new_n294));
  INV_X1    g093(.A(new_n202), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n290), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G8gat), .B(G36gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(G64gat), .B(G92gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(G226gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n301), .A2(new_n204), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT25), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT64), .ZN(new_n305));
  INV_X1    g104(.A(G183gat), .ZN(new_n306));
  INV_X1    g105(.A(G190gat), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(G183gat), .A2(G190gat), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT24), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n313));
  AND4_X1   g112(.A1(new_n308), .A2(new_n311), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(G169gat), .A2(G176gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT23), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT23), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n317), .B1(G169gat), .B2(G176gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(G169gat), .A2(G176gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n316), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n304), .B1(new_n314), .B2(new_n320), .ZN(new_n321));
  AND4_X1   g120(.A1(KEYINPUT25), .A2(new_n316), .A3(new_n318), .A4(new_n319), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT65), .ZN(new_n323));
  OAI211_X1 g122(.A(G183gat), .B(G190gat), .C1(new_n323), .C2(KEYINPUT24), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n309), .A2(KEYINPUT65), .A3(new_n310), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n324), .B(new_n325), .C1(G183gat), .C2(G190gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n306), .A2(KEYINPUT27), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT27), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(G183gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n328), .A2(new_n330), .A3(new_n307), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT28), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT27), .B(G183gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n334), .A2(KEYINPUT28), .A3(new_n307), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT26), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n319), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n338), .B1(G169gat), .B2(G176gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n315), .A2(new_n337), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n339), .A2(new_n340), .B1(G183gat), .B2(G190gat), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n321), .A2(new_n327), .B1(new_n336), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n303), .B1(new_n342), .B2(KEYINPUT29), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT71), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n344), .B1(new_n342), .B2(new_n303), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n308), .A2(new_n311), .A3(new_n312), .A4(new_n313), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n346), .A2(new_n316), .A3(new_n318), .A4(new_n319), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n347), .A2(new_n304), .B1(new_n326), .B2(new_n322), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n336), .A2(new_n341), .ZN(new_n349));
  OAI211_X1 g148(.A(KEYINPUT71), .B(new_n302), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n343), .A2(new_n345), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(new_n221), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n302), .B1(new_n348), .B2(new_n349), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n343), .A2(new_n353), .A3(new_n264), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n352), .A2(KEYINPUT72), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT72), .B1(new_n352), .B2(new_n354), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n300), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n300), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n352), .A2(new_n354), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT30), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT30), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n352), .A2(new_n361), .A3(new_n354), .A4(new_n358), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n357), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(KEYINPUT82), .B(KEYINPUT40), .ZN(new_n365));
  NAND2_X1  g164(.A1(G225gat), .A2(G233gat), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n267), .A2(new_n268), .B1(new_n270), .B2(new_n271), .ZN(new_n368));
  INV_X1    g167(.A(G155gat), .ZN(new_n369));
  AND2_X1   g168(.A1(new_n369), .A2(KEYINPUT75), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(KEYINPUT75), .ZN(new_n371));
  OAI22_X1  g170(.A1(new_n370), .A2(new_n371), .B1(new_n224), .B2(new_n223), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n234), .B1(new_n372), .B2(KEYINPUT2), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT3), .B1(new_n368), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(G120gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(G113gat), .ZN(new_n376));
  INV_X1    g175(.A(G113gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(G120gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G127gat), .B(G134gat), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT1), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n380), .B1(new_n381), .B2(new_n379), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT77), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n379), .A2(new_n381), .ZN(new_n386));
  INV_X1    g185(.A(new_n380), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT77), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n388), .A2(new_n389), .A3(new_n382), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n374), .A2(new_n252), .A3(new_n385), .A4(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n383), .A2(new_n384), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n273), .A2(new_n392), .A3(KEYINPUT4), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT66), .B1(new_n383), .B2(new_n384), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT66), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n388), .A2(new_n396), .A3(new_n382), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT4), .B1(new_n398), .B2(new_n273), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n367), .B1(new_n394), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n249), .A2(new_n385), .A3(new_n390), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n273), .A2(new_n392), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(new_n402), .A3(new_n366), .ZN(new_n403));
  OR2_X1    g202(.A1(new_n403), .A2(KEYINPUT81), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT39), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n405), .B1(new_n403), .B2(KEYINPUT81), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n400), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n405), .B(new_n367), .C1(new_n394), .C2(new_n399), .ZN(new_n408));
  XNOR2_X1  g207(.A(G1gat), .B(G29gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(KEYINPUT0), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(KEYINPUT79), .ZN(new_n411));
  XNOR2_X1  g210(.A(G57gat), .B(G85gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n408), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n365), .B1(new_n407), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT83), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n400), .A2(new_n404), .A3(new_n406), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n419), .A2(KEYINPUT40), .A3(new_n414), .A4(new_n408), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT4), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n421), .B1(new_n398), .B2(new_n273), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n402), .A2(KEYINPUT4), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n391), .B(new_n366), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT5), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n401), .A2(new_n402), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n425), .B1(new_n426), .B2(new_n367), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n399), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n367), .A2(KEYINPUT5), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n429), .A2(new_n391), .A3(new_n393), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n413), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n420), .A2(new_n433), .ZN(new_n434));
  OAI211_X1 g233(.A(KEYINPUT83), .B(new_n365), .C1(new_n407), .C2(new_n415), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n364), .A2(new_n418), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT38), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT37), .B1(new_n355), .B2(new_n356), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT37), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n352), .A2(new_n439), .A3(new_n354), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n440), .A2(new_n300), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n437), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT6), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n428), .A2(new_n431), .A3(new_n414), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n433), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n351), .A2(new_n264), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n343), .A2(new_n221), .A3(new_n353), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(KEYINPUT37), .A3(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n440), .A2(new_n448), .A3(new_n437), .A4(new_n300), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n432), .A2(KEYINPUT6), .A3(new_n413), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n445), .A2(new_n449), .A3(new_n450), .A4(new_n359), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n297), .B(new_n436), .C1(new_n442), .C2(new_n451), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n383), .A2(new_n384), .A3(KEYINPUT66), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n396), .B1(new_n388), .B2(new_n382), .ZN(new_n454));
  OAI22_X1  g253(.A1(new_n348), .A2(new_n349), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n321), .A2(new_n327), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n336), .A2(new_n341), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n456), .A2(new_n395), .A3(new_n397), .A4(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(G227gat), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n459), .A2(new_n204), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n455), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  XOR2_X1   g260(.A(KEYINPUT67), .B(KEYINPUT33), .Z(new_n462));
  INV_X1    g261(.A(KEYINPUT32), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(G15gat), .B(G43gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(KEYINPUT68), .ZN(new_n467));
  XNOR2_X1  g266(.A(G71gat), .B(G99gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n467), .B(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT69), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n463), .B1(new_n469), .B2(new_n462), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n461), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n471), .B1(new_n461), .B2(new_n472), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n470), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n460), .B1(new_n455), .B2(new_n458), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT34), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI211_X1 g278(.A(KEYINPUT34), .B(new_n460), .C1(new_n455), .C2(new_n458), .ZN(new_n480));
  OR2_X1    g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n479), .A2(new_n480), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n461), .A2(new_n472), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT69), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n473), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n483), .B1(new_n486), .B2(new_n470), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT36), .B1(new_n482), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n476), .A2(new_n481), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n486), .A2(new_n483), .A3(new_n470), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT36), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n357), .A2(new_n363), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n445), .A2(new_n450), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n290), .A2(new_n296), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n493), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n452), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n482), .A2(new_n487), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n500), .A2(new_n290), .A3(new_n296), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n364), .B1(new_n450), .B2(new_n445), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT35), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT35), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n500), .A2(new_n290), .A3(new_n296), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n504), .B1(new_n496), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT84), .B1(new_n499), .B2(new_n507), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n503), .A2(new_n506), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT84), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n452), .A2(new_n498), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  XOR2_X1   g312(.A(G57gat), .B(G64gat), .Z(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT9), .ZN(new_n515));
  XNOR2_X1  g314(.A(G71gat), .B(G78gat), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n519), .A2(KEYINPUT92), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n519), .A2(KEYINPUT92), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n516), .B(new_n514), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT93), .B(KEYINPUT21), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(G231gat), .A2(G233gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n525), .B(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(G127gat), .B(G155gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n530));
  OR2_X1    g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n530), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(G8gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(G15gat), .B(G22gat), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n535), .A2(G1gat), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT89), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT16), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n535), .B1(new_n539), .B2(G1gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n538), .B(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n523), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n542), .B1(KEYINPUT21), .B2(new_n543), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n533), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n533), .A2(new_n544), .ZN(new_n546));
  XNOR2_X1  g345(.A(G183gat), .B(G211gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT94), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n548), .B1(new_n545), .B2(new_n546), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G190gat), .B(G218gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT95), .B(G85gat), .ZN(new_n554));
  INV_X1    g353(.A(G92gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(G99gat), .A2(G106gat), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n558), .B1(KEYINPUT8), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n556), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  OR2_X1    g360(.A1(G99gat), .A2(G106gat), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n561), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n559), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n556), .A2(new_n560), .A3(new_n564), .A4(new_n557), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT96), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n563), .A2(new_n565), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT96), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G43gat), .B(G50gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT15), .ZN(new_n573));
  NAND2_X1  g372(.A1(G29gat), .A2(G36gat), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT14), .ZN(new_n575));
  INV_X1    g374(.A(G29gat), .ZN(new_n576));
  INV_X1    g375(.A(G36gat), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n573), .B1(new_n574), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n579), .A2(KEYINPUT87), .ZN(new_n583));
  MUX2_X1   g382(.A(KEYINPUT87), .B(new_n583), .S(new_n578), .Z(new_n584));
  OR2_X1    g383(.A1(new_n572), .A2(KEYINPUT15), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n584), .A2(new_n573), .A3(new_n585), .A4(new_n574), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT88), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n585), .A2(new_n573), .A3(new_n574), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT88), .B1(new_n589), .B2(new_n584), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n582), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT17), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n586), .A2(new_n587), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n589), .A2(KEYINPUT88), .A3(new_n584), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n581), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT17), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n571), .B1(new_n592), .B2(new_n597), .ZN(new_n598));
  AND2_X1   g397(.A1(G232gat), .A2(G233gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT41), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n568), .A2(new_n570), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n600), .B1(new_n601), .B2(new_n595), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n553), .B1(new_n598), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n595), .A2(new_n596), .ZN(new_n604));
  AOI211_X1 g403(.A(KEYINPUT17), .B(new_n581), .C1(new_n593), .C2(new_n594), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n601), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI22_X1  g405(.A1(new_n571), .A2(new_n591), .B1(KEYINPUT41), .B2(new_n599), .ZN(new_n607));
  INV_X1    g406(.A(new_n553), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT97), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n603), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT98), .ZN(new_n612));
  XOR2_X1   g411(.A(G134gat), .B(G162gat), .Z(new_n613));
  NOR2_X1   g412(.A1(new_n599), .A2(KEYINPUT41), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n611), .A2(new_n612), .A3(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n612), .B1(new_n611), .B2(new_n615), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n603), .A2(new_n609), .ZN(new_n619));
  OAI22_X1  g418(.A1(new_n617), .A2(new_n618), .B1(new_n610), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n611), .A2(new_n615), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT98), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n619), .A2(new_n610), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n622), .A2(new_n623), .A3(new_n616), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n552), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n538), .B(new_n541), .Z(new_n628));
  OAI21_X1  g427(.A(new_n628), .B1(new_n604), .B2(new_n605), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n591), .A2(new_n542), .ZN(new_n630));
  NAND2_X1  g429(.A1(G229gat), .A2(G233gat), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT18), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n629), .A2(KEYINPUT18), .A3(new_n630), .A4(new_n631), .ZN(new_n635));
  OAI21_X1  g434(.A(KEYINPUT90), .B1(new_n595), .B2(new_n628), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n595), .A2(new_n628), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n595), .A2(KEYINPUT90), .A3(new_n628), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n631), .B(KEYINPUT13), .Z(new_n641));
  AOI21_X1  g440(.A(KEYINPUT91), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT91), .ZN(new_n643));
  INV_X1    g442(.A(new_n641), .ZN(new_n644));
  AOI211_X1 g443(.A(new_n643), .B(new_n644), .C1(new_n638), .C2(new_n639), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n634), .B(new_n635), .C1(new_n642), .C2(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(G113gat), .B(G141gat), .Z(new_n647));
  XNOR2_X1  g446(.A(G169gat), .B(G197gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n649), .B(new_n650), .Z(new_n651));
  XOR2_X1   g450(.A(KEYINPUT86), .B(KEYINPUT12), .Z(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n646), .A2(new_n653), .ZN(new_n654));
  AND3_X1   g453(.A1(new_n595), .A2(KEYINPUT90), .A3(new_n628), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n655), .B1(new_n637), .B2(new_n636), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n643), .B1(new_n656), .B2(new_n644), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n640), .A2(KEYINPUT91), .A3(new_n641), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n653), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n659), .A2(new_n660), .A3(new_n634), .A4(new_n635), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n654), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT10), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n566), .A2(new_n523), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n569), .A2(new_n543), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n568), .A2(KEYINPUT10), .A3(new_n543), .A4(new_n570), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(G230gat), .A2(G233gat), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OR3_X1    g469(.A1(new_n664), .A2(new_n669), .A3(new_n665), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g471(.A(G120gat), .B(G148gat), .Z(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT99), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n674), .B(KEYINPUT100), .Z(new_n675));
  XOR2_X1   g474(.A(G176gat), .B(G204gat), .Z(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT101), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n675), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n672), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n678), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n670), .A2(new_n671), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  AND4_X1   g482(.A1(new_n513), .A2(new_n627), .A3(new_n662), .A4(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n495), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(G1gat), .ZN(G1324gat));
  INV_X1    g486(.A(new_n684), .ZN(new_n688));
  OAI21_X1  g487(.A(G8gat), .B1(new_n688), .B2(new_n494), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(KEYINPUT42), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT16), .B(G8gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT102), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n688), .A2(new_n494), .A3(new_n692), .ZN(new_n693));
  MUX2_X1   g492(.A(new_n690), .B(KEYINPUT42), .S(new_n693), .Z(G1325gat));
  INV_X1    g493(.A(new_n493), .ZN(new_n695));
  OAI21_X1  g494(.A(G15gat), .B1(new_n688), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(G15gat), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n684), .A2(new_n697), .A3(new_n500), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(G1326gat));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n497), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT103), .ZN(new_n701));
  XNOR2_X1  g500(.A(KEYINPUT43), .B(G22gat), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1327gat));
  INV_X1    g502(.A(new_n662), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n551), .A2(new_n704), .A3(new_n682), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n513), .A2(new_n626), .A3(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n707), .A2(new_n576), .A3(new_n685), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT45), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n710), .B1(new_n513), .B2(new_n626), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n710), .B(new_n626), .C1(new_n499), .C2(new_n507), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(KEYINPUT104), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n511), .A2(new_n506), .A3(new_n503), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT104), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n714), .A2(new_n715), .A3(new_n710), .A4(new_n626), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n705), .B1(new_n711), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT105), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n720), .B(new_n705), .C1(new_n711), .C2(new_n717), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n719), .A2(new_n685), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n709), .B1(new_n722), .B2(new_n576), .ZN(G1328gat));
  NAND3_X1  g522(.A1(new_n719), .A2(new_n364), .A3(new_n721), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT106), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT106), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n719), .A2(new_n726), .A3(new_n364), .A4(new_n721), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n725), .A2(G36gat), .A3(new_n727), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n706), .A2(G36gat), .A3(new_n494), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT46), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(G1329gat));
  OAI211_X1 g530(.A(new_n493), .B(new_n705), .C1(new_n711), .C2(new_n717), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(G43gat), .ZN(new_n733));
  INV_X1    g532(.A(G43gat), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n500), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(KEYINPUT47), .B1(new_n706), .B2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT107), .B1(new_n733), .B2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT107), .ZN(new_n739));
  AOI211_X1 g538(.A(new_n739), .B(new_n736), .C1(new_n732), .C2(G43gat), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n719), .A2(new_n493), .A3(new_n721), .ZN(new_n742));
  INV_X1    g541(.A(new_n735), .ZN(new_n743));
  AOI22_X1  g542(.A1(new_n742), .A2(G43gat), .B1(new_n707), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n741), .B1(new_n744), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g544(.A(G50gat), .B1(new_n718), .B2(new_n297), .ZN(new_n746));
  OR2_X1    g545(.A1(new_n297), .A2(G50gat), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n706), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n706), .A2(KEYINPUT108), .A3(new_n747), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n746), .B(KEYINPUT48), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n719), .A2(new_n497), .A3(new_n721), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n748), .B1(new_n753), .B2(G50gat), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n752), .B1(new_n754), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR4_X1   g554(.A1(new_n552), .A2(new_n626), .A3(new_n662), .A4(new_n683), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n714), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(new_n495), .ZN(new_n758));
  XNOR2_X1  g557(.A(KEYINPUT109), .B(G57gat), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(G1332gat));
  AOI211_X1 g559(.A(new_n494), .B(new_n757), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n761));
  NOR2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(G1333gat));
  OAI21_X1  g562(.A(G71gat), .B1(new_n757), .B2(new_n695), .ZN(new_n764));
  INV_X1    g563(.A(G71gat), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n500), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n764), .B1(new_n757), .B2(new_n766), .ZN(new_n767));
  XOR2_X1   g566(.A(new_n767), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g567(.A1(new_n757), .A2(new_n297), .ZN(new_n769));
  XNOR2_X1  g568(.A(KEYINPUT110), .B(G78gat), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n769), .B(new_n770), .ZN(G1335gat));
  AOI21_X1  g570(.A(new_n625), .B1(new_n509), .B2(new_n511), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n551), .A2(new_n662), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n772), .A2(KEYINPUT51), .A3(new_n773), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n778), .A2(new_n685), .A3(new_n554), .A4(new_n682), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n773), .A2(new_n682), .ZN(new_n780));
  INV_X1    g579(.A(new_n711), .ZN(new_n781));
  INV_X1    g580(.A(new_n717), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n783), .A2(new_n784), .A3(new_n685), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n784), .B1(new_n783), .B2(new_n685), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n779), .B1(new_n787), .B2(new_n554), .ZN(G1336gat));
  NAND3_X1  g587(.A1(new_n364), .A2(new_n682), .A3(new_n555), .ZN(new_n789));
  XOR2_X1   g588(.A(new_n789), .B(KEYINPUT112), .Z(new_n790));
  AOI21_X1  g589(.A(KEYINPUT52), .B1(new_n778), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n783), .A2(new_n364), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n791), .B1(new_n793), .B2(new_n555), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT113), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n777), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(new_n776), .ZN(new_n797));
  AOI22_X1  g596(.A1(new_n792), .A2(G92gat), .B1(new_n790), .B2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n794), .B1(new_n798), .B2(new_n799), .ZN(G1337gat));
  NOR2_X1   g599(.A1(new_n683), .A2(G99gat), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n778), .A2(new_n500), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n783), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT114), .B1(new_n803), .B2(new_n695), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(G99gat), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n803), .A2(KEYINPUT114), .A3(new_n695), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n802), .B1(new_n805), .B2(new_n806), .ZN(G1338gat));
  NAND2_X1  g606(.A1(new_n783), .A2(new_n497), .ZN(new_n808));
  XOR2_X1   g607(.A(KEYINPUT115), .B(G106gat), .Z(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n297), .A2(G106gat), .A3(new_n683), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT53), .B1(new_n778), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  AOI22_X1  g612(.A1(new_n808), .A2(new_n809), .B1(new_n797), .B2(new_n811), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(G1339gat));
  INV_X1    g615(.A(new_n651), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n640), .A2(new_n641), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n631), .B1(new_n629), .B2(new_n630), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n661), .A2(new_n682), .A3(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823));
  INV_X1    g622(.A(new_n669), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n666), .A2(new_n824), .A3(new_n667), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n670), .A2(KEYINPUT54), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n678), .B1(new_n670), .B2(KEYINPUT54), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n823), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n824), .B1(new_n666), .B2(new_n667), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n680), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n670), .A2(KEYINPUT54), .A3(new_n825), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n831), .A2(new_n832), .A3(KEYINPUT55), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n828), .A2(new_n681), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n834), .B1(new_n654), .B2(new_n661), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n622), .A2(new_n623), .A3(new_n616), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n623), .B1(new_n622), .B2(new_n616), .ZN(new_n837));
  OAI22_X1  g636(.A1(new_n822), .A2(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n661), .A2(new_n820), .ZN(new_n839));
  INV_X1    g638(.A(new_n834), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n620), .A2(new_n839), .A3(new_n624), .A4(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n551), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  AND4_X1   g641(.A1(new_n551), .A2(new_n625), .A3(new_n704), .A4(new_n683), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n844), .A2(new_n495), .A3(new_n364), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n501), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(new_n704), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(new_n377), .ZN(G1340gat));
  NOR2_X1   g647(.A1(new_n846), .A2(new_n683), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(new_n375), .ZN(G1341gat));
  NOR2_X1   g649(.A1(new_n846), .A2(new_n552), .ZN(new_n851));
  XOR2_X1   g650(.A(new_n851), .B(G127gat), .Z(G1342gat));
  NAND2_X1  g651(.A1(new_n845), .A2(new_n626), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT56), .ZN(new_n854));
  INV_X1    g653(.A(G134gat), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n501), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OR3_X1    g655(.A1(new_n853), .A2(KEYINPUT116), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT116), .B1(new_n853), .B2(new_n856), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n854), .A2(new_n855), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n857), .A2(new_n854), .A3(new_n855), .A4(new_n858), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(G1343gat));
  NOR2_X1   g662(.A1(new_n495), .A2(new_n364), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n695), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n865), .B(KEYINPUT117), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n497), .A2(KEYINPUT57), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n662), .A2(new_n840), .ZN(new_n868));
  AOI22_X1  g667(.A1(new_n868), .A2(new_n821), .B1(new_n620), .B2(new_n624), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n838), .A2(KEYINPUT118), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n871), .A2(new_n872), .A3(new_n841), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n552), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n551), .A2(new_n625), .A3(new_n704), .A4(new_n683), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n867), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n841), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n552), .B1(new_n877), .B2(new_n869), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n875), .ZN(new_n879));
  AOI21_X1  g678(.A(KEYINPUT57), .B1(new_n879), .B2(new_n497), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n662), .B(new_n866), .C1(new_n876), .C2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT120), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n883), .B1(new_n844), .B2(new_n297), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n843), .B1(new_n873), .B2(new_n552), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n884), .B1(new_n885), .B2(new_n867), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n886), .A2(new_n887), .A3(new_n662), .A4(new_n866), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n228), .B1(new_n882), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n297), .A2(new_n493), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n879), .A2(new_n864), .A3(new_n890), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n891), .A2(G141gat), .A3(new_n704), .ZN(new_n892));
  XNOR2_X1  g691(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT58), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n892), .B1(new_n881), .B2(G141gat), .ZN(new_n896));
  OAI22_X1  g695(.A1(new_n889), .A2(new_n894), .B1(new_n895), .B2(new_n896), .ZN(G1344gat));
  NAND3_X1  g696(.A1(new_n879), .A2(KEYINPUT57), .A3(new_n497), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n884), .A2(new_n898), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n866), .A2(new_n682), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n901), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n902));
  OAI21_X1  g701(.A(KEYINPUT59), .B1(new_n891), .B2(new_n683), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n229), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n886), .A2(new_n905), .A3(new_n900), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n902), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT121), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n902), .A2(new_n909), .A3(new_n904), .A4(new_n906), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(G1345gat));
  AND2_X1   g710(.A1(new_n886), .A2(new_n866), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n552), .A2(new_n226), .ZN(new_n913));
  XOR2_X1   g712(.A(new_n913), .B(KEYINPUT122), .Z(new_n914));
  NAND3_X1  g713(.A1(new_n845), .A2(new_n551), .A3(new_n890), .ZN(new_n915));
  AOI22_X1  g714(.A1(new_n912), .A2(new_n914), .B1(new_n915), .B2(new_n226), .ZN(G1346gat));
  NAND3_X1  g715(.A1(new_n886), .A2(new_n626), .A3(new_n866), .ZN(new_n917));
  OAI22_X1  g716(.A1(new_n917), .A2(KEYINPUT123), .B1(new_n224), .B2(new_n223), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n917), .A2(KEYINPUT123), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n890), .A2(new_n225), .ZN(new_n920));
  OAI22_X1  g719(.A1(new_n918), .A2(new_n919), .B1(new_n853), .B2(new_n920), .ZN(G1347gat));
  NAND4_X1  g720(.A1(new_n879), .A2(new_n495), .A3(new_n364), .A4(new_n501), .ZN(new_n922));
  INV_X1    g721(.A(G169gat), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n922), .A2(new_n923), .A3(new_n704), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n495), .B1(new_n842), .B2(new_n843), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT124), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n927), .B(new_n495), .C1(new_n842), .C2(new_n843), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n494), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n929), .A2(new_n501), .A3(new_n662), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n924), .B1(new_n930), .B2(new_n923), .ZN(G1348gat));
  OAI21_X1  g730(.A(G176gat), .B1(new_n922), .B2(new_n683), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n929), .A2(new_n501), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n683), .A2(G176gat), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(G1349gat));
  OAI21_X1  g734(.A(G183gat), .B1(new_n922), .B2(new_n552), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n551), .A2(new_n334), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n933), .B2(new_n937), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g738(.A(G190gat), .B1(new_n922), .B2(new_n625), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT61), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n626), .A2(new_n307), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n933), .B2(new_n942), .ZN(G1351gat));
  NAND4_X1  g742(.A1(new_n929), .A2(new_n213), .A3(new_n662), .A4(new_n890), .ZN(new_n944));
  INV_X1    g743(.A(new_n899), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n695), .A2(new_n495), .A3(new_n364), .ZN(new_n946));
  XOR2_X1   g745(.A(new_n946), .B(KEYINPUT125), .Z(new_n947));
  NOR3_X1   g746(.A1(new_n945), .A2(new_n704), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n944), .B1(new_n948), .B2(new_n213), .ZN(G1352gat));
  OR2_X1    g748(.A1(new_n945), .A2(new_n947), .ZN(new_n950));
  OAI21_X1  g749(.A(G204gat), .B1(new_n950), .B2(new_n683), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n926), .A2(new_n928), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n683), .A2(G204gat), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n952), .A2(new_n364), .A3(new_n890), .A4(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(KEYINPUT126), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n929), .A2(new_n956), .A3(new_n890), .A4(new_n953), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n955), .A2(KEYINPUT62), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(KEYINPUT62), .B1(new_n955), .B2(new_n957), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n951), .B1(new_n958), .B2(new_n959), .ZN(G1353gat));
  NAND4_X1  g759(.A1(new_n929), .A2(new_n216), .A3(new_n551), .A4(new_n890), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n552), .A2(new_n946), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n899), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n963), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n964));
  AOI21_X1  g763(.A(KEYINPUT63), .B1(new_n963), .B2(G211gat), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n965), .B2(KEYINPUT127), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT63), .ZN(new_n967));
  INV_X1    g766(.A(new_n962), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n968), .B1(new_n884), .B2(new_n898), .ZN(new_n969));
  OAI211_X1 g768(.A(KEYINPUT127), .B(new_n967), .C1(new_n969), .C2(new_n216), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n961), .B1(new_n966), .B2(new_n971), .ZN(G1354gat));
  OAI21_X1  g771(.A(G218gat), .B1(new_n950), .B2(new_n625), .ZN(new_n973));
  NAND4_X1  g772(.A1(new_n929), .A2(new_n217), .A3(new_n626), .A4(new_n890), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(G1355gat));
endmodule


