

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593;

  INV_X1 U323 ( .A(KEYINPUT72), .ZN(n379) );
  XNOR2_X1 U324 ( .A(n407), .B(KEYINPUT46), .ZN(n408) );
  INV_X1 U325 ( .A(n460), .ZN(n528) );
  XOR2_X1 U326 ( .A(n425), .B(n424), .Z(n291) );
  XOR2_X1 U327 ( .A(n375), .B(n441), .Z(n292) );
  XOR2_X1 U328 ( .A(G211GAT), .B(KEYINPUT21), .Z(n293) );
  XOR2_X1 U329 ( .A(KEYINPUT92), .B(n465), .Z(n294) );
  XNOR2_X1 U330 ( .A(KEYINPUT74), .B(G85GAT), .ZN(n357) );
  AND2_X1 U331 ( .A1(n415), .A2(n509), .ZN(n416) );
  XNOR2_X1 U332 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U333 ( .A(n382), .B(n381), .ZN(n386) );
  XNOR2_X1 U334 ( .A(n371), .B(n370), .ZN(n372) );
  NOR2_X1 U335 ( .A1(n418), .A2(n417), .ZN(n419) );
  NOR2_X1 U336 ( .A1(n471), .A2(n590), .ZN(n472) );
  NOR2_X1 U337 ( .A1(n554), .A2(n438), .ZN(n573) );
  XOR2_X1 U338 ( .A(KEYINPUT36), .B(n548), .Z(n590) );
  XNOR2_X1 U339 ( .A(n456), .B(KEYINPUT119), .ZN(n568) );
  XOR2_X1 U340 ( .A(n347), .B(n346), .Z(n554) );
  INV_X1 U341 ( .A(G43GAT), .ZN(n475) );
  XNOR2_X1 U342 ( .A(n474), .B(n473), .ZN(n507) );
  XNOR2_X1 U343 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n479) );
  XNOR2_X1 U344 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U345 ( .A(n480), .B(n479), .ZN(G1351GAT) );
  XNOR2_X1 U346 ( .A(n478), .B(n477), .ZN(G1330GAT) );
  XOR2_X1 U347 ( .A(G78GAT), .B(G71GAT), .Z(n296) );
  XNOR2_X1 U348 ( .A(G183GAT), .B(G127GAT), .ZN(n295) );
  XNOR2_X1 U349 ( .A(n296), .B(n295), .ZN(n310) );
  XOR2_X1 U350 ( .A(G57GAT), .B(KEYINPUT13), .Z(n387) );
  XOR2_X1 U351 ( .A(n387), .B(G155GAT), .Z(n299) );
  XNOR2_X1 U352 ( .A(G22GAT), .B(G15GAT), .ZN(n297) );
  XNOR2_X1 U353 ( .A(n297), .B(G1GAT), .ZN(n398) );
  XNOR2_X1 U354 ( .A(n398), .B(G211GAT), .ZN(n298) );
  XNOR2_X1 U355 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U356 ( .A(KEYINPUT77), .B(KEYINPUT12), .Z(n301) );
  NAND2_X1 U357 ( .A1(G231GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U358 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U359 ( .A(n303), .B(n302), .Z(n308) );
  XOR2_X1 U360 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n305) );
  XNOR2_X1 U361 ( .A(G8GAT), .B(G64GAT), .ZN(n304) );
  XNOR2_X1 U362 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U363 ( .A(n306), .B(KEYINPUT76), .ZN(n307) );
  XNOR2_X1 U364 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U365 ( .A(n310), .B(n309), .Z(n485) );
  INV_X1 U366 ( .A(n485), .ZN(n587) );
  XNOR2_X1 U367 ( .A(G197GAT), .B(KEYINPUT84), .ZN(n311) );
  XNOR2_X1 U368 ( .A(n293), .B(n311), .ZN(n425) );
  XOR2_X1 U369 ( .A(G155GAT), .B(KEYINPUT2), .Z(n313) );
  XNOR2_X1 U370 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n312) );
  XNOR2_X1 U371 ( .A(n313), .B(n312), .ZN(n337) );
  XNOR2_X1 U372 ( .A(n425), .B(n337), .ZN(n328) );
  XOR2_X1 U373 ( .A(G78GAT), .B(G148GAT), .Z(n315) );
  XNOR2_X1 U374 ( .A(KEYINPUT73), .B(G204GAT), .ZN(n314) );
  XNOR2_X1 U375 ( .A(n315), .B(n314), .ZN(n375) );
  XOR2_X1 U376 ( .A(G50GAT), .B(G162GAT), .Z(n369) );
  XOR2_X1 U377 ( .A(n375), .B(n369), .Z(n317) );
  XNOR2_X1 U378 ( .A(G218GAT), .B(G106GAT), .ZN(n316) );
  XNOR2_X1 U379 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U380 ( .A(KEYINPUT83), .B(KEYINPUT23), .Z(n319) );
  NAND2_X1 U381 ( .A1(G228GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U382 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U383 ( .A(n321), .B(n320), .Z(n326) );
  XOR2_X1 U384 ( .A(KEYINPUT24), .B(KEYINPUT85), .Z(n323) );
  XNOR2_X1 U385 ( .A(KEYINPUT82), .B(KEYINPUT22), .ZN(n322) );
  XNOR2_X1 U386 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U387 ( .A(G22GAT), .B(n324), .ZN(n325) );
  XNOR2_X1 U388 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U389 ( .A(n328), .B(n327), .ZN(n466) );
  XOR2_X1 U390 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n330) );
  XNOR2_X1 U391 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n329) );
  XNOR2_X1 U392 ( .A(n330), .B(n329), .ZN(n347) );
  XOR2_X1 U393 ( .A(KEYINPUT1), .B(G148GAT), .Z(n332) );
  XNOR2_X1 U394 ( .A(G120GAT), .B(G162GAT), .ZN(n331) );
  XNOR2_X1 U395 ( .A(n332), .B(n331), .ZN(n334) );
  XOR2_X1 U396 ( .A(G29GAT), .B(G85GAT), .Z(n333) );
  XNOR2_X1 U397 ( .A(n334), .B(n333), .ZN(n343) );
  XOR2_X1 U398 ( .A(G127GAT), .B(KEYINPUT0), .Z(n336) );
  XNOR2_X1 U399 ( .A(G113GAT), .B(G134GAT), .ZN(n335) );
  XNOR2_X1 U400 ( .A(n336), .B(n335), .ZN(n440) );
  XNOR2_X1 U401 ( .A(n440), .B(n337), .ZN(n341) );
  XOR2_X1 U402 ( .A(G57GAT), .B(KEYINPUT86), .Z(n339) );
  XNOR2_X1 U403 ( .A(KEYINPUT4), .B(KEYINPUT5), .ZN(n338) );
  XNOR2_X1 U404 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U405 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U406 ( .A(n343), .B(n342), .ZN(n345) );
  NAND2_X1 U407 ( .A1(G225GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U408 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U409 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n349) );
  XNOR2_X1 U410 ( .A(G43GAT), .B(G29GAT), .ZN(n348) );
  XNOR2_X1 U411 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U412 ( .A(KEYINPUT70), .B(n350), .Z(n402) );
  NAND2_X1 U413 ( .A1(G232GAT), .A2(G233GAT), .ZN(n356) );
  INV_X1 U414 ( .A(KEYINPUT11), .ZN(n351) );
  NAND2_X1 U415 ( .A1(n351), .A2(KEYINPUT64), .ZN(n354) );
  INV_X1 U416 ( .A(KEYINPUT64), .ZN(n352) );
  NAND2_X1 U417 ( .A1(n352), .A2(KEYINPUT11), .ZN(n353) );
  NAND2_X1 U418 ( .A1(n354), .A2(n353), .ZN(n355) );
  XOR2_X1 U419 ( .A(n356), .B(n355), .Z(n360) );
  INV_X1 U420 ( .A(n357), .ZN(n359) );
  XNOR2_X1 U421 ( .A(G99GAT), .B(G106GAT), .ZN(n358) );
  XNOR2_X1 U422 ( .A(n359), .B(n358), .ZN(n377) );
  XNOR2_X1 U423 ( .A(n360), .B(n377), .ZN(n368) );
  INV_X1 U424 ( .A(G218GAT), .ZN(n361) );
  NAND2_X1 U425 ( .A1(G92GAT), .A2(n361), .ZN(n364) );
  INV_X1 U426 ( .A(G92GAT), .ZN(n362) );
  NAND2_X1 U427 ( .A1(n362), .A2(G218GAT), .ZN(n363) );
  NAND2_X1 U428 ( .A1(n364), .A2(n363), .ZN(n366) );
  XNOR2_X1 U429 ( .A(G36GAT), .B(G190GAT), .ZN(n365) );
  XNOR2_X1 U430 ( .A(n366), .B(n365), .ZN(n428) );
  XNOR2_X1 U431 ( .A(G134GAT), .B(n428), .ZN(n367) );
  XNOR2_X1 U432 ( .A(n368), .B(n367), .ZN(n373) );
  XNOR2_X1 U433 ( .A(n369), .B(KEYINPUT9), .ZN(n371) );
  INV_X1 U434 ( .A(KEYINPUT10), .ZN(n370) );
  XNOR2_X1 U435 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U436 ( .A(n402), .B(n374), .ZN(n565) );
  XOR2_X1 U437 ( .A(G120GAT), .B(G71GAT), .Z(n441) );
  NAND2_X1 U438 ( .A1(G230GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U439 ( .A(n292), .B(n376), .ZN(n382) );
  BUF_X1 U440 ( .A(n377), .Z(n378) );
  XNOR2_X1 U441 ( .A(n378), .B(KEYINPUT32), .ZN(n380) );
  XOR2_X1 U442 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n384) );
  XNOR2_X1 U443 ( .A(G92GAT), .B(KEYINPUT71), .ZN(n383) );
  XNOR2_X1 U444 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U445 ( .A(n386), .B(n385), .Z(n389) );
  XOR2_X1 U446 ( .A(G176GAT), .B(G64GAT), .Z(n424) );
  XNOR2_X1 U447 ( .A(n424), .B(n387), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n389), .B(n388), .ZN(n580) );
  XNOR2_X1 U449 ( .A(KEYINPUT41), .B(n580), .ZN(n481) );
  XOR2_X1 U450 ( .A(KEYINPUT29), .B(KEYINPUT65), .Z(n391) );
  XNOR2_X1 U451 ( .A(KEYINPUT69), .B(KEYINPUT68), .ZN(n390) );
  XNOR2_X1 U452 ( .A(n391), .B(n390), .ZN(n406) );
  XOR2_X1 U453 ( .A(G141GAT), .B(G197GAT), .Z(n393) );
  XNOR2_X1 U454 ( .A(G36GAT), .B(G50GAT), .ZN(n392) );
  XNOR2_X1 U455 ( .A(n393), .B(n392), .ZN(n397) );
  XOR2_X1 U456 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n395) );
  XNOR2_X1 U457 ( .A(G113GAT), .B(KEYINPUT66), .ZN(n394) );
  XNOR2_X1 U458 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U459 ( .A(n397), .B(n396), .Z(n404) );
  XOR2_X1 U460 ( .A(G169GAT), .B(G8GAT), .Z(n432) );
  XOR2_X1 U461 ( .A(n432), .B(n398), .Z(n400) );
  NAND2_X1 U462 ( .A1(G229GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U463 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U464 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U465 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U466 ( .A(n406), .B(n405), .ZN(n575) );
  NAND2_X1 U467 ( .A1(n481), .A2(n575), .ZN(n407) );
  NAND2_X1 U468 ( .A1(n408), .A2(n485), .ZN(n409) );
  NOR2_X1 U469 ( .A1(n565), .A2(n409), .ZN(n410) );
  XOR2_X1 U470 ( .A(n410), .B(KEYINPUT47), .Z(n418) );
  INV_X1 U471 ( .A(KEYINPUT75), .ZN(n411) );
  XNOR2_X1 U472 ( .A(n411), .B(n565), .ZN(n548) );
  NOR2_X1 U473 ( .A1(n485), .A2(n590), .ZN(n412) );
  XNOR2_X1 U474 ( .A(KEYINPUT45), .B(n412), .ZN(n413) );
  NAND2_X1 U475 ( .A1(n413), .A2(n580), .ZN(n414) );
  XNOR2_X1 U476 ( .A(n414), .B(KEYINPUT109), .ZN(n415) );
  INV_X1 U477 ( .A(n575), .ZN(n509) );
  XNOR2_X1 U478 ( .A(n416), .B(KEYINPUT110), .ZN(n417) );
  XNOR2_X1 U479 ( .A(KEYINPUT48), .B(n419), .ZN(n536) );
  INV_X1 U480 ( .A(n536), .ZN(n436) );
  XNOR2_X1 U481 ( .A(KEYINPUT17), .B(KEYINPUT80), .ZN(n420) );
  XNOR2_X1 U482 ( .A(n420), .B(G183GAT), .ZN(n421) );
  XOR2_X1 U483 ( .A(n421), .B(KEYINPUT18), .Z(n423) );
  XNOR2_X1 U484 ( .A(KEYINPUT81), .B(KEYINPUT19), .ZN(n422) );
  XNOR2_X1 U485 ( .A(n423), .B(n422), .ZN(n454) );
  NAND2_X1 U486 ( .A1(G226GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U487 ( .A(n291), .B(n426), .ZN(n427) );
  XOR2_X1 U488 ( .A(n427), .B(KEYINPUT91), .Z(n430) );
  XNOR2_X1 U489 ( .A(n428), .B(KEYINPUT89), .ZN(n429) );
  XNOR2_X1 U490 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U491 ( .A(n431), .B(KEYINPUT90), .Z(n434) );
  XNOR2_X1 U492 ( .A(n432), .B(G204GAT), .ZN(n433) );
  XNOR2_X1 U493 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U494 ( .A(n454), .B(n435), .ZN(n460) );
  NAND2_X1 U495 ( .A1(n436), .A2(n528), .ZN(n437) );
  XNOR2_X1 U496 ( .A(n437), .B(KEYINPUT54), .ZN(n438) );
  NAND2_X1 U497 ( .A1(n466), .A2(n573), .ZN(n439) );
  XNOR2_X1 U498 ( .A(n439), .B(KEYINPUT55), .ZN(n455) );
  XOR2_X1 U499 ( .A(n441), .B(n440), .Z(n443) );
  XNOR2_X1 U500 ( .A(G99GAT), .B(G190GAT), .ZN(n442) );
  XNOR2_X1 U501 ( .A(n443), .B(n442), .ZN(n447) );
  XOR2_X1 U502 ( .A(KEYINPUT78), .B(G176GAT), .Z(n445) );
  NAND2_X1 U503 ( .A1(G227GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U504 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U505 ( .A(n447), .B(n446), .Z(n452) );
  XOR2_X1 U506 ( .A(KEYINPUT79), .B(KEYINPUT20), .Z(n449) );
  XNOR2_X1 U507 ( .A(G43GAT), .B(G15GAT), .ZN(n448) );
  XNOR2_X1 U508 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U509 ( .A(G169GAT), .B(n450), .ZN(n451) );
  XNOR2_X1 U510 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U511 ( .A(n454), .B(n453), .ZN(n537) );
  NAND2_X1 U512 ( .A1(n455), .A2(n537), .ZN(n456) );
  NAND2_X1 U513 ( .A1(n587), .A2(n568), .ZN(n458) );
  XNOR2_X1 U514 ( .A(G183GAT), .B(KEYINPUT120), .ZN(n457) );
  XNOR2_X1 U515 ( .A(n458), .B(n457), .ZN(G1350GAT) );
  NOR2_X1 U516 ( .A1(n466), .A2(n537), .ZN(n459) );
  XOR2_X1 U517 ( .A(KEYINPUT26), .B(n459), .Z(n572) );
  XNOR2_X1 U518 ( .A(KEYINPUT27), .B(n460), .ZN(n468) );
  NOR2_X1 U519 ( .A1(n572), .A2(n468), .ZN(n553) );
  NAND2_X1 U520 ( .A1(n528), .A2(n537), .ZN(n461) );
  NAND2_X1 U521 ( .A1(n466), .A2(n461), .ZN(n462) );
  XNOR2_X1 U522 ( .A(KEYINPUT25), .B(n462), .ZN(n463) );
  NOR2_X1 U523 ( .A1(n553), .A2(n463), .ZN(n464) );
  NOR2_X1 U524 ( .A1(n554), .A2(n464), .ZN(n465) );
  INV_X1 U525 ( .A(n537), .ZN(n469) );
  XNOR2_X1 U526 ( .A(n466), .B(KEYINPUT28), .ZN(n497) );
  NAND2_X1 U527 ( .A1(n554), .A2(n497), .ZN(n467) );
  NOR2_X1 U528 ( .A1(n468), .A2(n467), .ZN(n538) );
  NAND2_X1 U529 ( .A1(n469), .A2(n538), .ZN(n470) );
  NAND2_X1 U530 ( .A1(n294), .A2(n470), .ZN(n487) );
  NAND2_X1 U531 ( .A1(n485), .A2(n487), .ZN(n471) );
  XNOR2_X1 U532 ( .A(n472), .B(KEYINPUT37), .ZN(n523) );
  NAND2_X1 U533 ( .A1(n580), .A2(n575), .ZN(n489) );
  NOR2_X1 U534 ( .A1(n523), .A2(n489), .ZN(n474) );
  XNOR2_X1 U535 ( .A(KEYINPUT98), .B(KEYINPUT38), .ZN(n473) );
  NAND2_X1 U536 ( .A1(n507), .A2(n537), .ZN(n478) );
  XOR2_X1 U537 ( .A(KEYINPUT100), .B(KEYINPUT40), .Z(n476) );
  NAND2_X1 U538 ( .A1(n568), .A2(n548), .ZN(n480) );
  NAND2_X1 U539 ( .A1(n568), .A2(n481), .ZN(n484) );
  XOR2_X1 U540 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n482) );
  XNOR2_X1 U541 ( .A(n482), .B(G176GAT), .ZN(n483) );
  XNOR2_X1 U542 ( .A(n484), .B(n483), .ZN(G1349GAT) );
  NOR2_X1 U543 ( .A1(n485), .A2(n548), .ZN(n486) );
  XNOR2_X1 U544 ( .A(n486), .B(KEYINPUT16), .ZN(n488) );
  NAND2_X1 U545 ( .A1(n488), .A2(n487), .ZN(n511) );
  NOR2_X1 U546 ( .A1(n489), .A2(n511), .ZN(n498) );
  NAND2_X1 U547 ( .A1(n498), .A2(n554), .ZN(n490) );
  XNOR2_X1 U548 ( .A(n490), .B(KEYINPUT34), .ZN(n491) );
  XNOR2_X1 U549 ( .A(G1GAT), .B(n491), .ZN(G1324GAT) );
  XOR2_X1 U550 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n493) );
  NAND2_X1 U551 ( .A1(n498), .A2(n528), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U553 ( .A(G8GAT), .B(n494), .ZN(G1325GAT) );
  XOR2_X1 U554 ( .A(G15GAT), .B(KEYINPUT35), .Z(n496) );
  NAND2_X1 U555 ( .A1(n498), .A2(n537), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n496), .B(n495), .ZN(G1326GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n500) );
  INV_X1 U558 ( .A(n497), .ZN(n532) );
  NAND2_X1 U559 ( .A1(n498), .A2(n532), .ZN(n499) );
  XNOR2_X1 U560 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U561 ( .A(G22GAT), .B(n501), .ZN(G1327GAT) );
  XNOR2_X1 U562 ( .A(KEYINPUT99), .B(KEYINPUT39), .ZN(n505) );
  XOR2_X1 U563 ( .A(G29GAT), .B(KEYINPUT97), .Z(n503) );
  NAND2_X1 U564 ( .A1(n507), .A2(n554), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n505), .B(n504), .ZN(G1328GAT) );
  NAND2_X1 U567 ( .A1(n507), .A2(n528), .ZN(n506) );
  XNOR2_X1 U568 ( .A(n506), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U569 ( .A1(n507), .A2(n532), .ZN(n508) );
  XNOR2_X1 U570 ( .A(n508), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT102), .B(KEYINPUT42), .Z(n513) );
  NAND2_X1 U572 ( .A1(n481), .A2(n509), .ZN(n510) );
  XOR2_X1 U573 ( .A(KEYINPUT101), .B(n510), .Z(n524) );
  NOR2_X1 U574 ( .A1(n524), .A2(n511), .ZN(n519) );
  NAND2_X1 U575 ( .A1(n519), .A2(n554), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U577 ( .A(G57GAT), .B(n514), .Z(G1332GAT) );
  XOR2_X1 U578 ( .A(G64GAT), .B(KEYINPUT103), .Z(n516) );
  NAND2_X1 U579 ( .A1(n519), .A2(n528), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n516), .B(n515), .ZN(G1333GAT) );
  NAND2_X1 U581 ( .A1(n537), .A2(n519), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n517), .B(KEYINPUT104), .ZN(n518) );
  XNOR2_X1 U583 ( .A(G71GAT), .B(n518), .ZN(G1334GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT43), .B(KEYINPUT105), .Z(n521) );
  NAND2_X1 U585 ( .A1(n519), .A2(n532), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U587 ( .A(G78GAT), .B(n522), .Z(G1335GAT) );
  XOR2_X1 U588 ( .A(G85GAT), .B(KEYINPUT107), .Z(n527) );
  NOR2_X1 U589 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n525), .B(KEYINPUT106), .ZN(n533) );
  NAND2_X1 U591 ( .A1(n554), .A2(n533), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n527), .B(n526), .ZN(G1336GAT) );
  NAND2_X1 U593 ( .A1(n533), .A2(n528), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n529), .B(KEYINPUT108), .ZN(n530) );
  XNOR2_X1 U595 ( .A(G92GAT), .B(n530), .ZN(G1337GAT) );
  NAND2_X1 U596 ( .A1(n533), .A2(n537), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n531), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U598 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n534), .B(KEYINPUT44), .ZN(n535) );
  XNOR2_X1 U600 ( .A(G106GAT), .B(n535), .ZN(G1339GAT) );
  NAND2_X1 U601 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U602 ( .A1(n536), .A2(n539), .ZN(n549) );
  NAND2_X1 U603 ( .A1(n549), .A2(n575), .ZN(n540) );
  XNOR2_X1 U604 ( .A(G113GAT), .B(n540), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT112), .B(KEYINPUT49), .Z(n542) );
  NAND2_X1 U606 ( .A1(n549), .A2(n481), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(n544) );
  XOR2_X1 U608 ( .A(G120GAT), .B(KEYINPUT111), .Z(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(G1341GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT50), .B(KEYINPUT113), .Z(n546) );
  NAND2_X1 U611 ( .A1(n549), .A2(n587), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U613 ( .A(G127GAT), .B(n547), .ZN(G1342GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n551) );
  NAND2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U617 ( .A(G134GAT), .B(n552), .ZN(G1343GAT) );
  NAND2_X1 U618 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U619 ( .A1(n536), .A2(n555), .ZN(n564) );
  NAND2_X1 U620 ( .A1(n564), .A2(n575), .ZN(n556) );
  XNOR2_X1 U621 ( .A(G141GAT), .B(n556), .ZN(G1344GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT116), .B(KEYINPUT53), .Z(n558) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U625 ( .A(KEYINPUT115), .B(n559), .Z(n561) );
  NAND2_X1 U626 ( .A1(n564), .A2(n481), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1345GAT) );
  XOR2_X1 U628 ( .A(G155GAT), .B(KEYINPUT117), .Z(n563) );
  NAND2_X1 U629 ( .A1(n564), .A2(n587), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(G1346GAT) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(KEYINPUT118), .ZN(n567) );
  XNOR2_X1 U633 ( .A(G162GAT), .B(n567), .ZN(G1347GAT) );
  NAND2_X1 U634 ( .A1(n568), .A2(n575), .ZN(n569) );
  XNOR2_X1 U635 ( .A(G169GAT), .B(n569), .ZN(G1348GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT123), .B(KEYINPUT60), .Z(n571) );
  XNOR2_X1 U637 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n571), .B(n570), .ZN(n579) );
  XOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT59), .Z(n577) );
  INV_X1 U640 ( .A(n572), .ZN(n574) );
  NAND2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n589) );
  INV_X1 U642 ( .A(n589), .ZN(n586) );
  NAND2_X1 U643 ( .A1(n586), .A2(n575), .ZN(n576) );
  XNOR2_X1 U644 ( .A(n577), .B(n576), .ZN(n578) );
  XOR2_X1 U645 ( .A(n579), .B(n578), .Z(G1352GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n582) );
  OR2_X1 U647 ( .A1(n589), .A2(n580), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(n583) );
  XOR2_X1 U649 ( .A(n583), .B(KEYINPUT125), .Z(n585) );
  XNOR2_X1 U650 ( .A(G204GAT), .B(KEYINPUT124), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(G1353GAT) );
  NAND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n592) );
  XNOR2_X1 U655 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n591) );
  XNOR2_X1 U656 ( .A(n592), .B(n591), .ZN(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

