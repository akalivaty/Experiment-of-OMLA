

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576;

  XNOR2_X1 U323 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U324 ( .A(G169GAT), .B(G15GAT), .Z(n291) );
  XOR2_X1 U325 ( .A(G120GAT), .B(G71GAT), .Z(n423) );
  XNOR2_X1 U326 ( .A(n355), .B(n291), .ZN(n356) );
  AND2_X1 U327 ( .A1(n451), .A2(n407), .ZN(n409) );
  XOR2_X1 U328 ( .A(n539), .B(KEYINPUT28), .Z(n511) );
  XNOR2_X1 U329 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n446) );
  XNOR2_X1 U330 ( .A(n447), .B(n446), .ZN(G1330GAT) );
  XOR2_X1 U331 ( .A(KEYINPUT22), .B(KEYINPUT85), .Z(n293) );
  XNOR2_X1 U332 ( .A(KEYINPUT89), .B(KEYINPUT24), .ZN(n292) );
  XNOR2_X1 U333 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U334 ( .A(n294), .B(KEYINPUT88), .Z(n296) );
  XOR2_X1 U335 ( .A(G141GAT), .B(G22GAT), .Z(n432) );
  XNOR2_X1 U336 ( .A(G50GAT), .B(n432), .ZN(n295) );
  XNOR2_X1 U337 ( .A(n296), .B(n295), .ZN(n301) );
  XNOR2_X1 U338 ( .A(G106GAT), .B(G78GAT), .ZN(n297) );
  XNOR2_X1 U339 ( .A(n297), .B(G148GAT), .ZN(n411) );
  XOR2_X1 U340 ( .A(KEYINPUT23), .B(n411), .Z(n299) );
  NAND2_X1 U341 ( .A1(G228GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U342 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U343 ( .A(n301), .B(n300), .Z(n310) );
  XNOR2_X1 U344 ( .A(G211GAT), .B(G218GAT), .ZN(n302) );
  XNOR2_X1 U345 ( .A(n302), .B(KEYINPUT86), .ZN(n303) );
  XOR2_X1 U346 ( .A(n303), .B(KEYINPUT21), .Z(n305) );
  XNOR2_X1 U347 ( .A(G197GAT), .B(G204GAT), .ZN(n304) );
  XNOR2_X1 U348 ( .A(n305), .B(n304), .ZN(n321) );
  XOR2_X1 U349 ( .A(KEYINPUT2), .B(G162GAT), .Z(n307) );
  XNOR2_X1 U350 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n306) );
  XNOR2_X1 U351 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U352 ( .A(KEYINPUT87), .B(n308), .Z(n342) );
  XNOR2_X1 U353 ( .A(n321), .B(n342), .ZN(n309) );
  XNOR2_X1 U354 ( .A(n310), .B(n309), .ZN(n539) );
  XNOR2_X1 U355 ( .A(KEYINPUT27), .B(KEYINPUT96), .ZN(n325) );
  XOR2_X1 U356 ( .A(KEYINPUT18), .B(KEYINPUT84), .Z(n312) );
  XNOR2_X1 U357 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n311) );
  XNOR2_X1 U358 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U359 ( .A(KEYINPUT19), .B(n313), .Z(n359) );
  XNOR2_X1 U360 ( .A(G176GAT), .B(G92GAT), .ZN(n314) );
  XNOR2_X1 U361 ( .A(n314), .B(G64GAT), .ZN(n410) );
  XOR2_X1 U362 ( .A(n410), .B(G190GAT), .Z(n316) );
  XOR2_X1 U363 ( .A(G169GAT), .B(G8GAT), .Z(n429) );
  XNOR2_X1 U364 ( .A(G36GAT), .B(n429), .ZN(n315) );
  XNOR2_X1 U365 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U366 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n318) );
  NAND2_X1 U367 ( .A1(G226GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U368 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U369 ( .A(n320), .B(n319), .Z(n323) );
  XNOR2_X1 U370 ( .A(n321), .B(KEYINPUT93), .ZN(n322) );
  XNOR2_X1 U371 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U372 ( .A(n359), .B(n324), .ZN(n535) );
  INV_X1 U373 ( .A(n535), .ZN(n486) );
  XNOR2_X1 U374 ( .A(n325), .B(n486), .ZN(n365) );
  XOR2_X1 U375 ( .A(KEYINPUT6), .B(KEYINPUT90), .Z(n327) );
  XNOR2_X1 U376 ( .A(G120GAT), .B(G148GAT), .ZN(n326) );
  XNOR2_X1 U377 ( .A(n327), .B(n326), .ZN(n331) );
  XOR2_X1 U378 ( .A(KEYINPUT5), .B(G57GAT), .Z(n329) );
  XNOR2_X1 U379 ( .A(KEYINPUT1), .B(KEYINPUT4), .ZN(n328) );
  XNOR2_X1 U380 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U381 ( .A(n331), .B(n330), .Z(n336) );
  XOR2_X1 U382 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n333) );
  NAND2_X1 U383 ( .A1(G225GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U384 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U385 ( .A(G1GAT), .B(n334), .ZN(n335) );
  XNOR2_X1 U386 ( .A(n336), .B(n335), .ZN(n341) );
  XOR2_X1 U387 ( .A(G85GAT), .B(G134GAT), .Z(n339) );
  XNOR2_X1 U388 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n337) );
  XNOR2_X1 U389 ( .A(n337), .B(G127GAT), .ZN(n355) );
  XNOR2_X1 U390 ( .A(G141GAT), .B(n355), .ZN(n338) );
  XNOR2_X1 U391 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U392 ( .A(n341), .B(n340), .Z(n344) );
  XNOR2_X1 U393 ( .A(G29GAT), .B(n342), .ZN(n343) );
  XNOR2_X1 U394 ( .A(n344), .B(n343), .ZN(n538) );
  NAND2_X1 U395 ( .A1(n365), .A2(n538), .ZN(n345) );
  XOR2_X1 U396 ( .A(KEYINPUT97), .B(n345), .Z(n507) );
  NOR2_X1 U397 ( .A1(n511), .A2(n507), .ZN(n346) );
  XNOR2_X1 U398 ( .A(KEYINPUT98), .B(n346), .ZN(n360) );
  XOR2_X1 U399 ( .A(KEYINPUT20), .B(KEYINPUT65), .Z(n348) );
  XNOR2_X1 U400 ( .A(G176GAT), .B(KEYINPUT83), .ZN(n347) );
  XOR2_X1 U401 ( .A(n348), .B(n347), .Z(n352) );
  XOR2_X1 U402 ( .A(G99GAT), .B(n423), .Z(n350) );
  XOR2_X1 U403 ( .A(G190GAT), .B(G134GAT), .Z(n398) );
  XNOR2_X1 U404 ( .A(G43GAT), .B(n398), .ZN(n349) );
  XNOR2_X1 U405 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U406 ( .A(n352), .B(n351), .ZN(n354) );
  NAND2_X1 U407 ( .A1(G227GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U408 ( .A(n354), .B(n353), .ZN(n357) );
  XNOR2_X1 U409 ( .A(n359), .B(n358), .ZN(n542) );
  AND2_X1 U410 ( .A1(n360), .A2(n542), .ZN(n371) );
  NOR2_X1 U411 ( .A1(n542), .A2(n535), .ZN(n361) );
  XNOR2_X1 U412 ( .A(KEYINPUT99), .B(n361), .ZN(n362) );
  NAND2_X1 U413 ( .A1(n362), .A2(n539), .ZN(n363) );
  XNOR2_X1 U414 ( .A(n363), .B(KEYINPUT25), .ZN(n367) );
  INV_X1 U415 ( .A(n542), .ZN(n508) );
  NOR2_X1 U416 ( .A1(n508), .A2(n539), .ZN(n364) );
  XNOR2_X1 U417 ( .A(KEYINPUT26), .B(n364), .ZN(n558) );
  AND2_X1 U418 ( .A1(n365), .A2(n558), .ZN(n366) );
  NOR2_X1 U419 ( .A1(n367), .A2(n366), .ZN(n368) );
  NOR2_X1 U420 ( .A1(n538), .A2(n368), .ZN(n369) );
  XNOR2_X1 U421 ( .A(n369), .B(KEYINPUT100), .ZN(n370) );
  NOR2_X1 U422 ( .A1(n371), .A2(n370), .ZN(n372) );
  XNOR2_X1 U423 ( .A(n372), .B(KEYINPUT101), .ZN(n451) );
  XOR2_X1 U424 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n374) );
  XNOR2_X1 U425 ( .A(KEYINPUT15), .B(KEYINPUT79), .ZN(n373) );
  XNOR2_X1 U426 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U427 ( .A(G57GAT), .B(KEYINPUT13), .Z(n413) );
  XOR2_X1 U428 ( .A(n413), .B(G211GAT), .Z(n376) );
  XOR2_X1 U429 ( .A(G15GAT), .B(G1GAT), .Z(n428) );
  XNOR2_X1 U430 ( .A(G22GAT), .B(n428), .ZN(n375) );
  XNOR2_X1 U431 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U432 ( .A(n378), .B(n377), .Z(n380) );
  NAND2_X1 U433 ( .A1(G231GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U434 ( .A(n380), .B(n379), .ZN(n388) );
  XOR2_X1 U435 ( .A(G78GAT), .B(G155GAT), .Z(n382) );
  XNOR2_X1 U436 ( .A(G127GAT), .B(G71GAT), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n382), .B(n381), .ZN(n386) );
  XOR2_X1 U438 ( .A(KEYINPUT80), .B(G64GAT), .Z(n384) );
  XNOR2_X1 U439 ( .A(G8GAT), .B(G183GAT), .ZN(n383) );
  XNOR2_X1 U440 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U441 ( .A(n386), .B(n385), .Z(n387) );
  XNOR2_X1 U442 ( .A(n388), .B(n387), .ZN(n550) );
  XNOR2_X1 U443 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n389) );
  XNOR2_X1 U444 ( .A(n389), .B(G29GAT), .ZN(n390) );
  XOR2_X1 U445 ( .A(n390), .B(KEYINPUT8), .Z(n392) );
  XNOR2_X1 U446 ( .A(G43GAT), .B(G50GAT), .ZN(n391) );
  XNOR2_X1 U447 ( .A(n392), .B(n391), .ZN(n443) );
  XOR2_X1 U448 ( .A(KEYINPUT67), .B(KEYINPUT10), .Z(n394) );
  XNOR2_X1 U449 ( .A(G162GAT), .B(G106GAT), .ZN(n393) );
  XNOR2_X1 U450 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U451 ( .A(n443), .B(n395), .ZN(n406) );
  XOR2_X1 U452 ( .A(KEYINPUT11), .B(KEYINPUT78), .Z(n397) );
  XNOR2_X1 U453 ( .A(KEYINPUT77), .B(KEYINPUT9), .ZN(n396) );
  XNOR2_X1 U454 ( .A(n397), .B(n396), .ZN(n402) );
  XOR2_X1 U455 ( .A(G99GAT), .B(G85GAT), .Z(n412) );
  XOR2_X1 U456 ( .A(n412), .B(G92GAT), .Z(n400) );
  XNOR2_X1 U457 ( .A(n398), .B(G218GAT), .ZN(n399) );
  XNOR2_X1 U458 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U459 ( .A(n402), .B(n401), .Z(n404) );
  NAND2_X1 U460 ( .A1(G232GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U461 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n532) );
  XNOR2_X1 U463 ( .A(KEYINPUT36), .B(n532), .ZN(n573) );
  NOR2_X1 U464 ( .A1(n550), .A2(n573), .ZN(n407) );
  XNOR2_X1 U465 ( .A(KEYINPUT37), .B(KEYINPUT106), .ZN(n408) );
  XNOR2_X1 U466 ( .A(n409), .B(n408), .ZN(n484) );
  XNOR2_X1 U467 ( .A(n411), .B(n410), .ZN(n427) );
  XOR2_X1 U468 ( .A(n413), .B(n412), .Z(n415) );
  NAND2_X1 U469 ( .A1(G230GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U470 ( .A(n415), .B(n414), .ZN(n419) );
  XOR2_X1 U471 ( .A(KEYINPUT32), .B(KEYINPUT73), .Z(n417) );
  XNOR2_X1 U472 ( .A(KEYINPUT76), .B(KEYINPUT75), .ZN(n416) );
  XNOR2_X1 U473 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U474 ( .A(n419), .B(n418), .Z(n425) );
  XOR2_X1 U475 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n421) );
  XNOR2_X1 U476 ( .A(G204GAT), .B(KEYINPUT74), .ZN(n420) );
  XNOR2_X1 U477 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U478 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U479 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U480 ( .A(n427), .B(n426), .ZN(n565) );
  XOR2_X1 U481 ( .A(n429), .B(n428), .Z(n431) );
  NAND2_X1 U482 ( .A1(G229GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U483 ( .A(n431), .B(n430), .ZN(n433) );
  XOR2_X1 U484 ( .A(n433), .B(n432), .Z(n441) );
  XOR2_X1 U485 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n435) );
  XNOR2_X1 U486 ( .A(G197GAT), .B(G113GAT), .ZN(n434) );
  XNOR2_X1 U487 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U488 ( .A(KEYINPUT69), .B(KEYINPUT71), .Z(n437) );
  XNOR2_X1 U489 ( .A(KEYINPUT70), .B(KEYINPUT29), .ZN(n436) );
  XNOR2_X1 U490 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U491 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U492 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U493 ( .A(n443), .B(n442), .ZN(n560) );
  XOR2_X1 U494 ( .A(n560), .B(KEYINPUT72), .Z(n543) );
  NAND2_X1 U495 ( .A1(n565), .A2(n543), .ZN(n453) );
  NOR2_X1 U496 ( .A1(n484), .A2(n453), .ZN(n444) );
  XOR2_X1 U497 ( .A(KEYINPUT38), .B(n444), .Z(n445) );
  XNOR2_X1 U498 ( .A(KEYINPUT107), .B(n445), .ZN(n469) );
  NAND2_X1 U499 ( .A1(n469), .A2(n508), .ZN(n447) );
  XOR2_X1 U500 ( .A(KEYINPUT34), .B(KEYINPUT103), .Z(n456) );
  NAND2_X1 U501 ( .A1(n550), .A2(n532), .ZN(n450) );
  XNOR2_X1 U502 ( .A(KEYINPUT16), .B(KEYINPUT82), .ZN(n448) );
  XNOR2_X1 U503 ( .A(n448), .B(KEYINPUT81), .ZN(n449) );
  XNOR2_X1 U504 ( .A(n450), .B(n449), .ZN(n452) );
  NAND2_X1 U505 ( .A1(n452), .A2(n451), .ZN(n473) );
  NOR2_X1 U506 ( .A1(n453), .A2(n473), .ZN(n454) );
  XNOR2_X1 U507 ( .A(KEYINPUT102), .B(n454), .ZN(n462) );
  NAND2_X1 U508 ( .A1(n538), .A2(n462), .ZN(n455) );
  XNOR2_X1 U509 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U510 ( .A(G1GAT), .B(n457), .ZN(G1324GAT) );
  NAND2_X1 U511 ( .A1(n462), .A2(n486), .ZN(n458) );
  XNOR2_X1 U512 ( .A(n458), .B(KEYINPUT104), .ZN(n459) );
  XNOR2_X1 U513 ( .A(G8GAT), .B(n459), .ZN(G1325GAT) );
  XOR2_X1 U514 ( .A(G15GAT), .B(KEYINPUT35), .Z(n461) );
  NAND2_X1 U515 ( .A1(n508), .A2(n462), .ZN(n460) );
  XNOR2_X1 U516 ( .A(n461), .B(n460), .ZN(G1326GAT) );
  NAND2_X1 U517 ( .A1(n462), .A2(n511), .ZN(n463) );
  XNOR2_X1 U518 ( .A(n463), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U519 ( .A(KEYINPUT108), .B(KEYINPUT39), .Z(n465) );
  XNOR2_X1 U520 ( .A(G29GAT), .B(KEYINPUT105), .ZN(n464) );
  XNOR2_X1 U521 ( .A(n465), .B(n464), .ZN(n467) );
  NAND2_X1 U522 ( .A1(n469), .A2(n538), .ZN(n466) );
  XOR2_X1 U523 ( .A(n467), .B(n466), .Z(G1328GAT) );
  NAND2_X1 U524 ( .A1(n486), .A2(n469), .ZN(n468) );
  XNOR2_X1 U525 ( .A(G36GAT), .B(n468), .ZN(G1329GAT) );
  XOR2_X1 U526 ( .A(G50GAT), .B(KEYINPUT109), .Z(n471) );
  NAND2_X1 U527 ( .A1(n511), .A2(n469), .ZN(n470) );
  XNOR2_X1 U528 ( .A(n471), .B(n470), .ZN(G1331GAT) );
  XNOR2_X1 U529 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n475) );
  XOR2_X1 U530 ( .A(KEYINPUT41), .B(KEYINPUT64), .Z(n472) );
  XNOR2_X1 U531 ( .A(n565), .B(n472), .ZN(n527) );
  INV_X1 U532 ( .A(n527), .ZN(n545) );
  NAND2_X1 U533 ( .A1(n545), .A2(n560), .ZN(n483) );
  NOR2_X1 U534 ( .A1(n473), .A2(n483), .ZN(n479) );
  NAND2_X1 U535 ( .A1(n538), .A2(n479), .ZN(n474) );
  XNOR2_X1 U536 ( .A(n475), .B(n474), .ZN(G1332GAT) );
  NAND2_X1 U537 ( .A1(n479), .A2(n486), .ZN(n476) );
  XNOR2_X1 U538 ( .A(n476), .B(KEYINPUT110), .ZN(n477) );
  XNOR2_X1 U539 ( .A(G64GAT), .B(n477), .ZN(G1333GAT) );
  NAND2_X1 U540 ( .A1(n479), .A2(n508), .ZN(n478) );
  XNOR2_X1 U541 ( .A(n478), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U542 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n481) );
  NAND2_X1 U543 ( .A1(n479), .A2(n511), .ZN(n480) );
  XNOR2_X1 U544 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U545 ( .A(G78GAT), .B(n482), .Z(G1335GAT) );
  NOR2_X1 U546 ( .A1(n484), .A2(n483), .ZN(n491) );
  NAND2_X1 U547 ( .A1(n538), .A2(n491), .ZN(n485) );
  XNOR2_X1 U548 ( .A(G85GAT), .B(n485), .ZN(G1336GAT) );
  NAND2_X1 U549 ( .A1(n491), .A2(n486), .ZN(n487) );
  XNOR2_X1 U550 ( .A(n487), .B(KEYINPUT112), .ZN(n488) );
  XNOR2_X1 U551 ( .A(G92GAT), .B(n488), .ZN(G1337GAT) );
  XOR2_X1 U552 ( .A(G99GAT), .B(KEYINPUT113), .Z(n490) );
  NAND2_X1 U553 ( .A1(n491), .A2(n508), .ZN(n489) );
  XNOR2_X1 U554 ( .A(n490), .B(n489), .ZN(G1338GAT) );
  NAND2_X1 U555 ( .A1(n491), .A2(n511), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n492), .B(KEYINPUT44), .ZN(n493) );
  XNOR2_X1 U557 ( .A(G106GAT), .B(n493), .ZN(G1339GAT) );
  XOR2_X1 U558 ( .A(G113GAT), .B(KEYINPUT117), .Z(n513) );
  NOR2_X1 U559 ( .A1(n560), .A2(n527), .ZN(n495) );
  XNOR2_X1 U560 ( .A(KEYINPUT46), .B(KEYINPUT114), .ZN(n494) );
  XNOR2_X1 U561 ( .A(n495), .B(n494), .ZN(n496) );
  NOR2_X1 U562 ( .A1(n496), .A2(n550), .ZN(n497) );
  NAND2_X1 U563 ( .A1(n532), .A2(n497), .ZN(n498) );
  XNOR2_X1 U564 ( .A(n498), .B(KEYINPUT47), .ZN(n505) );
  XNOR2_X1 U565 ( .A(KEYINPUT115), .B(KEYINPUT45), .ZN(n499) );
  XNOR2_X1 U566 ( .A(n499), .B(KEYINPUT66), .ZN(n501) );
  INV_X1 U567 ( .A(n550), .ZN(n570) );
  NOR2_X1 U568 ( .A1(n573), .A2(n570), .ZN(n500) );
  XOR2_X1 U569 ( .A(n501), .B(n500), .Z(n502) );
  NAND2_X1 U570 ( .A1(n565), .A2(n502), .ZN(n503) );
  NOR2_X1 U571 ( .A1(n543), .A2(n503), .ZN(n504) );
  NOR2_X1 U572 ( .A1(n505), .A2(n504), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n506), .B(KEYINPUT48), .ZN(n534) );
  NOR2_X1 U574 ( .A1(n534), .A2(n507), .ZN(n522) );
  NAND2_X1 U575 ( .A1(n508), .A2(n522), .ZN(n509) );
  XNOR2_X1 U576 ( .A(KEYINPUT116), .B(n509), .ZN(n510) );
  NOR2_X1 U577 ( .A1(n511), .A2(n510), .ZN(n518) );
  NAND2_X1 U578 ( .A1(n518), .A2(n543), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(G1340GAT) );
  XOR2_X1 U580 ( .A(G120GAT), .B(KEYINPUT49), .Z(n515) );
  NAND2_X1 U581 ( .A1(n518), .A2(n545), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n515), .B(n514), .ZN(G1341GAT) );
  NAND2_X1 U583 ( .A1(n550), .A2(n518), .ZN(n516) );
  XNOR2_X1 U584 ( .A(n516), .B(KEYINPUT50), .ZN(n517) );
  XNOR2_X1 U585 ( .A(G127GAT), .B(n517), .ZN(G1342GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n520) );
  INV_X1 U587 ( .A(n532), .ZN(n553) );
  NAND2_X1 U588 ( .A1(n518), .A2(n553), .ZN(n519) );
  XNOR2_X1 U589 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U590 ( .A(G134GAT), .B(n521), .ZN(G1343GAT) );
  NAND2_X1 U591 ( .A1(n522), .A2(n558), .ZN(n531) );
  NOR2_X1 U592 ( .A1(n560), .A2(n531), .ZN(n524) );
  XNOR2_X1 U593 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n523) );
  XNOR2_X1 U594 ( .A(n524), .B(n523), .ZN(G1344GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT120), .B(KEYINPUT52), .Z(n526) );
  XNOR2_X1 U596 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n525) );
  XNOR2_X1 U597 ( .A(n526), .B(n525), .ZN(n529) );
  NOR2_X1 U598 ( .A1(n527), .A2(n531), .ZN(n528) );
  XOR2_X1 U599 ( .A(n529), .B(n528), .Z(G1345GAT) );
  NOR2_X1 U600 ( .A1(n570), .A2(n531), .ZN(n530) );
  XOR2_X1 U601 ( .A(G155GAT), .B(n530), .Z(G1346GAT) );
  NOR2_X1 U602 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U603 ( .A(G162GAT), .B(n533), .Z(G1347GAT) );
  NOR2_X1 U604 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U605 ( .A(KEYINPUT54), .B(n536), .Z(n537) );
  NOR2_X1 U606 ( .A1(n538), .A2(n537), .ZN(n559) );
  NAND2_X1 U607 ( .A1(n539), .A2(n559), .ZN(n540) );
  XOR2_X1 U608 ( .A(KEYINPUT55), .B(n540), .Z(n541) );
  NOR2_X1 U609 ( .A1(n542), .A2(n541), .ZN(n554) );
  NAND2_X1 U610 ( .A1(n543), .A2(n554), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n544), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U612 ( .A(G176GAT), .B(KEYINPUT56), .Z(n547) );
  NAND2_X1 U613 ( .A1(n554), .A2(n545), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(n549) );
  XOR2_X1 U615 ( .A(KEYINPUT121), .B(KEYINPUT57), .Z(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(G1349GAT) );
  NAND2_X1 U617 ( .A1(n550), .A2(n554), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n551), .B(KEYINPUT122), .ZN(n552) );
  XNOR2_X1 U619 ( .A(G183GAT), .B(n552), .ZN(G1350GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n556) );
  NAND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G190GAT), .B(n557), .ZN(G1351GAT) );
  NAND2_X1 U624 ( .A1(n559), .A2(n558), .ZN(n572) );
  NOR2_X1 U625 ( .A1(n560), .A2(n572), .ZN(n564) );
  XNOR2_X1 U626 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(KEYINPUT59), .ZN(n562) );
  XNOR2_X1 U628 ( .A(KEYINPUT60), .B(n562), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(G1352GAT) );
  NOR2_X1 U630 ( .A1(n572), .A2(n565), .ZN(n569) );
  XOR2_X1 U631 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n567) );
  XNOR2_X1 U632 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1353GAT) );
  NOR2_X1 U635 ( .A1(n570), .A2(n572), .ZN(n571) );
  XOR2_X1 U636 ( .A(G211GAT), .B(n571), .Z(G1354GAT) );
  NOR2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n575) );
  XNOR2_X1 U638 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U640 ( .A(G218GAT), .B(n576), .ZN(G1355GAT) );
endmodule

