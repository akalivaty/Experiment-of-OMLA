//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n548, new_n549, new_n550, new_n551, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n582, new_n583, new_n584, new_n585, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1168, new_n1169, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT65), .Z(G319));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  AND2_X1   g034(.A1(new_n459), .A2(G125), .ZN(new_n460));
  AND2_X1   g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(G2105), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n464));
  XOR2_X1   g039(.A(new_n464), .B(KEYINPUT67), .Z(new_n465));
  AND3_X1   g040(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(KEYINPUT3), .B1(KEYINPUT66), .B2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G137), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n462), .A2(new_n465), .A3(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(G160));
  OAI21_X1  g047(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(G112), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n473), .B1(new_n474), .B2(G2105), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n468), .A2(new_n463), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n475), .B1(new_n476), .B2(G124), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n469), .A2(G136), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  INV_X1    g055(.A(KEYINPUT4), .ZN(new_n481));
  NAND4_X1  g056(.A1(new_n459), .A2(new_n481), .A3(G138), .A4(new_n463), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT68), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n482), .B(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n481), .B1(new_n469), .B2(G138), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G2105), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n490), .B1(new_n476), .B2(G126), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G164));
  INV_X1    g068(.A(KEYINPUT72), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT5), .B1(new_n494), .B2(G543), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n494), .B2(G543), .ZN(new_n496));
  XNOR2_X1  g071(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n497));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT74), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT74), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT73), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n503), .A2(KEYINPUT73), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n500), .B(G543), .C1(new_n502), .C2(new_n504), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n496), .B1(new_n499), .B2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT69), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT69), .A2(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n506), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n513), .B1(new_n514), .B2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(KEYINPUT71), .A3(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT70), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n519), .B1(new_n510), .B2(KEYINPUT6), .ZN(new_n520));
  NOR4_X1   g095(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT70), .A4(new_n516), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n512), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n511), .A2(new_n523), .ZN(G166));
  INV_X1    g099(.A(KEYINPUT76), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g101(.A(KEYINPUT76), .B(new_n518), .C1(new_n520), .C2(new_n521), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n526), .A2(G543), .A3(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G51), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT75), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n532), .B(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XOR2_X1   g110(.A(new_n535), .B(KEYINPUT7), .Z(new_n536));
  OR2_X1    g111(.A1(KEYINPUT69), .A2(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(KEYINPUT69), .A2(G651), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n537), .A2(KEYINPUT6), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(KEYINPUT70), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n510), .A2(new_n519), .A3(KEYINPUT6), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n540), .A2(new_n541), .B1(new_n515), .B2(new_n517), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n542), .A2(new_n506), .ZN(new_n543));
  XNOR2_X1  g118(.A(KEYINPUT77), .B(G89), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n536), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n534), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n531), .A2(new_n546), .ZN(G168));
  AOI22_X1  g122(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n510), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n549), .B1(G90), .B2(new_n543), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n529), .A2(G52), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  AOI22_X1  g128(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  OR2_X1    g129(.A1(new_n554), .A2(new_n510), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n526), .A2(G43), .A3(G543), .A4(new_n527), .ZN(new_n556));
  INV_X1    g131(.A(G81), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n542), .A2(new_n506), .ZN(new_n558));
  OAI211_X1 g133(.A(new_n555), .B(new_n556), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  INV_X1    g140(.A(KEYINPUT78), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n542), .A2(new_n506), .A3(G91), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(new_n506), .B2(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n567), .B1(new_n570), .B2(new_n514), .ZN(new_n571));
  AND2_X1   g146(.A1(G53), .A2(G543), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n526), .A2(new_n527), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(KEYINPUT9), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n526), .A2(new_n575), .A3(new_n527), .A4(new_n572), .ZN(new_n576));
  AOI211_X1 g151(.A(new_n566), .B(new_n571), .C1(new_n574), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n574), .A2(new_n576), .ZN(new_n578));
  INV_X1    g153(.A(new_n571), .ZN(new_n579));
  AOI21_X1  g154(.A(KEYINPUT78), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n577), .A2(new_n580), .ZN(G299));
  OAI21_X1  g156(.A(KEYINPUT79), .B1(new_n531), .B2(new_n546), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT79), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n530), .A2(new_n534), .A3(new_n583), .A4(new_n545), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G286));
  OR2_X1    g161(.A1(new_n511), .A2(new_n523), .ZN(G303));
  NAND2_X1  g162(.A1(new_n543), .A2(G87), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n589));
  INV_X1    g164(.A(G49), .ZN(new_n590));
  OAI211_X1 g165(.A(new_n588), .B(new_n589), .C1(new_n590), .C2(new_n528), .ZN(G288));
  NAND2_X1  g166(.A1(new_n506), .A2(G61), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n592), .A2(KEYINPUT80), .B1(G73), .B2(G543), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(KEYINPUT80), .B2(new_n592), .ZN(new_n594));
  INV_X1    g169(.A(new_n510), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n506), .A2(G86), .ZN(new_n597));
  AND2_X1   g172(.A1(G48), .A2(G543), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n542), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n596), .A2(new_n599), .ZN(G305));
  NAND2_X1  g175(.A1(new_n529), .A2(G47), .ZN(new_n601));
  AND2_X1   g176(.A1(new_n506), .A2(G60), .ZN(new_n602));
  AND2_X1   g177(.A1(G72), .A2(G543), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n595), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n543), .A2(G85), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n601), .A2(new_n604), .A3(new_n605), .ZN(G290));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NOR2_X1   g182(.A1(G301), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT81), .ZN(new_n609));
  INV_X1    g184(.A(G66), .ZN(new_n610));
  AOI211_X1 g185(.A(new_n610), .B(new_n496), .C1(new_n499), .C2(new_n505), .ZN(new_n611));
  AND2_X1   g186(.A1(G79), .A2(G543), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n609), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n612), .B1(new_n506), .B2(G66), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(KEYINPUT81), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n613), .A2(new_n615), .A3(G651), .ZN(new_n616));
  NAND4_X1  g191(.A1(new_n526), .A2(G54), .A3(G543), .A4(new_n527), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT10), .ZN(new_n618));
  INV_X1    g193(.A(G92), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n558), .B2(new_n619), .ZN(new_n620));
  NAND4_X1  g195(.A1(new_n542), .A2(new_n506), .A3(KEYINPUT10), .A4(G92), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n616), .A2(new_n617), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT82), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n608), .B1(new_n624), .B2(new_n607), .ZN(G284));
  AOI21_X1  g200(.A(new_n608), .B1(new_n624), .B2(new_n607), .ZN(G321));
  NOR2_X1   g201(.A1(G299), .A2(G868), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n627), .B1(G868), .B2(new_n585), .ZN(G297));
  XOR2_X1   g203(.A(G297), .B(KEYINPUT83), .Z(G280));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n624), .B1(new_n630), .B2(G860), .ZN(G148));
  NAND2_X1  g206(.A1(new_n624), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G868), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n633), .A2(KEYINPUT84), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(KEYINPUT84), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n634), .B(new_n635), .C1(G868), .C2(new_n560), .ZN(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g212(.A1(new_n469), .A2(G135), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n476), .A2(G123), .ZN(new_n639));
  OR2_X1    g214(.A1(G99), .A2(G2105), .ZN(new_n640));
  OAI211_X1 g215(.A(new_n640), .B(G2104), .C1(G111), .C2(new_n463), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n638), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2096), .Z(new_n643));
  NAND3_X1  g218(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT12), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT13), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2100), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT85), .ZN(G156));
  INV_X1    g224(.A(KEYINPUT14), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n650), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n653), .B2(new_n652), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n655), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  AND3_X1   g238(.A1(new_n662), .A2(G14), .A3(new_n663), .ZN(G401));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n665), .B1(new_n668), .B2(KEYINPUT18), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT86), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2100), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT18), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n668), .A2(KEYINPUT17), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n666), .A2(new_n667), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(G2096), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n671), .B(new_n676), .ZN(G227));
  XOR2_X1   g252(.A(G1971), .B(G1976), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1956), .B(G2474), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1961), .B(G1966), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT20), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n680), .A2(new_n681), .ZN(new_n685));
  NOR3_X1   g260(.A1(new_n679), .A2(new_n682), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(new_n679), .B2(new_n685), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1991), .B(G1996), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1981), .B(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(G229));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G6), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n596), .A2(new_n599), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(new_n695), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT89), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT32), .B(G1981), .Z(new_n701));
  OR2_X1    g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n695), .A2(G23), .ZN(new_n704));
  INV_X1    g279(.A(G288), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(new_n705), .B2(new_n695), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT33), .B(G1976), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT90), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n706), .A2(new_n709), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n695), .A2(G22), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G166), .B2(new_n695), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n713), .A2(G1971), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n713), .A2(G1971), .ZN(new_n715));
  NOR4_X1   g290(.A1(new_n710), .A2(new_n711), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n702), .A2(new_n703), .A3(new_n716), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n717), .A2(KEYINPUT34), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(KEYINPUT34), .ZN(new_n719));
  NOR2_X1   g294(.A1(G16), .A2(G24), .ZN(new_n720));
  INV_X1    g295(.A(G290), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(G16), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n722), .A2(G1986), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(G1986), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n469), .A2(G131), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT87), .Z(new_n726));
  OAI21_X1  g301(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n727));
  INV_X1    g302(.A(G107), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(G2105), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n476), .B2(G119), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  MUX2_X1   g306(.A(G25), .B(new_n731), .S(G29), .Z(new_n732));
  XOR2_X1   g307(.A(KEYINPUT35), .B(G1991), .Z(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT88), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n732), .B(new_n734), .ZN(new_n735));
  NOR3_X1   g310(.A1(new_n723), .A2(new_n724), .A3(new_n735), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n718), .A2(new_n719), .A3(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT36), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n695), .A2(G20), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT97), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT23), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n578), .A2(new_n579), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(new_n566), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n578), .A2(KEYINPUT78), .A3(new_n579), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n742), .B1(new_n746), .B2(new_n695), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G1956), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n695), .A2(G19), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n560), .B2(new_n695), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(G1341), .Z(new_n751));
  INV_X1    g326(.A(G29), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G32), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n469), .A2(G141), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT94), .ZN(new_n755));
  AND3_X1   g330(.A1(new_n463), .A2(G105), .A3(G2104), .ZN(new_n756));
  NAND3_X1  g331(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT26), .ZN(new_n758));
  AOI211_X1 g333(.A(new_n756), .B(new_n758), .C1(new_n476), .C2(G129), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n753), .B1(new_n761), .B2(new_n752), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT27), .B(G1996), .Z(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT95), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n762), .B(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G2090), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n752), .A2(G35), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G162), .B2(new_n752), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT29), .Z(new_n769));
  OAI21_X1  g344(.A(new_n765), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n766), .B2(new_n769), .ZN(new_n771));
  NOR2_X1   g346(.A1(G164), .A2(new_n752), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G27), .B2(new_n752), .ZN(new_n773));
  INV_X1    g348(.A(G2078), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n752), .A2(G26), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT28), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n469), .A2(G140), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n476), .A2(G128), .ZN(new_n780));
  OAI21_X1  g355(.A(KEYINPUT92), .B1(G104), .B2(G2105), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  NOR3_X1   g357(.A1(KEYINPUT92), .A2(G104), .A3(G2105), .ZN(new_n783));
  OAI221_X1 g358(.A(G2104), .B1(G116), .B2(new_n463), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n779), .A2(new_n780), .A3(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n778), .B1(new_n786), .B2(new_n752), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G2067), .ZN(new_n788));
  NOR3_X1   g363(.A1(new_n775), .A2(new_n776), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n469), .A2(G139), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT93), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n459), .A2(G127), .ZN(new_n792));
  NAND2_X1  g367(.A1(G115), .A2(G2104), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n463), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT25), .ZN(new_n795));
  NAND2_X1  g370(.A1(G103), .A2(G2104), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n795), .B1(new_n796), .B2(G2105), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n463), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n794), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n791), .A2(new_n799), .ZN(new_n800));
  MUX2_X1   g375(.A(G33), .B(new_n800), .S(G29), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G2072), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n642), .A2(new_n752), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT96), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT30), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n805), .A2(G28), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n752), .B1(new_n805), .B2(G28), .ZN(new_n807));
  AND2_X1   g382(.A1(KEYINPUT31), .A2(G11), .ZN(new_n808));
  NOR2_X1   g383(.A1(KEYINPUT31), .A2(G11), .ZN(new_n809));
  OAI22_X1  g384(.A1(new_n806), .A2(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(G34), .ZN(new_n811));
  AOI21_X1  g386(.A(G29), .B1(new_n811), .B2(KEYINPUT24), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(KEYINPUT24), .B2(new_n811), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n471), .B2(new_n752), .ZN(new_n814));
  INV_X1    g389(.A(G2084), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NOR4_X1   g391(.A1(new_n802), .A2(new_n804), .A3(new_n810), .A4(new_n816), .ZN(new_n817));
  AND4_X1   g392(.A1(new_n751), .A2(new_n771), .A3(new_n789), .A4(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n695), .A2(G4), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n624), .B2(new_n695), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT91), .B(G1348), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n820), .B(new_n821), .Z(new_n822));
  NOR2_X1   g397(.A1(G168), .A2(new_n695), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n695), .B2(G21), .ZN(new_n824));
  INV_X1    g399(.A(G1966), .ZN(new_n825));
  INV_X1    g400(.A(G1961), .ZN(new_n826));
  NOR2_X1   g401(.A1(G171), .A2(new_n695), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(G5), .B2(new_n695), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n824), .A2(new_n825), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(new_n826), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n824), .A2(new_n825), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n818), .A2(new_n822), .A3(new_n829), .A4(new_n832), .ZN(new_n833));
  NOR3_X1   g408(.A1(new_n739), .A2(new_n748), .A3(new_n833), .ZN(G311));
  OR3_X1    g409(.A1(new_n739), .A2(new_n748), .A3(new_n833), .ZN(G150));
  NAND2_X1  g410(.A1(new_n624), .A2(G559), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT38), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n838));
  INV_X1    g413(.A(G93), .ZN(new_n839));
  OAI22_X1  g414(.A1(new_n838), .A2(new_n510), .B1(new_n558), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(new_n529), .B2(G55), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n559), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n837), .B(new_n842), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n843), .A2(KEYINPUT39), .ZN(new_n844));
  INV_X1    g419(.A(G860), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(KEYINPUT39), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n841), .A2(new_n845), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT37), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(G145));
  XNOR2_X1  g425(.A(new_n731), .B(KEYINPUT100), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n645), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n476), .A2(G130), .ZN(new_n853));
  OR2_X1    g428(.A1(G106), .A2(G2105), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n854), .B(G2104), .C1(G118), .C2(new_n463), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(G142), .B2(new_n469), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n852), .B(new_n857), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n858), .A2(KEYINPUT102), .ZN(new_n859));
  INV_X1    g434(.A(new_n491), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n482), .B(KEYINPUT68), .ZN(new_n861));
  OAI21_X1  g436(.A(KEYINPUT98), .B1(new_n861), .B2(new_n485), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT98), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n484), .A2(new_n486), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n860), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n786), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n761), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n791), .A2(KEYINPUT99), .A3(new_n799), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT99), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n800), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n867), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(new_n868), .B2(new_n867), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n859), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n479), .B(new_n642), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n471), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n875), .B1(new_n859), .B2(new_n872), .ZN(new_n876));
  AOI21_X1  g451(.A(G37), .B1(new_n873), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT101), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n872), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n872), .A2(new_n878), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(new_n880), .A3(new_n858), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n881), .B(new_n875), .C1(new_n880), .C2(new_n858), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g459(.A(new_n623), .B1(new_n577), .B2(new_n580), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT104), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n746), .A2(KEYINPUT104), .A3(new_n623), .ZN(new_n888));
  INV_X1    g463(.A(new_n623), .ZN(new_n889));
  AOI21_X1  g464(.A(KEYINPUT103), .B1(G299), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT103), .ZN(new_n891));
  NOR4_X1   g466(.A1(new_n577), .A2(new_n580), .A3(new_n891), .A4(new_n623), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n887), .B(new_n888), .C1(new_n890), .C2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT41), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n744), .A2(new_n745), .A3(new_n889), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n891), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n744), .A2(KEYINPUT103), .A3(new_n745), .A4(new_n889), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI22_X1  g473(.A1(new_n893), .A2(new_n894), .B1(new_n898), .B2(new_n885), .ZN(new_n899));
  INV_X1    g474(.A(new_n842), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n632), .B(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n896), .A2(new_n897), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n885), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  OR3_X1    g480(.A1(new_n902), .A2(new_n905), .A3(KEYINPUT42), .ZN(new_n906));
  XNOR2_X1  g481(.A(G166), .B(KEYINPUT105), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(new_n721), .ZN(new_n908));
  XNOR2_X1  g483(.A(G305), .B(new_n705), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n908), .A2(new_n909), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT42), .B1(new_n902), .B2(new_n905), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n906), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n913), .B1(new_n906), .B2(new_n914), .ZN(new_n916));
  OAI21_X1  g491(.A(G868), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n917), .B1(G868), .B2(new_n841), .ZN(G295));
  OAI21_X1  g493(.A(new_n917), .B1(G868), .B2(new_n841), .ZN(G331));
  INV_X1    g494(.A(G37), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT106), .ZN(new_n921));
  AOI21_X1  g496(.A(G301), .B1(new_n582), .B2(new_n584), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(G171), .A2(G168), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n923), .A2(new_n900), .A3(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n842), .B1(new_n922), .B2(new_n924), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n904), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n921), .B(new_n929), .C1(new_n899), .C2(new_n928), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(new_n911), .B2(new_n912), .ZN(new_n932));
  OR2_X1    g507(.A1(new_n908), .A2(new_n909), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n933), .A2(new_n910), .A3(KEYINPUT107), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n930), .A2(new_n935), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n926), .A2(new_n927), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n885), .B(KEYINPUT104), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT41), .B1(new_n938), .B2(new_n903), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n903), .A2(KEYINPUT41), .A3(new_n885), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n921), .B1(new_n941), .B2(new_n929), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n920), .B1(new_n936), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT108), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI211_X1 g520(.A(KEYINPUT108), .B(new_n920), .C1(new_n936), .C2(new_n942), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n941), .A2(new_n913), .A3(new_n929), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n941), .A2(KEYINPUT109), .A3(new_n913), .A4(new_n929), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n945), .A2(KEYINPUT43), .A3(new_n946), .A4(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT110), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n929), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n928), .A2(KEYINPUT110), .A3(new_n904), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n904), .A2(new_n894), .B1(new_n938), .B2(new_n898), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n955), .B(new_n956), .C1(new_n928), .C2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(G37), .B1(new_n958), .B2(new_n935), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n951), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n952), .A2(new_n953), .A3(new_n962), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n951), .A2(new_n959), .A3(KEYINPUT43), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n945), .A2(new_n946), .A3(new_n951), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n964), .B1(new_n965), .B2(new_n961), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n963), .B1(new_n966), .B2(new_n953), .ZN(G397));
  INV_X1    g542(.A(KEYINPUT120), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n862), .A2(new_n864), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n491), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT113), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT50), .ZN(new_n972));
  INV_X1    g547(.A(G1384), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n970), .A2(new_n971), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(KEYINPUT111), .B(G40), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n471), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n492), .A2(new_n973), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n977), .B1(new_n978), .B2(KEYINPUT50), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n974), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n970), .A2(new_n973), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT113), .B1(new_n981), .B2(KEYINPUT50), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n821), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n865), .A2(G1384), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n976), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n985), .A2(G2067), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n968), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n986), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n974), .A2(new_n979), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n971), .B1(new_n984), .B2(new_n972), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI211_X1 g566(.A(KEYINPUT120), .B(new_n988), .C1(new_n991), .C2(new_n821), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n987), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n623), .B1(new_n993), .B2(KEYINPUT60), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT60), .ZN(new_n995));
  AOI211_X1 g570(.A(new_n995), .B(new_n889), .C1(new_n987), .C2(new_n992), .ZN(new_n996));
  OAI22_X1  g571(.A1(new_n994), .A2(new_n996), .B1(KEYINPUT60), .B2(new_n993), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n984), .A2(KEYINPUT45), .ZN(new_n998));
  AOI21_X1  g573(.A(G1384), .B1(new_n487), .B2(new_n491), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n976), .B1(new_n999), .B2(KEYINPUT45), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g576(.A(KEYINPUT56), .B(G2072), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n998), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n977), .B1(new_n999), .B2(new_n972), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1004), .B1(new_n984), .B2(new_n972), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1003), .B1(new_n1006), .B2(G1956), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT119), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n743), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT57), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n1009), .B(KEYINPUT57), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1000), .B1(new_n984), .B2(KEYINPUT45), .ZN(new_n1014));
  INV_X1    g589(.A(G1956), .ZN(new_n1015));
  AOI22_X1  g590(.A1(new_n1014), .A2(new_n1002), .B1(new_n1005), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n1012), .A2(new_n1017), .A3(KEYINPUT61), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT61), .B1(new_n1012), .B2(new_n1017), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT122), .ZN(new_n1021));
  INV_X1    g596(.A(G1996), .ZN(new_n1022));
  XOR2_X1   g597(.A(KEYINPUT58), .B(G1341), .Z(new_n1023));
  AOI22_X1  g598(.A1(new_n1014), .A2(new_n1022), .B1(new_n985), .B2(new_n1023), .ZN(new_n1024));
  OR3_X1    g599(.A1(new_n1024), .A2(KEYINPUT121), .A3(new_n559), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT121), .B1(new_n1024), .B2(new_n559), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(new_n1026), .A3(KEYINPUT59), .ZN(new_n1027));
  OR2_X1    g602(.A1(new_n1026), .A2(KEYINPUT59), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1020), .A2(new_n1021), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1012), .A2(new_n1017), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT61), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1012), .A2(new_n1017), .A3(KEYINPUT61), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1032), .A2(new_n1027), .A3(new_n1028), .A4(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT122), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n997), .A2(new_n1029), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n993), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n623), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n1037), .A2(new_n1038), .B1(new_n1011), .B2(new_n1007), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G8), .ZN(new_n1041));
  NOR2_X1   g616(.A1(G168), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n982), .A2(new_n815), .A3(new_n974), .A4(new_n979), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n984), .A2(KEYINPUT45), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT45), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n976), .B1(new_n978), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n825), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1043), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1044), .A2(new_n1048), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(G8), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1042), .A2(KEYINPUT51), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT124), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1041), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT124), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1052), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1053), .A2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1043), .B1(new_n1054), .B2(KEYINPUT123), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1050), .A2(KEYINPUT123), .A3(G8), .ZN(new_n1060));
  OAI21_X1  g635(.A(KEYINPUT51), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1049), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n1063));
  XOR2_X1   g638(.A(KEYINPUT112), .B(G1971), .Z(new_n1064));
  NOR2_X1   g639(.A1(new_n1014), .A2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1005), .A2(G2090), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1063), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  OAI221_X1 g642(.A(KEYINPUT118), .B1(new_n1005), .B2(G2090), .C1(new_n1064), .C2(new_n1014), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(new_n1068), .A3(G8), .ZN(new_n1069));
  NOR2_X1   g644(.A1(G166), .A2(new_n1041), .ZN(new_n1070));
  XOR2_X1   g645(.A(KEYINPUT114), .B(KEYINPUT55), .Z(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT55), .ZN(new_n1073));
  OAI22_X1  g648(.A1(G166), .A2(new_n1041), .B1(KEYINPUT114), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1069), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n985), .A2(G8), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n697), .B(G1981), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1078), .B1(new_n1079), .B2(KEYINPUT49), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT115), .ZN(new_n1081));
  OR2_X1    g656(.A1(G305), .A2(G1981), .ZN(new_n1082));
  NAND2_X1  g657(.A1(G305), .A2(G1981), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT49), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1081), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AOI211_X1 g661(.A(KEYINPUT115), .B(KEYINPUT49), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1080), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n989), .A2(new_n990), .A3(G2090), .ZN(new_n1089));
  OAI211_X1 g664(.A(G8), .B(new_n1075), .C1(new_n1089), .C2(new_n1065), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n705), .A2(G1976), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n985), .A2(new_n1091), .A3(G8), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n705), .A2(G1976), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1092), .A2(KEYINPUT52), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1094), .B1(KEYINPUT52), .B2(new_n1092), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1077), .A2(new_n1088), .A3(new_n1090), .A4(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(G301), .B(KEYINPUT54), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1014), .A2(new_n774), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT53), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1100), .B1(G1961), .B2(new_n991), .ZN(new_n1101));
  NAND2_X1  g676(.A1(G160), .A2(G40), .ZN(new_n1102));
  OAI211_X1 g677(.A(KEYINPUT53), .B(new_n774), .C1(new_n1102), .C2(KEYINPUT125), .ZN(new_n1103));
  AOI211_X1 g678(.A(new_n1103), .B(new_n1045), .C1(KEYINPUT125), .C2(new_n1102), .ZN(new_n1104));
  AOI211_X1 g679(.A(new_n1097), .B(new_n1101), .C1(new_n998), .C2(new_n1104), .ZN(new_n1105));
  NOR4_X1   g680(.A1(new_n1045), .A2(new_n1099), .A3(new_n1047), .A4(G2078), .ZN(new_n1106));
  OR2_X1    g681(.A1(new_n1101), .A2(new_n1106), .ZN(new_n1107));
  AND2_X1   g682(.A1(new_n1107), .A2(new_n1097), .ZN(new_n1108));
  NOR4_X1   g683(.A1(new_n1062), .A2(new_n1096), .A3(new_n1105), .A4(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1040), .A2(new_n1109), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT62), .B1(new_n1111), .B2(new_n1049), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1062), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT126), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1107), .A2(G171), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1096), .A2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1112), .A2(new_n1114), .A3(new_n1115), .A4(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1117), .B1(new_n1062), .B2(new_n1113), .ZN(new_n1119));
  AOI211_X1 g694(.A(KEYINPUT62), .B(new_n1049), .C1(new_n1058), .C2(new_n1061), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT126), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1082), .ZN(new_n1122));
  NOR2_X1   g697(.A1(G288), .A2(G1976), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1122), .B1(new_n1088), .B2(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1078), .B(KEYINPUT116), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1088), .A2(new_n1095), .ZN(new_n1126));
  OAI22_X1  g701(.A1(new_n1124), .A2(new_n1125), .B1(new_n1126), .B2(new_n1090), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT117), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT117), .ZN(new_n1129));
  OAI221_X1 g704(.A(new_n1129), .B1(new_n1126), .B2(new_n1090), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT63), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1054), .A2(new_n585), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1131), .B1(new_n1096), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1126), .ZN(new_n1134));
  OAI21_X1  g709(.A(G8), .B1(new_n1089), .B2(new_n1065), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n1076), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1132), .A2(new_n1131), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1134), .A2(new_n1090), .A3(new_n1136), .A4(new_n1137), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n1128), .A2(new_n1130), .B1(new_n1133), .B2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1110), .A2(new_n1118), .A3(new_n1121), .A4(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n760), .B(new_n1022), .ZN(new_n1141));
  INV_X1    g716(.A(G2067), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n785), .B(new_n1142), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n731), .B(new_n733), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1144), .B(new_n1145), .C1(G1986), .C2(G290), .ZN(new_n1146));
  AND2_X1   g721(.A1(G290), .A2(G1986), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1045), .B(new_n976), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1140), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1045), .A2(new_n976), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1150), .B1(new_n761), .B2(new_n1143), .ZN(new_n1151));
  OR3_X1    g726(.A1(new_n1150), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1152));
  OAI21_X1  g727(.A(KEYINPUT46), .B1(new_n1150), .B2(G1996), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1151), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  XOR2_X1   g729(.A(new_n1154), .B(KEYINPUT47), .Z(new_n1155));
  NAND4_X1  g730(.A1(new_n1144), .A2(new_n726), .A3(new_n730), .A4(new_n733), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n786), .A2(new_n1142), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1150), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1150), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1150), .A2(G1986), .A3(G290), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1159), .B1(KEYINPUT48), .B2(new_n1160), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n1160), .A2(KEYINPUT48), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1158), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1155), .A2(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1164), .B(KEYINPUT127), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1149), .A2(new_n1165), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g741(.A(G319), .ZN(new_n1168));
  NOR4_X1   g742(.A1(G229), .A2(new_n1168), .A3(G401), .A4(G227), .ZN(new_n1169));
  AND2_X1   g743(.A1(new_n883), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g744(.A1(new_n1170), .A2(new_n962), .A3(new_n952), .ZN(G225));
  INV_X1    g745(.A(G225), .ZN(G308));
endmodule


