//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 0 0 0 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n538, new_n540, new_n541, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n554, new_n555,
    new_n556, new_n557, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n601, new_n603, new_n604, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1155, new_n1156, new_n1157, new_n1159, new_n1160, new_n1161,
    new_n1162;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  XNOR2_X1  g013(.A(KEYINPUT66), .B(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  XNOR2_X1  g015(.A(KEYINPUT67), .B(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G125), .ZN(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n464));
  NAND2_X1  g039(.A1(G101), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n466), .B1(new_n460), .B2(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n464), .B1(new_n467), .B2(G2105), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n470), .A2(new_n472), .A3(G137), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(new_n465), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(KEYINPUT68), .A3(new_n459), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n463), .B1(new_n468), .B2(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n470), .A2(new_n472), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(new_n459), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n477), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  NOR2_X1   g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(new_n459), .B2(G112), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n479), .B(new_n481), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  NAND3_X1  g060(.A1(new_n459), .A2(G102), .A3(G2104), .ZN(new_n486));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(new_n469), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(new_n460), .B2(G126), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n486), .B1(new_n489), .B2(new_n459), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n470), .A2(new_n472), .A3(G138), .A4(new_n459), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n460), .A2(KEYINPUT4), .A3(G138), .A4(new_n459), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n490), .A2(new_n495), .ZN(G164));
  AND2_X1   g071(.A1(KEYINPUT6), .A2(G651), .ZN(new_n497));
  NOR2_X1   g072(.A1(KEYINPUT6), .A2(G651), .ZN(new_n498));
  OR2_X1    g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G50), .ZN(new_n501));
  INV_X1    g076(.A(G88), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G543), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n504), .B(new_n506), .C1(new_n497), .C2(new_n498), .ZN(new_n507));
  OAI22_X1  g082(.A1(new_n500), .A2(new_n501), .B1(new_n502), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n504), .A2(new_n506), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G62), .ZN(new_n511));
  NAND2_X1  g086(.A1(G75), .A2(G543), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n508), .A2(new_n513), .ZN(G166));
  NAND3_X1  g089(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n515));
  XOR2_X1   g090(.A(new_n515), .B(KEYINPUT69), .Z(new_n516));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT7), .ZN(new_n518));
  INV_X1    g093(.A(G89), .ZN(new_n519));
  XOR2_X1   g094(.A(KEYINPUT70), .B(G51), .Z(new_n520));
  OAI221_X1 g095(.A(new_n518), .B1(new_n519), .B2(new_n507), .C1(new_n500), .C2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n516), .A2(new_n521), .ZN(G168));
  AOI22_X1  g097(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n523), .A2(new_n509), .ZN(new_n524));
  INV_X1    g099(.A(G52), .ZN(new_n525));
  INV_X1    g100(.A(G90), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n500), .A2(new_n525), .B1(new_n526), .B2(new_n507), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n524), .A2(new_n527), .ZN(G171));
  OAI211_X1 g103(.A(G43), .B(G543), .C1(new_n497), .C2(new_n498), .ZN(new_n529));
  INV_X1    g104(.A(G81), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n507), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(G68), .A2(G543), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n504), .A2(new_n506), .ZN(new_n533));
  INV_X1    g108(.A(G56), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n531), .B1(G651), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G860), .ZN(G153));
  AND3_X1   g112(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G36), .ZN(G176));
  NAND2_X1  g114(.A1(G1), .A2(G3), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT8), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n538), .A2(new_n541), .ZN(G188));
  OAI211_X1 g117(.A(G53), .B(G543), .C1(new_n497), .C2(new_n498), .ZN(new_n543));
  XOR2_X1   g118(.A(new_n543), .B(KEYINPUT9), .Z(new_n544));
  INV_X1    g119(.A(new_n507), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G91), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n510), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n547), .B2(new_n509), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(G299));
  INV_X1    g125(.A(G171), .ZN(G301));
  OR2_X1    g126(.A1(new_n516), .A2(new_n521), .ZN(G286));
  OR2_X1    g127(.A1(new_n508), .A2(new_n513), .ZN(G303));
  AND2_X1   g128(.A1(new_n499), .A2(G543), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G49), .ZN(new_n555));
  OAI21_X1  g130(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n545), .A2(G87), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(G288));
  INV_X1    g133(.A(G61), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT71), .B1(new_n533), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(G73), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT71), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n504), .A2(new_n506), .A3(new_n562), .A4(G61), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G651), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n554), .A2(G48), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n545), .A2(G86), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(G305));
  AOI22_X1  g143(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n569), .A2(new_n509), .ZN(new_n570));
  INV_X1    g145(.A(G47), .ZN(new_n571));
  INV_X1    g146(.A(G85), .ZN(new_n572));
  OAI22_X1  g147(.A1(new_n500), .A2(new_n571), .B1(new_n572), .B2(new_n507), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G290));
  NAND2_X1  g150(.A1(G301), .A2(G868), .ZN(new_n576));
  INV_X1    g151(.A(G92), .ZN(new_n577));
  OR3_X1    g152(.A1(new_n507), .A2(KEYINPUT72), .A3(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(KEYINPUT72), .B1(new_n507), .B2(new_n577), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT10), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(G79), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G66), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n533), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n554), .A2(G54), .B1(new_n585), .B2(G651), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n578), .A2(KEYINPUT10), .A3(new_n579), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n582), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT73), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n588), .B(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT74), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n588), .B(KEYINPUT73), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(KEYINPUT74), .ZN(new_n594));
  AND2_X1   g169(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n576), .B1(new_n595), .B2(G868), .ZN(G321));
  XOR2_X1   g171(.A(G321), .B(KEYINPUT75), .Z(G284));
  NAND2_X1  g172(.A1(G286), .A2(G868), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n598), .B1(G868), .B2(new_n549), .ZN(G297));
  XNOR2_X1  g174(.A(G297), .B(KEYINPUT76), .ZN(G280));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n595), .B1(new_n601), .B2(G860), .ZN(G148));
  NAND3_X1  g177(.A1(new_n592), .A2(new_n594), .A3(new_n601), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G868), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G868), .B2(new_n536), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT77), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g182(.A1(new_n478), .A2(G123), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n480), .A2(G135), .ZN(new_n609));
  NOR2_X1   g184(.A1(G99), .A2(G2105), .ZN(new_n610));
  OAI21_X1  g185(.A(G2104), .B1(new_n459), .B2(G111), .ZN(new_n611));
  OAI211_X1 g186(.A(new_n608), .B(new_n609), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT78), .Z(new_n613));
  OR2_X1    g188(.A1(new_n613), .A2(G2096), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n459), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT13), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(G2100), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n613), .A2(G2096), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n614), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT79), .Z(G156));
  XOR2_X1   g196(.A(KEYINPUT15), .B(G2435), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2438), .ZN(new_n623));
  XOR2_X1   g198(.A(G2427), .B(G2430), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT81), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n623), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(KEYINPUT14), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2451), .B(G2454), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2443), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2446), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n627), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(KEYINPUT82), .B(KEYINPUT83), .Z(new_n632));
  XNOR2_X1  g207(.A(G1341), .B(G1348), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n631), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n635), .B(new_n636), .Z(new_n637));
  AND2_X1   g212(.A1(new_n637), .A2(G14), .ZN(G401));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2067), .B(G2678), .Z(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(new_n643), .A3(KEYINPUT17), .ZN(new_n644));
  INV_X1    g219(.A(KEYINPUT18), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2072), .B(G2078), .Z(new_n647));
  AOI21_X1  g222(.A(new_n647), .B1(new_n642), .B2(KEYINPUT18), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n646), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2096), .B(G2100), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT84), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n649), .B(new_n651), .ZN(G227));
  XNOR2_X1  g227(.A(G1971), .B(G1976), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT19), .ZN(new_n654));
  XOR2_X1   g229(.A(G1956), .B(G2474), .Z(new_n655));
  XOR2_X1   g230(.A(G1961), .B(G1966), .Z(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n655), .A2(new_n656), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT20), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n654), .A2(new_n657), .A3(new_n659), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n662), .B(new_n663), .C1(new_n661), .C2(new_n660), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT21), .B(G1986), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G1991), .B(G1996), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT22), .B(G1981), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(G229));
  INV_X1    g247(.A(G16), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(G4), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n674), .B1(new_n595), .B2(new_n673), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n675), .A2(KEYINPUT89), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(KEYINPUT89), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G1348), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT25), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n460), .A2(G127), .ZN(new_n682));
  NAND2_X1  g257(.A1(G115), .A2(G2104), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n459), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  AOI211_X1 g259(.A(new_n681), .B(new_n684), .C1(G139), .C2(new_n480), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT91), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G29), .ZN(new_n688));
  OAI21_X1  g263(.A(KEYINPUT90), .B1(G29), .B2(G33), .ZN(new_n689));
  NOR2_X1   g264(.A1(G29), .A2(G33), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT90), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g267(.A1(new_n688), .A2(G2072), .A3(new_n689), .A4(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT93), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI22_X1  g270(.A1(new_n687), .A2(G29), .B1(new_n691), .B2(new_n690), .ZN(new_n696));
  NAND4_X1  g271(.A1(new_n696), .A2(KEYINPUT93), .A3(G2072), .A4(new_n689), .ZN(new_n697));
  INV_X1    g272(.A(G2090), .ZN(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G35), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G162), .B2(new_n699), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT29), .Z(new_n702));
  AOI22_X1  g277(.A1(new_n695), .A2(new_n697), .B1(new_n698), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n699), .A2(G26), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n478), .A2(G128), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n480), .A2(G140), .ZN(new_n706));
  OR2_X1    g281(.A1(G104), .A2(G2105), .ZN(new_n707));
  OAI211_X1 g282(.A(new_n707), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n705), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n704), .B1(new_n710), .B2(new_n699), .ZN(new_n711));
  MUX2_X1   g286(.A(new_n704), .B(new_n711), .S(KEYINPUT28), .Z(new_n712));
  INV_X1    g287(.A(G2067), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n673), .A2(G21), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G168), .B2(new_n673), .ZN(new_n716));
  INV_X1    g291(.A(G1966), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  OR2_X1    g293(.A1(G29), .A2(G32), .ZN(new_n719));
  AOI22_X1  g294(.A1(G129), .A2(new_n478), .B1(new_n480), .B2(G141), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n459), .A2(G105), .A3(G2104), .ZN(new_n721));
  NAND3_X1  g296(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT26), .Z(new_n723));
  NAND3_X1  g298(.A1(new_n720), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n719), .B1(new_n724), .B2(new_n699), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT27), .B(G1996), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT30), .B(G28), .Z(new_n727));
  OAI22_X1  g302(.A1(new_n725), .A2(new_n726), .B1(G29), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(G16), .A2(G19), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n536), .B2(G16), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n728), .B1(G1341), .B2(new_n730), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n703), .A2(new_n714), .A3(new_n718), .A4(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(G2072), .B1(new_n696), .B2(new_n689), .ZN(new_n733));
  NAND2_X1  g308(.A1(G160), .A2(G29), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT92), .B(KEYINPUT24), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(G34), .Z(new_n736));
  OAI21_X1  g311(.A(new_n734), .B1(G29), .B2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G2084), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n733), .A2(new_n739), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n730), .A2(G1341), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n702), .A2(new_n698), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT31), .B(G11), .Z(new_n743));
  NAND2_X1  g318(.A1(new_n699), .A2(G27), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G164), .B2(new_n699), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G2078), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n673), .A2(KEYINPUT23), .A3(G20), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT23), .ZN(new_n748));
  INV_X1    g323(.A(G20), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(G16), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n747), .B(new_n750), .C1(new_n549), .C2(new_n673), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G1956), .ZN(new_n752));
  NOR4_X1   g327(.A1(new_n742), .A2(new_n743), .A3(new_n746), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n725), .A2(new_n726), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n740), .A2(new_n741), .A3(new_n753), .A4(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n732), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n673), .A2(G23), .ZN(new_n757));
  INV_X1    g332(.A(G288), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n758), .B2(new_n673), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT33), .B(G1976), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT86), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n759), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n673), .A2(G22), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G166), .B2(new_n673), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(G1971), .Z(new_n765));
  AND2_X1   g340(.A1(new_n673), .A2(G6), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G305), .B2(G16), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT32), .B(G1981), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n762), .A2(new_n765), .A3(new_n769), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT34), .Z(new_n771));
  NOR2_X1   g346(.A1(G16), .A2(G24), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n574), .B(KEYINPUT85), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(G16), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G1986), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n699), .A2(G25), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n478), .A2(G119), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n480), .A2(G131), .ZN(new_n778));
  OR2_X1    g353(.A1(G95), .A2(G2105), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n779), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n777), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n776), .B1(new_n782), .B2(new_n699), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT35), .B(G1991), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n783), .B(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT36), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(KEYINPUT88), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n775), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n771), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT87), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n790), .B(KEYINPUT88), .C1(new_n791), .C2(new_n787), .ZN(new_n792));
  OAI21_X1  g367(.A(KEYINPUT88), .B1(new_n791), .B2(new_n787), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n771), .A2(new_n793), .A3(new_n789), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n756), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(KEYINPUT94), .B1(G5), .B2(G16), .ZN(new_n796));
  OR3_X1    g371(.A1(KEYINPUT94), .A2(G5), .A3(G16), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n796), .B(new_n797), .C1(G301), .C2(new_n673), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(G1961), .Z(new_n799));
  NOR2_X1   g374(.A1(new_n612), .A2(new_n699), .ZN(new_n800));
  NOR4_X1   g375(.A1(new_n679), .A2(new_n795), .A3(new_n799), .A4(new_n800), .ZN(G311));
  NOR2_X1   g376(.A1(new_n679), .A2(new_n795), .ZN(new_n802));
  INV_X1    g377(.A(new_n799), .ZN(new_n803));
  INV_X1    g378(.A(new_n800), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(G150));
  NAND2_X1  g380(.A1(new_n510), .A2(G67), .ZN(new_n806));
  NAND2_X1  g381(.A1(G80), .A2(G543), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n509), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  OAI211_X1 g383(.A(G55), .B(G543), .C1(new_n497), .C2(new_n498), .ZN(new_n809));
  INV_X1    g384(.A(G93), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n507), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(G860), .B1(new_n808), .B2(new_n811), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT37), .Z(new_n813));
  NAND2_X1  g388(.A1(new_n595), .A2(G559), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n806), .A2(new_n807), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n811), .B1(new_n815), .B2(G651), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n535), .A2(G651), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(new_n531), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n536), .B1(new_n808), .B2(new_n811), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n814), .B(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n813), .B1(new_n823), .B2(G860), .ZN(G145));
  INV_X1    g399(.A(KEYINPUT40), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n724), .B(new_n710), .ZN(new_n826));
  INV_X1    g401(.A(new_n495), .ZN(new_n827));
  INV_X1    g402(.A(new_n486), .ZN(new_n828));
  INV_X1    g403(.A(G126), .ZN(new_n829));
  OAI22_X1  g404(.A1(new_n477), .A2(new_n829), .B1(new_n487), .B2(new_n469), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n828), .B1(new_n830), .B2(G2105), .ZN(new_n831));
  AOI21_X1  g406(.A(KEYINPUT95), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT95), .ZN(new_n833));
  NOR3_X1   g408(.A1(new_n490), .A2(new_n495), .A3(new_n833), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n826), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n724), .B(new_n709), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n832), .A2(new_n834), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(new_n686), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n836), .A2(new_n839), .A3(new_n685), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT98), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT97), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT96), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n478), .A2(new_n846), .A3(G130), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n460), .A2(G2105), .ZN(new_n848));
  INV_X1    g423(.A(G130), .ZN(new_n849));
  OAI21_X1  g424(.A(KEYINPUT96), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n480), .A2(G142), .ZN(new_n851));
  OR2_X1    g426(.A1(G106), .A2(G2105), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n852), .B(G2104), .C1(G118), .C2(new_n459), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n847), .A2(new_n850), .A3(new_n851), .A4(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n616), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(new_n782), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n855), .A2(new_n782), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n845), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n858), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n860), .A2(KEYINPUT97), .A3(new_n856), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n843), .A2(new_n844), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n844), .B1(new_n843), .B2(new_n862), .ZN(new_n864));
  OAI22_X1  g439(.A1(new_n863), .A2(new_n864), .B1(new_n862), .B2(new_n843), .ZN(new_n865));
  XNOR2_X1  g440(.A(G162), .B(G160), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n612), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(G37), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT99), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n843), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n841), .A2(KEYINPUT99), .A3(new_n842), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n871), .A2(new_n856), .A3(new_n860), .A4(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n867), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n873), .B(new_n874), .C1(new_n863), .C2(new_n864), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n868), .A2(new_n869), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n876), .A2(KEYINPUT100), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n878));
  AOI21_X1  g453(.A(G37), .B1(new_n865), .B2(new_n867), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n878), .B1(new_n879), .B2(new_n875), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n825), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n876), .A2(KEYINPUT100), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n879), .A2(new_n878), .A3(new_n875), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(KEYINPUT40), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(new_n884), .ZN(G395));
  NAND3_X1  g460(.A1(new_n595), .A2(new_n601), .A3(new_n820), .ZN(new_n886));
  INV_X1    g461(.A(new_n587), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT10), .B1(new_n578), .B2(new_n579), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n889), .A2(KEYINPUT101), .A3(new_n549), .A4(new_n586), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n549), .A2(KEYINPUT101), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT101), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n892), .B1(new_n544), .B2(new_n548), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n588), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT41), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n890), .A2(new_n894), .A3(KEYINPUT41), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n603), .A2(new_n819), .A3(new_n818), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n886), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  AOI22_X1  g476(.A1(new_n886), .A2(new_n900), .B1(new_n890), .B2(new_n894), .ZN(new_n902));
  OAI21_X1  g477(.A(KEYINPUT42), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n886), .A2(new_n900), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n895), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT42), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n886), .A2(new_n899), .A3(new_n900), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n758), .A2(G303), .ZN(new_n909));
  NAND2_X1  g484(.A1(G166), .A2(G288), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI22_X1  g486(.A1(new_n564), .A2(G651), .B1(G86), .B2(new_n545), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n911), .A2(new_n566), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n909), .A2(G305), .A3(new_n910), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  XOR2_X1   g490(.A(new_n574), .B(KEYINPUT102), .Z(new_n916));
  XNOR2_X1  g491(.A(new_n915), .B(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n903), .A2(new_n908), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n918), .B1(new_n903), .B2(new_n908), .ZN(new_n920));
  OAI21_X1  g495(.A(G868), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n921), .B1(G868), .B2(new_n816), .ZN(G295));
  OAI21_X1  g497(.A(new_n921), .B1(G868), .B2(new_n816), .ZN(G331));
  AND3_X1   g498(.A1(G301), .A2(new_n818), .A3(new_n819), .ZN(new_n924));
  AOI21_X1  g499(.A(G301), .B1(new_n818), .B2(new_n819), .ZN(new_n925));
  OAI21_X1  g500(.A(G286), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n820), .A2(G171), .ZN(new_n927));
  NAND3_X1  g502(.A1(G301), .A2(new_n818), .A3(new_n819), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(G168), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n930), .A2(new_n897), .A3(new_n898), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT103), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n930), .A2(new_n897), .A3(KEYINPUT103), .A4(new_n898), .ZN(new_n934));
  OR2_X1    g509(.A1(new_n930), .A2(new_n895), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n933), .A2(new_n917), .A3(new_n934), .A4(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n869), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n930), .A2(new_n895), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n938), .B1(new_n931), .B2(new_n932), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n917), .B1(new_n939), .B2(new_n934), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT43), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n935), .A2(new_n931), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n918), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n943), .A2(new_n936), .A3(new_n944), .A4(new_n869), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n944), .B1(new_n937), .B2(new_n940), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n943), .A2(new_n936), .A3(new_n869), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n947), .B1(new_n944), .B2(new_n948), .ZN(new_n949));
  MUX2_X1   g524(.A(new_n946), .B(new_n949), .S(KEYINPUT44), .Z(G397));
  INV_X1    g525(.A(KEYINPUT45), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n951), .B1(new_n838), .B2(G1384), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n461), .A2(new_n462), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(G2105), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT68), .B1(new_n474), .B2(new_n459), .ZN(new_n955));
  AOI211_X1 g530(.A(new_n464), .B(G2105), .C1(new_n473), .C2(new_n465), .ZN(new_n956));
  OAI211_X1 g531(.A(G40), .B(new_n954), .C1(new_n955), .C2(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n952), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n709), .B(new_n713), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n959), .B(KEYINPUT105), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n724), .B(G1996), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n781), .B(new_n785), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(G290), .A2(G1986), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n965), .A2(KEYINPUT104), .ZN(new_n966));
  NAND2_X1  g541(.A1(G290), .A2(G1986), .ZN(new_n967));
  XOR2_X1   g542(.A(new_n966), .B(new_n967), .Z(new_n968));
  OAI21_X1  g543(.A(new_n958), .B1(new_n964), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G1384), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n970), .B1(new_n490), .B2(new_n495), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n951), .ZN(new_n972));
  INV_X1    g547(.A(G40), .ZN(new_n973));
  AOI211_X1 g548(.A(new_n973), .B(new_n463), .C1(new_n468), .C2(new_n475), .ZN(new_n974));
  INV_X1    g549(.A(G2078), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n975), .A2(KEYINPUT53), .ZN(new_n976));
  OAI211_X1 g551(.A(KEYINPUT45), .B(new_n970), .C1(new_n490), .C2(new_n495), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n972), .A2(new_n974), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n971), .A2(new_n979), .ZN(new_n980));
  OAI211_X1 g555(.A(KEYINPUT50), .B(new_n970), .C1(new_n490), .C2(new_n495), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n957), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n978), .B1(new_n982), .B2(G1961), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT123), .ZN(new_n984));
  OAI211_X1 g559(.A(KEYINPUT45), .B(new_n970), .C1(new_n832), .C2(new_n834), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n957), .B1(new_n951), .B2(new_n971), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n985), .A2(new_n986), .A3(new_n975), .ZN(new_n987));
  NAND2_X1  g562(.A1(KEYINPUT124), .A2(KEYINPUT53), .ZN(new_n988));
  OR2_X1    g563(.A1(KEYINPUT124), .A2(KEYINPUT53), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT123), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n978), .B(new_n991), .C1(new_n982), .C2(G1961), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n984), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(G171), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT125), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT125), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n993), .A2(new_n996), .A3(G171), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n982), .A2(G1961), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n998), .B(KEYINPUT126), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n952), .A2(new_n974), .A3(new_n985), .A4(new_n976), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n999), .A2(G301), .A3(new_n1000), .A4(new_n990), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n995), .A2(new_n997), .A3(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(KEYINPUT122), .B(KEYINPUT54), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n999), .A2(new_n1000), .A3(new_n990), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(G171), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1006), .B(KEYINPUT54), .C1(G171), .C2(new_n993), .ZN(new_n1007));
  AOI21_X1  g582(.A(G1971), .B1(new_n985), .B2(new_n986), .ZN(new_n1008));
  XOR2_X1   g583(.A(KEYINPUT106), .B(G2090), .Z(new_n1009));
  AOI211_X1 g584(.A(new_n957), .B(new_n1009), .C1(new_n980), .C2(new_n981), .ZN(new_n1010));
  OAI21_X1  g585(.A(G8), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g586(.A(KEYINPUT55), .B(G8), .C1(new_n508), .C2(new_n513), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n1012), .B(KEYINPUT107), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n1014));
  INV_X1    g589(.A(G8), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1014), .B1(G166), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT108), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g593(.A(KEYINPUT108), .B(new_n1014), .C1(G166), .C2(new_n1015), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1013), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1011), .B(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G1981), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT110), .B1(new_n564), .B2(G651), .ZN(new_n1023));
  OAI21_X1  g598(.A(G305), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT110), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n565), .A2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1026), .A2(G1981), .A3(new_n566), .A4(new_n912), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1024), .A2(new_n1027), .A3(KEYINPUT111), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT49), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n957), .A2(new_n971), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1030), .A2(new_n1015), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT49), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1024), .A2(new_n1027), .A3(KEYINPUT111), .A4(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1029), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G1976), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1031), .B1(new_n1035), .B2(G288), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT52), .ZN(new_n1037));
  XOR2_X1   g612(.A(KEYINPUT109), .B(G1976), .Z(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT52), .B1(G288), .B2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1031), .B(new_n1039), .C1(new_n1035), .C2(G288), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1034), .A2(new_n1037), .A3(new_n1040), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1021), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n982), .A2(new_n738), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n972), .A2(new_n974), .A3(new_n977), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n717), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1015), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(G286), .A2(G8), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT121), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT51), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1047), .ZN(new_n1050));
  OR3_X1    g625(.A1(new_n1046), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1049), .B1(new_n1046), .B2(new_n1050), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1046), .A2(G286), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1004), .A2(new_n1007), .A3(new_n1042), .A4(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n549), .B(KEYINPUT57), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT115), .B(G2072), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1058), .B(KEYINPUT56), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n985), .A2(new_n986), .A3(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n982), .A2(G1956), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1057), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT118), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT61), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1065), .B(new_n1057), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n985), .A2(new_n986), .A3(new_n1059), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1068), .B(new_n1056), .C1(G1956), .C2(new_n982), .ZN(new_n1069));
  AND2_X1   g644(.A1(KEYINPUT119), .A2(KEYINPUT61), .ZN(new_n1070));
  OR2_X1    g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1062), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1067), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G1996), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n985), .A2(new_n986), .A3(new_n1074), .ZN(new_n1075));
  XOR2_X1   g650(.A(KEYINPUT58), .B(G1341), .Z(new_n1076));
  OAI21_X1  g651(.A(new_n1076), .B1(new_n957), .B2(new_n971), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OAI211_X1 g654(.A(KEYINPUT116), .B(new_n1076), .C1(new_n957), .C2(new_n971), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1075), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT117), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1075), .A2(new_n1083), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1082), .A2(new_n536), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1082), .A2(KEYINPUT59), .A3(new_n536), .A4(new_n1084), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT120), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1073), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1067), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT120), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1030), .A2(new_n713), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n982), .B2(G1348), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT60), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1096), .B1(new_n590), .B2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n590), .A2(new_n1097), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1098), .B(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1091), .A2(new_n1094), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1069), .A2(new_n593), .A3(new_n1096), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1102), .A2(new_n1062), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1055), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1013), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1011), .A2(new_n1105), .A3(KEYINPUT113), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1013), .A2(new_n1018), .A3(KEYINPUT113), .A4(new_n1019), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1107), .B(G8), .C1(new_n1008), .C2(new_n1010), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1106), .A2(new_n1108), .A3(KEYINPUT63), .ZN(new_n1109));
  AOI211_X1 g684(.A(new_n1015), .B(G286), .C1(new_n1043), .C2(new_n1045), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1110), .A2(new_n1037), .A3(new_n1034), .A4(new_n1040), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT114), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1106), .A2(new_n1108), .A3(KEYINPUT63), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT114), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n1114), .A2(new_n1111), .A3(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  OR2_X1    g692(.A1(new_n1011), .A2(new_n1105), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1011), .A2(new_n1105), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1041), .A2(new_n1118), .A3(new_n1119), .A4(new_n1110), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT112), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT63), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1021), .A2(KEYINPUT112), .A3(new_n1041), .A4(new_n1110), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1122), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1117), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1118), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1127), .A2(new_n1041), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT62), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1051), .A2(new_n1129), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1130), .A2(new_n1021), .A3(new_n1041), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1054), .A2(KEYINPUT62), .B1(new_n995), .B2(new_n997), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1128), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1034), .A2(new_n1035), .A3(new_n758), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(G1981), .B2(G305), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n1031), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1126), .A2(new_n1133), .A3(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n969), .B1(new_n1104), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n958), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n962), .A2(new_n785), .A3(new_n782), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n710), .A2(new_n713), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1139), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT46), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1143), .B1(new_n1139), .B2(G1996), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n958), .B1(new_n960), .B2(new_n724), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n958), .A2(KEYINPUT46), .A3(new_n1074), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  XOR2_X1   g722(.A(new_n1147), .B(KEYINPUT47), .Z(new_n1148));
  NAND2_X1  g723(.A1(new_n964), .A2(new_n958), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n958), .A2(new_n965), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1150), .B(KEYINPUT48), .ZN(new_n1151));
  AOI211_X1 g726(.A(new_n1142), .B(new_n1148), .C1(new_n1149), .C2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1138), .A2(new_n1152), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g728(.A1(new_n670), .A2(G319), .A3(new_n671), .ZN(new_n1155));
  INV_X1    g729(.A(new_n1155), .ZN(new_n1156));
  AOI21_X1  g730(.A(G227), .B1(new_n637), .B2(G14), .ZN(new_n1157));
  NAND4_X1  g731(.A1(new_n946), .A2(new_n876), .A3(new_n1156), .A4(new_n1157), .ZN(G225));
  INV_X1    g732(.A(KEYINPUT127), .ZN(new_n1159));
  NAND2_X1  g733(.A1(G225), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g734(.A(new_n1155), .B1(new_n941), .B2(new_n945), .ZN(new_n1161));
  NAND4_X1  g735(.A1(new_n1161), .A2(KEYINPUT127), .A3(new_n876), .A4(new_n1157), .ZN(new_n1162));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1162), .ZN(G308));
endmodule


