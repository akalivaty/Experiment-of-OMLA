

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761;

  INV_X1 U374 ( .A(n513), .ZN(n692) );
  XNOR2_X1 U375 ( .A(n744), .B(n432), .ZN(n658) );
  XNOR2_X2 U376 ( .A(n510), .B(n509), .ZN(n540) );
  NAND2_X1 U377 ( .A1(n374), .A2(n371), .ZN(n370) );
  XNOR2_X2 U378 ( .A(n446), .B(n445), .ZN(n513) );
  XNOR2_X2 U379 ( .A(n464), .B(n355), .ZN(n567) );
  XNOR2_X2 U380 ( .A(n596), .B(KEYINPUT40), .ZN(n761) );
  AND2_X2 U381 ( .A1(n618), .A2(n680), .ZN(n596) );
  NAND2_X1 U382 ( .A1(n671), .A2(n543), .ZN(n382) );
  AND2_X1 U383 ( .A1(n576), .A2(n575), .ZN(n593) );
  XNOR2_X1 U384 ( .A(n419), .B(n418), .ZN(n551) );
  XNOR2_X1 U385 ( .A(n452), .B(G134), .ZN(n490) );
  XNOR2_X1 U386 ( .A(KEYINPUT8), .B(KEYINPUT71), .ZN(n409) );
  XNOR2_X2 U387 ( .A(n385), .B(KEYINPUT35), .ZN(n636) );
  NAND2_X1 U388 ( .A1(n353), .A2(n352), .ZN(n525) );
  INV_X1 U389 ( .A(n524), .ZN(n352) );
  INV_X1 U390 ( .A(n636), .ZN(n353) );
  INV_X1 U391 ( .A(n541), .ZN(n354) );
  XNOR2_X1 U392 ( .A(n523), .B(n522), .ZN(n760) );
  XNOR2_X1 U393 ( .A(n375), .B(KEYINPUT87), .ZN(n374) );
  BUF_X1 U394 ( .A(n567), .Z(n617) );
  XNOR2_X2 U395 ( .A(n629), .B(n628), .ZN(n361) );
  XNOR2_X2 U396 ( .A(n370), .B(n545), .ZN(n360) );
  XNOR2_X2 U397 ( .A(n475), .B(KEYINPUT0), .ZN(n528) );
  INV_X1 U398 ( .A(KEYINPUT77), .ZN(n387) );
  NAND2_X1 U399 ( .A1(n395), .A2(n627), .ZN(n393) );
  OR2_X1 U400 ( .A1(n396), .A2(n623), .ZN(n395) );
  OR2_X1 U401 ( .A1(n622), .A2(n624), .ZN(n396) );
  INV_X1 U402 ( .A(n667), .ZN(n368) );
  XNOR2_X1 U403 ( .A(n364), .B(n363), .ZN(n379) );
  INV_X1 U404 ( .A(KEYINPUT108), .ZN(n363) );
  NOR2_X1 U405 ( .A1(n382), .A2(n387), .ZN(n376) );
  INV_X1 U406 ( .A(KEYINPUT2), .ZN(n391) );
  XNOR2_X1 U407 ( .A(n607), .B(KEYINPUT48), .ZN(n608) );
  NOR2_X1 U408 ( .A1(n606), .A2(n605), .ZN(n609) );
  NOR2_X1 U409 ( .A1(n692), .A2(n611), .ZN(n573) );
  XNOR2_X1 U410 ( .A(n417), .B(n416), .ZN(n418) );
  INV_X1 U411 ( .A(n570), .ZN(n507) );
  XOR2_X1 U412 ( .A(KEYINPUT106), .B(n506), .Z(n710) );
  AND2_X1 U413 ( .A1(n593), .A2(n707), .ZN(n595) );
  XNOR2_X1 U414 ( .A(n630), .B(n633), .ZN(n634) );
  NAND2_X1 U415 ( .A1(n366), .A2(n365), .ZN(n364) );
  INV_X1 U416 ( .A(n665), .ZN(n365) );
  NOR2_X1 U417 ( .A1(G953), .A2(G237), .ZN(n480) );
  INV_X1 U418 ( .A(G128), .ZN(n423) );
  XNOR2_X1 U419 ( .A(KEYINPUT73), .B(G131), .ZN(n483) );
  XNOR2_X1 U420 ( .A(G113), .B(G143), .ZN(n477) );
  XNOR2_X1 U421 ( .A(n454), .B(n453), .ZN(n456) );
  XNOR2_X1 U422 ( .A(KEYINPUT4), .B(G146), .ZN(n454) );
  NAND2_X1 U423 ( .A1(G234), .A2(G237), .ZN(n469) );
  NAND2_X1 U424 ( .A1(n373), .A2(n372), .ZN(n371) );
  NAND2_X1 U425 ( .A1(n377), .A2(n387), .ZN(n373) );
  XNOR2_X1 U426 ( .A(n467), .B(KEYINPUT79), .ZN(n468) );
  XNOR2_X1 U427 ( .A(n531), .B(KEYINPUT1), .ZN(n511) );
  XNOR2_X1 U428 ( .A(KEYINPUT5), .B(G146), .ZN(n435) );
  XOR2_X1 U429 ( .A(KEYINPUT70), .B(G101), .Z(n438) );
  XNOR2_X1 U430 ( .A(G116), .B(G113), .ZN(n439) );
  XNOR2_X1 U431 ( .A(G119), .B(G128), .ZN(n407) );
  XNOR2_X1 U432 ( .A(n400), .B(KEYINPUT72), .ZN(n745) );
  XNOR2_X1 U433 ( .A(G146), .B(G125), .ZN(n399) );
  NAND2_X2 U434 ( .A1(n392), .A2(n390), .ZN(n629) );
  NAND2_X1 U435 ( .A1(n389), .A2(n388), .ZN(n390) );
  NOR2_X1 U436 ( .A1(n746), .A2(n391), .ZN(n388) );
  OR2_X2 U437 ( .A1(n623), .A2(n622), .ZN(n746) );
  AND2_X1 U438 ( .A1(n532), .A2(n574), .ZN(n575) );
  XOR2_X1 U439 ( .A(KEYINPUT22), .B(KEYINPUT66), .Z(n509) );
  INV_X2 U440 ( .A(G953), .ZN(n747) );
  XNOR2_X1 U441 ( .A(n362), .B(n530), .ZN(n684) );
  INV_X1 U442 ( .A(KEYINPUT56), .ZN(n356) );
  NAND2_X1 U443 ( .A1(n358), .A2(n653), .ZN(n357) );
  XNOR2_X1 U444 ( .A(n359), .B(n634), .ZN(n358) );
  AND2_X1 U445 ( .A1(G210), .A2(n465), .ZN(n355) );
  XNOR2_X1 U446 ( .A(G902), .B(KEYINPUT15), .ZN(n624) );
  XNOR2_X1 U447 ( .A(n357), .B(n356), .ZN(G51) );
  NAND2_X1 U448 ( .A1(n649), .A2(G210), .ZN(n359) );
  XNOR2_X1 U449 ( .A(n370), .B(n545), .ZN(n734) );
  XNOR2_X1 U450 ( .A(n629), .B(n628), .ZN(n649) );
  XNOR2_X1 U451 ( .A(n384), .B(n449), .ZN(n704) );
  NAND2_X1 U452 ( .A1(n528), .A2(n698), .ZN(n362) );
  NAND2_X1 U453 ( .A1(n369), .A2(n368), .ZN(n367) );
  NAND2_X1 U454 ( .A1(n367), .A2(n581), .ZN(n366) );
  INV_X1 U455 ( .A(n684), .ZN(n369) );
  NAND2_X1 U456 ( .A1(n376), .A2(n544), .ZN(n372) );
  NAND2_X1 U457 ( .A1(n378), .A2(n379), .ZN(n375) );
  NAND2_X1 U458 ( .A1(n381), .A2(n544), .ZN(n377) );
  NAND2_X1 U459 ( .A1(n525), .A2(KEYINPUT44), .ZN(n378) );
  NAND2_X1 U460 ( .A1(n511), .A2(n694), .ZN(n529) );
  XNOR2_X2 U461 ( .A(n380), .B(n434), .ZN(n531) );
  NAND2_X1 U462 ( .A1(n658), .A2(n499), .ZN(n380) );
  INV_X1 U463 ( .A(n382), .ZN(n381) );
  XNOR2_X1 U464 ( .A(n383), .B(n476), .ZN(n386) );
  NAND2_X1 U465 ( .A1(n536), .A2(n704), .ZN(n383) );
  NAND2_X1 U466 ( .A1(n448), .A2(n555), .ZN(n384) );
  XNOR2_X1 U467 ( .A(n528), .B(KEYINPUT94), .ZN(n536) );
  NAND2_X1 U468 ( .A1(n386), .A2(n578), .ZN(n385) );
  INV_X1 U469 ( .A(n734), .ZN(n389) );
  NAND2_X1 U470 ( .A1(n360), .A2(n627), .ZN(n394) );
  NOR2_X1 U471 ( .A1(n734), .A2(n746), .ZN(n687) );
  AND2_X2 U472 ( .A1(n394), .A2(n393), .ZN(n392) );
  XOR2_X1 U473 ( .A(n483), .B(n425), .Z(n397) );
  INV_X1 U474 ( .A(G125), .ZN(n453) );
  INV_X1 U475 ( .A(KEYINPUT86), .ZN(n607) );
  INV_X1 U476 ( .A(KEYINPUT10), .ZN(n398) );
  XNOR2_X1 U477 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U478 ( .A(n405), .B(n404), .ZN(n406) );
  NOR2_X1 U479 ( .A1(n710), .A2(n507), .ZN(n508) );
  XNOR2_X1 U480 ( .A(n489), .B(n488), .ZN(n527) );
  INV_X1 U481 ( .A(KEYINPUT74), .ZN(n401) );
  XNOR2_X1 U482 ( .A(n401), .B(G140), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n426), .B(KEYINPUT23), .ZN(n405) );
  XOR2_X1 U484 ( .A(KEYINPUT97), .B(KEYINPUT24), .Z(n403) );
  XNOR2_X1 U485 ( .A(KEYINPUT98), .B(KEYINPUT96), .ZN(n402) );
  XNOR2_X1 U486 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U487 ( .A(n745), .B(n406), .ZN(n414) );
  XOR2_X1 U488 ( .A(G110), .B(G137), .Z(n408) );
  XNOR2_X1 U489 ( .A(n408), .B(n407), .ZN(n412) );
  NAND2_X1 U490 ( .A1(n747), .A2(G234), .ZN(n410) );
  XNOR2_X1 U491 ( .A(n410), .B(n409), .ZN(n491) );
  NAND2_X1 U492 ( .A1(G221), .A2(n491), .ZN(n411) );
  XOR2_X1 U493 ( .A(n412), .B(n411), .Z(n413) );
  XNOR2_X1 U494 ( .A(n414), .B(n413), .ZN(n643) );
  NOR2_X1 U495 ( .A1(G902), .A2(n643), .ZN(n419) );
  NAND2_X1 U496 ( .A1(G234), .A2(n624), .ZN(n415) );
  XNOR2_X1 U497 ( .A(KEYINPUT20), .B(n415), .ZN(n420) );
  NAND2_X1 U498 ( .A1(G217), .A2(n420), .ZN(n417) );
  XNOR2_X1 U499 ( .A(KEYINPUT25), .B(KEYINPUT80), .ZN(n416) );
  NAND2_X1 U500 ( .A1(G221), .A2(n420), .ZN(n421) );
  XOR2_X1 U501 ( .A(KEYINPUT21), .B(n421), .Z(n688) );
  INV_X1 U502 ( .A(KEYINPUT99), .ZN(n422) );
  XNOR2_X1 U503 ( .A(n688), .B(n422), .ZN(n570) );
  AND2_X1 U504 ( .A1(n551), .A2(n570), .ZN(n694) );
  XNOR2_X2 U505 ( .A(G143), .B(KEYINPUT82), .ZN(n424) );
  XNOR2_X2 U506 ( .A(n424), .B(n423), .ZN(n452) );
  XNOR2_X1 U507 ( .A(KEYINPUT4), .B(G137), .ZN(n425) );
  XNOR2_X2 U508 ( .A(n490), .B(n397), .ZN(n444) );
  XNOR2_X1 U509 ( .A(n426), .B(KEYINPUT95), .ZN(n427) );
  XNOR2_X2 U510 ( .A(n444), .B(n427), .ZN(n744) );
  XNOR2_X1 U511 ( .A(G104), .B(G110), .ZN(n428) );
  XNOR2_X1 U512 ( .A(n428), .B(G107), .ZN(n729) );
  XNOR2_X1 U513 ( .A(n438), .B(KEYINPUT76), .ZN(n429) );
  XNOR2_X1 U514 ( .A(n729), .B(n429), .ZN(n459) );
  NAND2_X1 U515 ( .A1(n747), .A2(G227), .ZN(n430) );
  XNOR2_X1 U516 ( .A(n430), .B(G146), .ZN(n431) );
  XNOR2_X1 U517 ( .A(n459), .B(n431), .ZN(n432) );
  INV_X1 U518 ( .A(G902), .ZN(n499) );
  INV_X1 U519 ( .A(KEYINPUT75), .ZN(n433) );
  XNOR2_X1 U520 ( .A(n433), .B(G469), .ZN(n434) );
  XNOR2_X1 U521 ( .A(n529), .B(KEYINPUT109), .ZN(n448) );
  NAND2_X1 U522 ( .A1(n480), .A2(G210), .ZN(n436) );
  XNOR2_X1 U523 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U524 ( .A(n438), .B(n437), .ZN(n442) );
  XNOR2_X1 U525 ( .A(n439), .B(KEYINPUT3), .ZN(n441) );
  XOR2_X1 U526 ( .A(KEYINPUT90), .B(G119), .Z(n440) );
  XNOR2_X1 U527 ( .A(n441), .B(n440), .ZN(n462) );
  XNOR2_X1 U528 ( .A(n442), .B(n462), .ZN(n443) );
  XNOR2_X1 U529 ( .A(n444), .B(n443), .ZN(n638) );
  NAND2_X1 U530 ( .A1(n638), .A2(n499), .ZN(n446) );
  XNOR2_X1 U531 ( .A(G472), .B(KEYINPUT100), .ZN(n445) );
  XNOR2_X1 U532 ( .A(KEYINPUT105), .B(KEYINPUT6), .ZN(n447) );
  XNOR2_X1 U533 ( .A(n692), .B(n447), .ZN(n537) );
  INV_X1 U534 ( .A(n537), .ZN(n555) );
  XNOR2_X1 U535 ( .A(KEYINPUT110), .B(KEYINPUT33), .ZN(n449) );
  NAND2_X1 U536 ( .A1(G224), .A2(n747), .ZN(n450) );
  XNOR2_X1 U537 ( .A(n450), .B(KEYINPUT17), .ZN(n451) );
  XNOR2_X1 U538 ( .A(n452), .B(n451), .ZN(n458) );
  INV_X1 U539 ( .A(KEYINPUT18), .ZN(n455) );
  XNOR2_X1 U540 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U541 ( .A(n458), .B(n457), .ZN(n460) );
  XNOR2_X1 U542 ( .A(n460), .B(n459), .ZN(n463) );
  XNOR2_X1 U543 ( .A(KEYINPUT16), .B(G122), .ZN(n461) );
  XNOR2_X1 U544 ( .A(n462), .B(n461), .ZN(n730) );
  XNOR2_X1 U545 ( .A(n463), .B(n730), .ZN(n630) );
  NAND2_X1 U546 ( .A1(n630), .A2(n624), .ZN(n464) );
  OR2_X1 U547 ( .A1(G237), .A2(G902), .ZN(n465) );
  NAND2_X1 U548 ( .A1(n465), .A2(G214), .ZN(n466) );
  XOR2_X1 U549 ( .A(n466), .B(KEYINPUT91), .Z(n706) );
  NAND2_X1 U550 ( .A1(n567), .A2(n706), .ZN(n546) );
  XNOR2_X1 U551 ( .A(KEYINPUT19), .B(KEYINPUT68), .ZN(n467) );
  XNOR2_X1 U552 ( .A(n546), .B(n468), .ZN(n563) );
  XNOR2_X1 U553 ( .A(n469), .B(KEYINPUT14), .ZN(n471) );
  NAND2_X1 U554 ( .A1(G952), .A2(n471), .ZN(n470) );
  XNOR2_X1 U555 ( .A(KEYINPUT92), .B(n470), .ZN(n721) );
  NOR2_X1 U556 ( .A1(G953), .A2(n721), .ZN(n550) );
  NAND2_X1 U557 ( .A1(G902), .A2(n471), .ZN(n547) );
  NOR2_X1 U558 ( .A1(G898), .A2(n747), .ZN(n472) );
  XNOR2_X1 U559 ( .A(KEYINPUT93), .B(n472), .ZN(n732) );
  NOR2_X1 U560 ( .A1(n547), .A2(n732), .ZN(n473) );
  NOR2_X1 U561 ( .A1(n550), .A2(n473), .ZN(n474) );
  NOR2_X2 U562 ( .A1(n563), .A2(n474), .ZN(n475) );
  INV_X1 U563 ( .A(KEYINPUT34), .ZN(n476) );
  XOR2_X1 U564 ( .A(G122), .B(G104), .Z(n478) );
  XNOR2_X1 U565 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U566 ( .A(n745), .B(n479), .ZN(n487) );
  XOR2_X1 U567 ( .A(G140), .B(KEYINPUT11), .Z(n482) );
  NAND2_X1 U568 ( .A1(G214), .A2(n480), .ZN(n481) );
  XNOR2_X1 U569 ( .A(n482), .B(n481), .ZN(n485) );
  XNOR2_X1 U570 ( .A(n483), .B(KEYINPUT12), .ZN(n484) );
  XNOR2_X1 U571 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U572 ( .A(n487), .B(n486), .ZN(n650) );
  NAND2_X1 U573 ( .A1(n650), .A2(n499), .ZN(n489) );
  XNOR2_X1 U574 ( .A(KEYINPUT13), .B(G475), .ZN(n488) );
  INV_X1 U575 ( .A(n527), .ZN(n504) );
  XOR2_X1 U576 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n493) );
  NAND2_X1 U577 ( .A1(G217), .A2(n491), .ZN(n492) );
  XNOR2_X1 U578 ( .A(n493), .B(n492), .ZN(n497) );
  XOR2_X1 U579 ( .A(KEYINPUT102), .B(G122), .Z(n495) );
  XNOR2_X1 U580 ( .A(G116), .B(G107), .ZN(n494) );
  XNOR2_X1 U581 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U582 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U583 ( .A(n490), .B(n498), .ZN(n647) );
  NAND2_X1 U584 ( .A1(n647), .A2(n499), .ZN(n503) );
  XNOR2_X1 U585 ( .A(KEYINPUT103), .B(KEYINPUT104), .ZN(n501) );
  INV_X1 U586 ( .A(G478), .ZN(n500) );
  XNOR2_X1 U587 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U588 ( .A(n503), .B(n502), .ZN(n526) );
  AND2_X1 U589 ( .A1(n504), .A2(n526), .ZN(n578) );
  INV_X1 U590 ( .A(n526), .ZN(n505) );
  AND2_X1 U591 ( .A1(n527), .A2(n505), .ZN(n506) );
  NAND2_X1 U592 ( .A1(n528), .A2(n508), .ZN(n510) );
  BUF_X1 U593 ( .A(n511), .Z(n512) );
  NOR2_X1 U594 ( .A1(n512), .A2(n513), .ZN(n514) );
  NAND2_X1 U595 ( .A1(n540), .A2(n514), .ZN(n515) );
  XNOR2_X1 U596 ( .A(n515), .B(KEYINPUT65), .ZN(n516) );
  INV_X1 U597 ( .A(n551), .ZN(n572) );
  NAND2_X1 U598 ( .A1(n516), .A2(n572), .ZN(n542) );
  INV_X1 U599 ( .A(KEYINPUT107), .ZN(n517) );
  XNOR2_X1 U600 ( .A(n551), .B(n517), .ZN(n689) );
  INV_X1 U601 ( .A(n689), .ZN(n519) );
  AND2_X1 U602 ( .A1(n512), .A2(n537), .ZN(n518) );
  AND2_X1 U603 ( .A1(n519), .A2(n518), .ZN(n520) );
  NAND2_X1 U604 ( .A1(n540), .A2(n520), .ZN(n523) );
  INV_X1 U605 ( .A(KEYINPUT81), .ZN(n521) );
  XNOR2_X1 U606 ( .A(n521), .B(KEYINPUT32), .ZN(n522) );
  NAND2_X1 U607 ( .A1(n542), .A2(n760), .ZN(n524) );
  AND2_X1 U608 ( .A1(n527), .A2(n526), .ZN(n683) );
  NOR2_X1 U609 ( .A1(n527), .A2(n526), .ZN(n680) );
  NOR2_X1 U610 ( .A1(n683), .A2(n680), .ZN(n712) );
  XOR2_X1 U611 ( .A(KEYINPUT31), .B(KEYINPUT101), .Z(n530) );
  NOR2_X1 U612 ( .A1(n529), .A2(n692), .ZN(n698) );
  NAND2_X1 U613 ( .A1(n694), .A2(n692), .ZN(n534) );
  BUF_X1 U614 ( .A(n531), .Z(n532) );
  INV_X1 U615 ( .A(n532), .ZN(n533) );
  NOR2_X1 U616 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U617 ( .A1(n536), .A2(n535), .ZN(n667) );
  NAND2_X1 U618 ( .A1(n689), .A2(n537), .ZN(n538) );
  NOR2_X1 U619 ( .A1(n538), .A2(n512), .ZN(n539) );
  AND2_X1 U620 ( .A1(n540), .A2(n539), .ZN(n665) );
  INV_X1 U621 ( .A(n760), .ZN(n541) );
  NOR2_X1 U622 ( .A1(n636), .A2(n541), .ZN(n544) );
  BUF_X1 U623 ( .A(n542), .Z(n671) );
  INV_X1 U624 ( .A(KEYINPUT44), .ZN(n543) );
  XNOR2_X1 U625 ( .A(KEYINPUT85), .B(KEYINPUT45), .ZN(n545) );
  INV_X1 U626 ( .A(KEYINPUT111), .ZN(n557) );
  INV_X1 U627 ( .A(n680), .ZN(n553) );
  OR2_X1 U628 ( .A1(n747), .A2(n547), .ZN(n548) );
  NOR2_X1 U629 ( .A1(G900), .A2(n548), .ZN(n549) );
  NOR2_X1 U630 ( .A1(n550), .A2(n549), .ZN(n568) );
  NOR2_X1 U631 ( .A1(n551), .A2(n568), .ZN(n552) );
  NAND2_X1 U632 ( .A1(n552), .A2(n688), .ZN(n561) );
  NOR2_X1 U633 ( .A1(n553), .A2(n561), .ZN(n554) );
  NAND2_X1 U634 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U635 ( .A(n557), .B(n556), .ZN(n610) );
  NOR2_X1 U636 ( .A1(n546), .A2(n610), .ZN(n558) );
  XNOR2_X1 U637 ( .A(KEYINPUT36), .B(n558), .ZN(n559) );
  NAND2_X1 U638 ( .A1(n559), .A2(n512), .ZN(n560) );
  XNOR2_X1 U639 ( .A(n560), .B(KEYINPUT114), .ZN(n758) );
  NOR2_X1 U640 ( .A1(n561), .A2(n692), .ZN(n562) );
  XNOR2_X1 U641 ( .A(n562), .B(KEYINPUT28), .ZN(n600) );
  INV_X1 U642 ( .A(n563), .ZN(n564) );
  AND2_X1 U643 ( .A1(n532), .A2(n564), .ZN(n585) );
  NAND2_X1 U644 ( .A1(n600), .A2(n585), .ZN(n565) );
  NAND2_X1 U645 ( .A1(n565), .A2(KEYINPUT47), .ZN(n566) );
  NAND2_X1 U646 ( .A1(n566), .A2(KEYINPUT83), .ZN(n580) );
  INV_X1 U647 ( .A(n568), .ZN(n569) );
  NAND2_X1 U648 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U649 ( .A1(n572), .A2(n571), .ZN(n576) );
  INV_X1 U650 ( .A(n706), .ZN(n611) );
  XNOR2_X1 U651 ( .A(n573), .B(KEYINPUT30), .ZN(n574) );
  NAND2_X1 U652 ( .A1(n617), .A2(n593), .ZN(n577) );
  XNOR2_X1 U653 ( .A(KEYINPUT113), .B(n577), .ZN(n579) );
  NAND2_X1 U654 ( .A1(n579), .A2(n578), .ZN(n678) );
  NAND2_X1 U655 ( .A1(n580), .A2(n678), .ZN(n591) );
  INV_X1 U656 ( .A(n712), .ZN(n581) );
  AND2_X1 U657 ( .A1(n585), .A2(n581), .ZN(n582) );
  NAND2_X1 U658 ( .A1(n600), .A2(n582), .ZN(n583) );
  NOR2_X1 U659 ( .A1(KEYINPUT47), .A2(n583), .ZN(n584) );
  XOR2_X1 U660 ( .A(n584), .B(KEYINPUT78), .Z(n589) );
  AND2_X1 U661 ( .A1(n600), .A2(n585), .ZN(n674) );
  NOR2_X1 U662 ( .A1(n674), .A2(KEYINPUT83), .ZN(n586) );
  OR2_X1 U663 ( .A1(n712), .A2(n586), .ZN(n587) );
  NAND2_X1 U664 ( .A1(KEYINPUT47), .A2(n587), .ZN(n588) );
  NAND2_X1 U665 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U666 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U667 ( .A1(n758), .A2(n592), .ZN(n606) );
  XOR2_X1 U668 ( .A(KEYINPUT38), .B(n617), .Z(n597) );
  BUF_X1 U669 ( .A(n597), .Z(n707) );
  INV_X1 U670 ( .A(KEYINPUT39), .ZN(n594) );
  XNOR2_X1 U671 ( .A(n595), .B(n594), .ZN(n618) );
  NAND2_X1 U672 ( .A1(n597), .A2(n706), .ZN(n711) );
  NOR2_X1 U673 ( .A1(n711), .A2(n710), .ZN(n599) );
  INV_X1 U674 ( .A(KEYINPUT41), .ZN(n598) );
  XNOR2_X1 U675 ( .A(n599), .B(n598), .ZN(n722) );
  AND2_X1 U676 ( .A1(n600), .A2(n532), .ZN(n601) );
  AND2_X1 U677 ( .A1(n722), .A2(n601), .ZN(n602) );
  XNOR2_X1 U678 ( .A(n602), .B(KEYINPUT42), .ZN(n756) );
  NOR2_X1 U679 ( .A1(n761), .A2(n756), .ZN(n603) );
  XNOR2_X1 U680 ( .A(KEYINPUT46), .B(n603), .ZN(n604) );
  INV_X1 U681 ( .A(n604), .ZN(n605) );
  XNOR2_X1 U682 ( .A(n609), .B(n608), .ZN(n623) );
  INV_X1 U683 ( .A(n610), .ZN(n613) );
  NOR2_X1 U684 ( .A1(n512), .A2(n611), .ZN(n612) );
  NAND2_X1 U685 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U686 ( .A(KEYINPUT43), .B(n614), .ZN(n615) );
  XOR2_X1 U687 ( .A(KEYINPUT112), .B(n615), .Z(n616) );
  NOR2_X1 U688 ( .A1(n617), .A2(n616), .ZN(n686) );
  INV_X1 U689 ( .A(n686), .ZN(n621) );
  NAND2_X1 U690 ( .A1(n618), .A2(n683), .ZN(n620) );
  INV_X1 U691 ( .A(KEYINPUT115), .ZN(n619) );
  XNOR2_X1 U692 ( .A(n620), .B(n619), .ZN(n757) );
  NAND2_X1 U693 ( .A1(n621), .A2(n757), .ZN(n622) );
  XOR2_X1 U694 ( .A(KEYINPUT84), .B(n624), .Z(n625) );
  NAND2_X1 U695 ( .A1(n625), .A2(KEYINPUT2), .ZN(n626) );
  XOR2_X1 U696 ( .A(KEYINPUT67), .B(n626), .Z(n627) );
  INV_X1 U697 ( .A(KEYINPUT64), .ZN(n628) );
  XOR2_X1 U698 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n632) );
  XNOR2_X1 U699 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n631) );
  XOR2_X1 U700 ( .A(n632), .B(n631), .Z(n633) );
  INV_X1 U701 ( .A(G952), .ZN(n635) );
  NAND2_X1 U702 ( .A1(n635), .A2(G953), .ZN(n653) );
  BUF_X1 U703 ( .A(n636), .Z(n637) );
  XOR2_X1 U704 ( .A(n637), .B(G122), .Z(G24) );
  NAND2_X1 U705 ( .A1(n361), .A2(G472), .ZN(n640) );
  XNOR2_X1 U706 ( .A(n638), .B(KEYINPUT62), .ZN(n639) );
  XNOR2_X1 U707 ( .A(n640), .B(n639), .ZN(n641) );
  NAND2_X1 U708 ( .A1(n641), .A2(n653), .ZN(n642) );
  XNOR2_X1 U709 ( .A(n642), .B(KEYINPUT63), .ZN(G57) );
  BUF_X1 U710 ( .A(n649), .Z(n657) );
  NAND2_X1 U711 ( .A1(n657), .A2(G217), .ZN(n644) );
  XNOR2_X1 U712 ( .A(n644), .B(n643), .ZN(n645) );
  INV_X1 U713 ( .A(n653), .ZN(n663) );
  NOR2_X1 U714 ( .A1(n645), .A2(n663), .ZN(G66) );
  NAND2_X1 U715 ( .A1(n361), .A2(G478), .ZN(n646) );
  XOR2_X1 U716 ( .A(n647), .B(n646), .Z(n648) );
  NOR2_X1 U717 ( .A1(n648), .A2(n663), .ZN(G63) );
  NAND2_X1 U718 ( .A1(n361), .A2(G475), .ZN(n652) );
  XOR2_X1 U719 ( .A(n650), .B(KEYINPUT59), .Z(n651) );
  XNOR2_X1 U720 ( .A(n652), .B(n651), .ZN(n654) );
  NAND2_X1 U721 ( .A1(n654), .A2(n653), .ZN(n656) );
  XNOR2_X1 U722 ( .A(KEYINPUT69), .B(KEYINPUT60), .ZN(n655) );
  XNOR2_X1 U723 ( .A(n656), .B(n655), .ZN(G60) );
  NAND2_X1 U724 ( .A1(n657), .A2(G469), .ZN(n662) );
  BUF_X1 U725 ( .A(n658), .Z(n659) );
  XNOR2_X1 U726 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n660) );
  XNOR2_X1 U727 ( .A(n659), .B(n660), .ZN(n661) );
  XNOR2_X1 U728 ( .A(n662), .B(n661), .ZN(n664) );
  NOR2_X1 U729 ( .A1(n664), .A2(n663), .ZN(G54) );
  XOR2_X1 U730 ( .A(G101), .B(n665), .Z(G3) );
  NAND2_X1 U731 ( .A1(n680), .A2(n667), .ZN(n666) );
  XNOR2_X1 U732 ( .A(G104), .B(n666), .ZN(G6) );
  XOR2_X1 U733 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n669) );
  NAND2_X1 U734 ( .A1(n667), .A2(n683), .ZN(n668) );
  XNOR2_X1 U735 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U736 ( .A(G107), .B(n670), .ZN(G9) );
  INV_X1 U737 ( .A(n671), .ZN(n672) );
  XOR2_X1 U738 ( .A(G110), .B(n672), .Z(n673) );
  XNOR2_X1 U739 ( .A(KEYINPUT116), .B(n673), .ZN(G12) );
  XOR2_X1 U740 ( .A(G128), .B(KEYINPUT29), .Z(n676) );
  NAND2_X1 U741 ( .A1(n674), .A2(n683), .ZN(n675) );
  XNOR2_X1 U742 ( .A(n676), .B(n675), .ZN(G30) );
  XOR2_X1 U743 ( .A(G143), .B(KEYINPUT117), .Z(n677) );
  XNOR2_X1 U744 ( .A(n678), .B(n677), .ZN(G45) );
  NAND2_X1 U745 ( .A1(n674), .A2(n680), .ZN(n679) );
  XNOR2_X1 U746 ( .A(n679), .B(G146), .ZN(G48) );
  NAND2_X1 U747 ( .A1(n684), .A2(n680), .ZN(n681) );
  XNOR2_X1 U748 ( .A(n681), .B(KEYINPUT118), .ZN(n682) );
  XNOR2_X1 U749 ( .A(G113), .B(n682), .ZN(G15) );
  NAND2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U751 ( .A(n685), .B(G116), .ZN(G18) );
  XOR2_X1 U752 ( .A(G140), .B(n686), .Z(G42) );
  XOR2_X1 U753 ( .A(KEYINPUT2), .B(n687), .Z(n726) );
  INV_X1 U754 ( .A(n722), .ZN(n702) );
  NOR2_X1 U755 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U756 ( .A(KEYINPUT119), .B(n690), .Z(n691) );
  XNOR2_X1 U757 ( .A(KEYINPUT49), .B(n691), .ZN(n693) );
  NAND2_X1 U758 ( .A1(n693), .A2(n692), .ZN(n697) );
  NOR2_X1 U759 ( .A1(n694), .A2(n512), .ZN(n695) );
  XNOR2_X1 U760 ( .A(n695), .B(KEYINPUT50), .ZN(n696) );
  NOR2_X1 U761 ( .A1(n697), .A2(n696), .ZN(n699) );
  NOR2_X1 U762 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U763 ( .A(KEYINPUT51), .B(n700), .Z(n701) );
  NOR2_X1 U764 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U765 ( .A(n703), .B(KEYINPUT120), .ZN(n718) );
  BUF_X1 U766 ( .A(n704), .Z(n705) );
  INV_X1 U767 ( .A(n705), .ZN(n716) );
  NOR2_X1 U768 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U769 ( .A(KEYINPUT121), .B(n708), .Z(n709) );
  NOR2_X1 U770 ( .A1(n710), .A2(n709), .ZN(n714) );
  NOR2_X1 U771 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U772 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U773 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U774 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U775 ( .A(n719), .B(KEYINPUT52), .ZN(n720) );
  NOR2_X1 U776 ( .A1(n721), .A2(n720), .ZN(n724) );
  AND2_X1 U777 ( .A1(n705), .A2(n722), .ZN(n723) );
  OR2_X1 U778 ( .A1(n724), .A2(n723), .ZN(n725) );
  OR2_X1 U779 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U780 ( .A1(n727), .A2(G953), .ZN(n728) );
  XNOR2_X1 U781 ( .A(n728), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U782 ( .A(G101), .B(n729), .ZN(n731) );
  XNOR2_X1 U783 ( .A(n731), .B(n730), .ZN(n733) );
  NAND2_X1 U784 ( .A1(n733), .A2(n732), .ZN(n743) );
  NOR2_X1 U785 ( .A1(n360), .A2(G953), .ZN(n741) );
  XOR2_X1 U786 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n736) );
  NAND2_X1 U787 ( .A1(G224), .A2(G953), .ZN(n735) );
  XNOR2_X1 U788 ( .A(n736), .B(n735), .ZN(n737) );
  XNOR2_X1 U789 ( .A(KEYINPUT122), .B(n737), .ZN(n738) );
  NAND2_X1 U790 ( .A1(n738), .A2(G898), .ZN(n739) );
  XOR2_X1 U791 ( .A(KEYINPUT124), .B(n739), .Z(n740) );
  NOR2_X1 U792 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U793 ( .A(n743), .B(n742), .ZN(G69) );
  XOR2_X1 U794 ( .A(n744), .B(n745), .Z(n749) );
  XNOR2_X1 U795 ( .A(n746), .B(n749), .ZN(n748) );
  NAND2_X1 U796 ( .A1(n748), .A2(n747), .ZN(n754) );
  XNOR2_X1 U797 ( .A(n749), .B(G227), .ZN(n750) );
  NAND2_X1 U798 ( .A1(n750), .A2(G900), .ZN(n751) );
  XOR2_X1 U799 ( .A(KEYINPUT125), .B(n751), .Z(n752) );
  NAND2_X1 U800 ( .A1(G953), .A2(n752), .ZN(n753) );
  NAND2_X1 U801 ( .A1(n754), .A2(n753), .ZN(G72) );
  XOR2_X1 U802 ( .A(G137), .B(KEYINPUT126), .Z(n755) );
  XNOR2_X1 U803 ( .A(n756), .B(n755), .ZN(G39) );
  XNOR2_X1 U804 ( .A(G134), .B(n757), .ZN(G36) );
  XOR2_X1 U805 ( .A(G125), .B(n758), .Z(n759) );
  XNOR2_X1 U806 ( .A(KEYINPUT37), .B(n759), .ZN(G27) );
  XNOR2_X1 U807 ( .A(G119), .B(n354), .ZN(G21) );
  XOR2_X1 U808 ( .A(G131), .B(n761), .Z(G33) );
endmodule

