//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 0 1 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 0 0 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n562, new_n563, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(G220));
  XOR2_X1   g012(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  AND2_X1   g017(.A1(G2072), .A2(G2078), .ZN(new_n443));
  NAND3_X1  g018(.A1(new_n443), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT66), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n466), .ZN(new_n468));
  OAI21_X1  g043(.A(KEYINPUT67), .B1(new_n468), .B2(new_n463), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n469), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n462), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n462), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n464), .A2(new_n466), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n462), .ZN(new_n477));
  INV_X1    g052(.A(G137), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n472), .A2(new_n479), .ZN(G160));
  NOR2_X1   g055(.A1(new_n468), .A2(new_n463), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(new_n462), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n481), .A2(G2105), .ZN(new_n483));
  AOI22_X1  g058(.A1(G124), .A2(new_n482), .B1(new_n483), .B2(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT68), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n484), .A2(new_n487), .ZN(G162));
  OAI211_X1 g063(.A(G126), .B(G2105), .C1(new_n468), .C2(new_n463), .ZN(new_n489));
  OR2_X1    g064(.A1(G102), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G114), .C2(new_n462), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g067(.A(G138), .B(new_n462), .C1(new_n468), .C2(new_n463), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR3_X1   g070(.A1(new_n495), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n467), .A2(new_n469), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n492), .B1(new_n494), .B2(new_n497), .ZN(G164));
  AND2_X1   g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NOR2_X1   g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  OAI21_X1  g075(.A(G62), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT70), .ZN(new_n502));
  NAND2_X1  g077(.A1(G75), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(new_n510), .A3(G62), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  OAI21_X1  g087(.A(G651), .B1(new_n504), .B2(new_n512), .ZN(new_n513));
  OR2_X1    g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n514), .A2(new_n515), .B1(new_n507), .B2(new_n508), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT69), .B(G88), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n506), .B1(new_n514), .B2(new_n515), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G50), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n513), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n501), .A2(KEYINPUT70), .B1(G75), .B2(G543), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n524), .B1(new_n525), .B2(new_n511), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n518), .A2(new_n520), .ZN(new_n527));
  OAI21_X1  g102(.A(KEYINPUT71), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n523), .A2(new_n528), .ZN(G166));
  AND2_X1   g104(.A1(KEYINPUT6), .A2(G651), .ZN(new_n530));
  NOR2_X1   g105(.A1(KEYINPUT6), .A2(G651), .ZN(new_n531));
  OAI21_X1  g106(.A(G543), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g109(.A(KEYINPUT72), .B(G543), .C1(new_n530), .C2(new_n531), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G51), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n516), .A2(G89), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n541));
  AND4_X1   g116(.A1(new_n537), .A2(new_n538), .A3(new_n540), .A4(new_n541), .ZN(G168));
  AOI22_X1  g117(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G90), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n500), .A2(new_n499), .B1(new_n530), .B2(new_n531), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n543), .A2(new_n524), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(G52), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n547), .B1(new_n534), .B2(new_n535), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n546), .A2(new_n548), .ZN(G171));
  NAND2_X1  g124(.A1(new_n514), .A2(new_n515), .ZN(new_n550));
  XNOR2_X1  g125(.A(KEYINPUT73), .B(G81), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n550), .A2(new_n509), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n554), .B1(new_n509), .B2(G56), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n552), .B1(new_n555), .B2(new_n524), .ZN(new_n556));
  INV_X1    g131(.A(G43), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n557), .B1(new_n534), .B2(new_n535), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n565), .B1(new_n507), .B2(new_n508), .ZN(new_n566));
  AND2_X1   g141(.A1(G78), .A2(G543), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n550), .A2(new_n509), .A3(G91), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n570), .B1(new_n519), .B2(G53), .ZN(new_n571));
  OAI211_X1 g146(.A(G53), .B(G543), .C1(new_n530), .C2(new_n531), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(KEYINPUT9), .ZN(new_n573));
  OAI211_X1 g148(.A(new_n568), .B(new_n569), .C1(new_n571), .C2(new_n573), .ZN(G299));
  INV_X1    g149(.A(G171), .ZN(G301));
  NAND4_X1  g150(.A1(new_n537), .A2(new_n538), .A3(new_n540), .A4(new_n541), .ZN(G286));
  INV_X1    g151(.A(G166), .ZN(G303));
  NAND2_X1  g152(.A1(new_n516), .A2(G87), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n519), .A2(G49), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n499), .A2(new_n500), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n585), .A2(G651), .B1(G48), .B2(new_n519), .ZN(new_n586));
  INV_X1    g161(.A(G86), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n545), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(KEYINPUT74), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT74), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n590), .B1(new_n545), .B2(new_n587), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n586), .A2(new_n589), .A3(new_n591), .ZN(G305));
  INV_X1    g167(.A(G60), .ZN(new_n593));
  INV_X1    g168(.A(G72), .ZN(new_n594));
  OAI22_X1  g169(.A1(new_n583), .A2(new_n593), .B1(new_n594), .B2(new_n506), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(KEYINPUT75), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT75), .ZN(new_n597));
  OAI221_X1 g172(.A(new_n597), .B1(new_n594), .B2(new_n506), .C1(new_n583), .C2(new_n593), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n596), .A2(G651), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n516), .A2(G85), .ZN(new_n600));
  XNOR2_X1  g175(.A(KEYINPUT76), .B(G47), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n536), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(G290));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n545), .B2(new_n605), .ZN(new_n606));
  NAND4_X1  g181(.A1(new_n550), .A2(new_n509), .A3(KEYINPUT10), .A4(G92), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g183(.A(KEYINPUT72), .B1(new_n550), .B2(G543), .ZN(new_n609));
  INV_X1    g184(.A(new_n535), .ZN(new_n610));
  OAI21_X1  g185(.A(G54), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n583), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G651), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n608), .A2(new_n611), .A3(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(new_n617), .B2(G171), .ZN(G284));
  OAI21_X1  g194(.A(new_n618), .B1(new_n617), .B2(G171), .ZN(G321));
  NAND2_X1  g195(.A1(G299), .A2(new_n617), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G168), .B2(new_n617), .ZN(G297));
  OAI21_X1  g197(.A(new_n621), .B1(G168), .B2(new_n617), .ZN(G280));
  AND3_X1   g198(.A1(new_n608), .A2(new_n611), .A3(new_n615), .ZN(new_n624));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G860), .ZN(G148));
  NOR2_X1   g201(.A1(new_n559), .A2(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n624), .A2(new_n625), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(G868), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT77), .Z(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n483), .A2(G135), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n482), .A2(G123), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n462), .A2(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT79), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT80), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2096), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n467), .A2(new_n469), .A3(new_n474), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT12), .Z(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT78), .B(KEYINPUT13), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2100), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n641), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n639), .A2(new_n644), .ZN(G156));
  XNOR2_X1  g220(.A(G2427), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2430), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(new_n650), .A3(KEYINPUT14), .ZN(new_n651));
  XOR2_X1   g226(.A(G1341), .B(G1348), .Z(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n651), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2451), .B(G2454), .Z(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n655), .A2(new_n658), .ZN(new_n660));
  AND3_X1   g235(.A1(new_n659), .A2(G14), .A3(new_n660), .ZN(G401));
  XOR2_X1   g236(.A(G2067), .B(G2678), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT82), .ZN(new_n663));
  NOR2_X1   g238(.A1(G2072), .A2(G2078), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n443), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2084), .B(G2090), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n663), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT18), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n663), .A2(new_n665), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n665), .B(KEYINPUT17), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n669), .B(new_n666), .C1(new_n663), .C2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n666), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n663), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n668), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2096), .B(G2100), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT83), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n674), .B(new_n676), .ZN(G227));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1956), .B(G2474), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1961), .B(G1966), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(new_n682), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n681), .A2(new_n682), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n686), .A2(KEYINPUT20), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(KEYINPUT20), .ZN(new_n688));
  OAI221_X1 g263(.A(new_n683), .B1(new_n680), .B2(new_n684), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G1991), .B(G1996), .Z(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n691), .A2(new_n693), .ZN(new_n696));
  AND3_X1   g271(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n695), .B1(new_n694), .B2(new_n696), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(G229));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G35), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G162), .B2(new_n700), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT29), .ZN(new_n703));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NOR2_X1   g279(.A1(G286), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT90), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G16), .B2(G21), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(KEYINPUT90), .B2(new_n705), .ZN(new_n709));
  INV_X1    g284(.A(G1966), .ZN(new_n710));
  OAI22_X1  g285(.A1(new_n703), .A2(G2090), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT31), .B(G11), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT30), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G28), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT91), .Z(new_n715));
  OAI21_X1  g290(.A(new_n700), .B1(new_n713), .B2(G28), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n712), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI22_X1  g292(.A1(new_n483), .A2(G141), .B1(G105), .B2(new_n474), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n482), .A2(G129), .ZN(new_n719));
  NAND3_X1  g294(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT26), .Z(new_n721));
  NAND3_X1  g296(.A1(new_n718), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n723), .A2(new_n700), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n700), .B2(G32), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT27), .B(G1996), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT89), .ZN(new_n727));
  OAI22_X1  g302(.A1(new_n725), .A2(new_n727), .B1(new_n700), .B2(new_n637), .ZN(new_n728));
  AOI211_X1 g303(.A(new_n717), .B(new_n728), .C1(new_n727), .C2(new_n725), .ZN(new_n729));
  NOR2_X1   g304(.A1(G27), .A2(G29), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G164), .B2(G29), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT94), .B(G2078), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT95), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n731), .B(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT24), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n700), .B1(new_n735), .B2(G34), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n735), .B2(G34), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G160), .B2(G29), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n738), .A2(G2084), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n709), .A2(new_n710), .ZN(new_n740));
  NAND4_X1  g315(.A1(new_n729), .A2(new_n734), .A3(new_n739), .A4(new_n740), .ZN(new_n741));
  AOI211_X1 g316(.A(new_n711), .B(new_n741), .C1(G2084), .C2(new_n738), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n703), .A2(G2090), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n704), .A2(G20), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT23), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n572), .B(new_n570), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n568), .A2(new_n569), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n745), .B1(new_n748), .B2(new_n704), .ZN(new_n749));
  INV_X1    g324(.A(G1956), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n743), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT96), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n704), .A2(G5), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G171), .B2(new_n704), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT92), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G1961), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT93), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n756), .A2(G1961), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n700), .A2(G26), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT28), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n483), .A2(G140), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n482), .A2(G128), .ZN(new_n763));
  OR2_X1    g338(.A1(G104), .A2(G2105), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n764), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n762), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n761), .B1(new_n767), .B2(new_n700), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT87), .B(G2067), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(G16), .A2(G19), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n559), .B2(G16), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G1341), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n772), .A2(G1341), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n770), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(G4), .A2(G16), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT86), .Z(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n616), .B2(new_n704), .ZN(new_n778));
  INV_X1    g353(.A(G1348), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(G29), .A2(G33), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT88), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT25), .Z(new_n784));
  INV_X1    g359(.A(G139), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n784), .B1(new_n477), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n467), .A2(new_n469), .A3(G127), .ZN(new_n787));
  NAND2_X1  g362(.A1(G115), .A2(G2104), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n462), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n782), .B1(new_n790), .B2(G29), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G2072), .ZN(new_n792));
  NOR4_X1   g367(.A1(new_n759), .A2(new_n775), .A3(new_n780), .A4(new_n792), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n742), .A2(new_n753), .A3(new_n758), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n704), .A2(G6), .ZN(new_n795));
  INV_X1    g370(.A(G305), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n795), .B1(new_n796), .B2(new_n704), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT32), .B(G1981), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n704), .A2(G23), .ZN(new_n800));
  AND3_X1   g375(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(new_n704), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT85), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT33), .B(G1976), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n799), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n704), .A2(G22), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G166), .B2(new_n704), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(G1971), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n803), .A2(new_n804), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n808), .A2(G1971), .ZN(new_n812));
  NOR4_X1   g387(.A1(new_n806), .A2(new_n810), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT34), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n814), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n700), .A2(G25), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n483), .A2(G131), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n482), .A2(G119), .ZN(new_n819));
  OR2_X1    g394(.A1(G95), .A2(G2105), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n820), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n818), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n817), .B1(new_n823), .B2(new_n700), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT35), .B(G1991), .Z(new_n825));
  XOR2_X1   g400(.A(new_n824), .B(new_n825), .Z(new_n826));
  AND2_X1   g401(.A1(new_n704), .A2(G24), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(G290), .B2(G16), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  AND2_X1   g404(.A1(new_n829), .A2(G1986), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n829), .A2(G1986), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n826), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n815), .A2(new_n816), .A3(new_n832), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT36), .Z(new_n834));
  NOR2_X1   g409(.A1(new_n794), .A2(new_n834), .ZN(G311));
  INV_X1    g410(.A(G311), .ZN(G150));
  OAI21_X1  g411(.A(G55), .B1(new_n609), .B2(new_n610), .ZN(new_n837));
  NAND2_X1  g412(.A1(G80), .A2(G543), .ZN(new_n838));
  INV_X1    g413(.A(G67), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n838), .B1(new_n583), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(G651), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n516), .A2(G93), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n837), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(G860), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT37), .Z(new_n845));
  NOR2_X1   g420(.A1(new_n616), .A2(new_n625), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT38), .Z(new_n847));
  INV_X1    g422(.A(KEYINPUT98), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(new_n559), .B2(KEYINPUT97), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT97), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(new_n556), .B2(new_n558), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(new_n843), .ZN(new_n852));
  INV_X1    g427(.A(G56), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n553), .B1(new_n583), .B2(new_n853), .ZN(new_n854));
  AOI22_X1  g429(.A1(new_n854), .A2(G651), .B1(new_n516), .B2(new_n551), .ZN(new_n855));
  OAI21_X1  g430(.A(G43), .B1(new_n609), .B2(new_n610), .ZN(new_n856));
  AND4_X1   g431(.A1(KEYINPUT97), .A2(new_n855), .A3(new_n856), .A4(new_n848), .ZN(new_n857));
  NOR3_X1   g432(.A1(new_n849), .A2(new_n852), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n855), .A2(new_n856), .A3(KEYINPUT97), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(KEYINPUT98), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n855), .A2(new_n856), .A3(KEYINPUT97), .A4(new_n848), .ZN(new_n861));
  AOI22_X1  g436(.A1(new_n860), .A2(new_n861), .B1(new_n843), .B2(new_n851), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n847), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n865), .A2(KEYINPUT39), .ZN(new_n866));
  INV_X1    g441(.A(G860), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(new_n865), .B2(KEYINPUT39), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n845), .B1(new_n866), .B2(new_n868), .ZN(G145));
  NAND2_X1  g444(.A1(new_n483), .A2(G142), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n482), .A2(G130), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n462), .A2(G118), .ZN(new_n872));
  OAI21_X1  g447(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n870), .B(new_n871), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n641), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n641), .A2(new_n874), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n723), .A2(new_n790), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n722), .B1(new_n789), .B2(new_n786), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n877), .A2(new_n880), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(G164), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n766), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n822), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n881), .A2(new_n886), .A3(new_n882), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n637), .A2(G160), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n637), .A2(G160), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n891), .A2(G162), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(G162), .B1(new_n891), .B2(new_n892), .ZN(new_n894));
  NOR3_X1   g469(.A1(new_n890), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n895), .A2(G37), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n890), .B1(new_n893), .B2(new_n894), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g474(.A(new_n863), .B(new_n628), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n616), .A2(new_n748), .ZN(new_n901));
  AOI21_X1  g476(.A(KEYINPUT99), .B1(new_n624), .B2(G299), .ZN(new_n902));
  AOI22_X1  g477(.A1(new_n606), .A2(new_n607), .B1(G651), .B2(new_n614), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n903), .A2(G299), .A3(KEYINPUT99), .A4(new_n611), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n901), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n900), .A2(new_n906), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n907), .A2(KEYINPUT100), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT99), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(new_n616), .B2(new_n748), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n904), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT41), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n912), .B1(new_n616), .B2(new_n748), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT101), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n906), .A2(new_n912), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT101), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n911), .A2(new_n917), .A3(new_n913), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n907), .B(KEYINPUT100), .C1(new_n900), .C2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(G166), .A2(new_n796), .ZN(new_n921));
  NAND2_X1  g496(.A1(G290), .A2(new_n801), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n599), .A2(G288), .A3(new_n600), .A4(new_n602), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n523), .A2(new_n528), .A3(G305), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n921), .A2(new_n922), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n922), .A2(new_n923), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n523), .A2(new_n528), .A3(G305), .ZN(new_n927));
  AOI21_X1  g502(.A(G305), .B1(new_n523), .B2(new_n528), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT42), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n925), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT102), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n933));
  AOI22_X1  g508(.A1(new_n921), .A2(new_n924), .B1(new_n922), .B2(new_n923), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n925), .A2(new_n929), .A3(KEYINPUT102), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n931), .B1(new_n938), .B2(new_n930), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n908), .A2(new_n920), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n939), .B1(new_n908), .B2(new_n920), .ZN(new_n941));
  OAI21_X1  g516(.A(G868), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n843), .A2(new_n617), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(G295));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n943), .ZN(G331));
  INV_X1    g520(.A(KEYINPUT104), .ZN(new_n946));
  INV_X1    g521(.A(new_n548), .ZN(new_n947));
  NAND2_X1  g522(.A1(G77), .A2(G543), .ZN(new_n948));
  INV_X1    g523(.A(G64), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n948), .B1(new_n583), .B2(new_n949), .ZN(new_n950));
  AOI22_X1  g525(.A1(new_n950), .A2(G651), .B1(new_n516), .B2(G90), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n946), .B1(new_n947), .B2(new_n951), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n546), .A2(new_n548), .A3(KEYINPUT104), .ZN(new_n953));
  OAI21_X1  g528(.A(G168), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n947), .A2(new_n951), .A3(new_n946), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT104), .B1(new_n546), .B2(new_n548), .ZN(new_n956));
  NAND3_X1  g531(.A1(G286), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n958), .B1(new_n858), .B2(new_n862), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n852), .B1(new_n849), .B2(new_n857), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n860), .A2(new_n843), .A3(new_n851), .A4(new_n861), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n960), .A2(new_n961), .A3(new_n954), .A4(new_n957), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT105), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AOI22_X1  g541(.A1(new_n910), .A2(new_n904), .B1(new_n748), .B2(new_n616), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n967), .B1(new_n959), .B2(new_n962), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n965), .B1(new_n963), .B2(new_n964), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n937), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G37), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n959), .A2(new_n962), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT105), .B1(new_n919), .B2(new_n974), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n975), .A2(new_n938), .A3(new_n969), .A4(new_n966), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n972), .A2(new_n973), .A3(new_n976), .ZN(new_n977));
  XOR2_X1   g552(.A(KEYINPUT103), .B(KEYINPUT43), .Z(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT106), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n970), .A2(new_n937), .A3(new_n971), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n914), .B1(new_n967), .B2(KEYINPUT41), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n983), .A2(new_n962), .A3(new_n959), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n937), .B1(new_n984), .B2(new_n968), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n985), .A2(new_n973), .A3(new_n978), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n981), .B1(new_n982), .B2(new_n986), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n985), .A2(new_n973), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n988), .A2(new_n976), .A3(KEYINPUT106), .A4(new_n978), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n980), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n975), .A2(new_n969), .A3(new_n966), .ZN(new_n991));
  AOI21_X1  g566(.A(G37), .B1(new_n991), .B2(new_n937), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n992), .A2(new_n976), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n988), .A2(new_n976), .ZN(new_n994));
  AOI22_X1  g569(.A1(new_n993), .A2(new_n978), .B1(KEYINPUT43), .B2(new_n994), .ZN(new_n995));
  MUX2_X1   g570(.A(new_n990), .B(new_n995), .S(KEYINPUT44), .Z(G397));
  INV_X1    g571(.A(G40), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n472), .A2(new_n997), .A3(new_n479), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n1000), .B1(G164), .B2(G1384), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1996), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n722), .B(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G2067), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n766), .B(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n823), .A2(new_n825), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n823), .A2(new_n825), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1004), .A2(new_n1006), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(G290), .B(G1986), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1002), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT63), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1013));
  OR2_X1    g588(.A1(G164), .A2(G1384), .ZN(new_n1014));
  XNOR2_X1  g589(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  OAI211_X1 g591(.A(KEYINPUT108), .B(new_n1013), .C1(new_n1014), .C2(new_n1016), .ZN(new_n1017));
  NOR4_X1   g592(.A1(G164), .A2(KEYINPUT108), .A3(G1384), .A4(new_n1016), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n998), .ZN(new_n1021));
  XNOR2_X1  g596(.A(KEYINPUT109), .B(G2090), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(G164), .A2(G1384), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT45), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1025), .A2(new_n1001), .A3(new_n998), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  OAI22_X1  g602(.A1(new_n1021), .A2(new_n1023), .B1(G1971), .B2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n523), .A2(new_n528), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1029));
  OR2_X1    g604(.A1(new_n1029), .A2(KEYINPUT110), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(KEYINPUT110), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n1032));
  INV_X1    g607(.A(G8), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1032), .B1(G166), .B2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1030), .A2(new_n1031), .A3(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1028), .A2(new_n1035), .A3(G8), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n585), .A2(G651), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n519), .A2(G48), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(G1981), .B1(new_n1039), .B2(new_n588), .ZN(new_n1040));
  XOR2_X1   g615(.A(KEYINPUT112), .B(G1981), .Z(new_n1041));
  NAND4_X1  g616(.A1(new_n586), .A2(new_n589), .A3(new_n591), .A4(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT113), .ZN(new_n1044));
  OR2_X1    g619(.A1(new_n1044), .A2(KEYINPUT49), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n998), .A2(new_n1024), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1047), .A2(new_n1033), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1044), .A2(KEYINPUT49), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1045), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n801), .A2(G1976), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1046), .A2(G8), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT111), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1046), .A2(KEYINPUT111), .A3(G8), .A4(new_n1051), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1054), .A2(KEYINPUT52), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G1976), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT52), .B1(G288), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1048), .A2(new_n1051), .A3(new_n1058), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1050), .A2(new_n1056), .A3(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1027), .A2(G1971), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1016), .B1(G164), .B2(G1384), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n998), .B(new_n1062), .C1(new_n1014), .C2(KEYINPUT50), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1063), .A2(new_n1023), .ZN(new_n1064));
  OAI21_X1  g639(.A(G8), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1035), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1036), .A2(new_n1060), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1026), .A2(new_n710), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n999), .A2(G2084), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT108), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1072), .B1(new_n1024), .B2(new_n1015), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1018), .B1(new_n1073), .B2(new_n1013), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1069), .B1(new_n1071), .B2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(G286), .A2(new_n1033), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1075), .A2(KEYINPUT116), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT116), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1012), .B1(new_n1068), .B2(new_n1080), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1074), .A2(new_n999), .A3(new_n1023), .ZN(new_n1082));
  OAI21_X1  g657(.A(G8), .B1(new_n1082), .B2(new_n1061), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT63), .B1(new_n1083), .B2(new_n1066), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1035), .B1(new_n1028), .B2(G8), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1050), .A2(new_n1056), .A3(new_n1059), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT114), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT114), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1050), .A2(new_n1056), .A3(new_n1089), .A4(new_n1059), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1086), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT117), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1085), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AOI211_X1 g668(.A(KEYINPUT117), .B(new_n1086), .C1(new_n1088), .C2(new_n1090), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1081), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1063), .A2(new_n750), .ZN(new_n1096));
  XOR2_X1   g671(.A(G299), .B(KEYINPUT57), .Z(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT56), .B(G2072), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1025), .A2(new_n1001), .A3(new_n998), .A4(new_n1098), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1096), .A2(new_n1097), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1027), .A2(new_n1098), .B1(new_n750), .B2(new_n1063), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT118), .B1(new_n1102), .B2(new_n1097), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1097), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1021), .A2(new_n779), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1047), .A2(new_n1005), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n616), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1101), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1103), .A2(KEYINPUT61), .A3(new_n1101), .A4(new_n1106), .ZN(new_n1112));
  XOR2_X1   g687(.A(KEYINPUT122), .B(KEYINPUT61), .Z(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1100), .B2(new_n1104), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n559), .A2(KEYINPUT121), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1025), .A2(new_n1003), .A3(new_n1001), .A4(new_n998), .ZN(new_n1116));
  OR2_X1    g691(.A1(new_n1116), .A2(KEYINPUT119), .ZN(new_n1117));
  XNOR2_X1  g692(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1118), .B(G1341), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1116), .A2(KEYINPUT119), .B1(new_n1046), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1115), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI211_X1 g698(.A(KEYINPUT59), .B(new_n1115), .C1(new_n1117), .C2(new_n1120), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1112), .B(new_n1114), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT60), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1108), .A2(KEYINPUT60), .A3(new_n1109), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n624), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1108), .A2(KEYINPUT60), .A3(new_n616), .A4(new_n1109), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1126), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1111), .B1(new_n1125), .B2(new_n1130), .ZN(new_n1131));
  OAI211_X1 g706(.A(G168), .B(new_n1069), .C1(new_n1071), .C2(new_n1074), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT51), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1132), .A2(new_n1133), .A3(G8), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1020), .A2(new_n1070), .B1(new_n710), .B2(new_n1026), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1033), .B1(new_n1135), .B2(G168), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1075), .A2(G286), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1134), .B1(new_n1138), .B2(KEYINPUT51), .ZN(new_n1139));
  XNOR2_X1  g714(.A(KEYINPUT123), .B(G1961), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1141), .B1(new_n1020), .B2(new_n998), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(G2078), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1025), .A2(new_n1144), .A3(new_n1001), .A4(new_n998), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(KEYINPUT53), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1143), .A2(new_n1146), .A3(G301), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT53), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1145), .B(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(G171), .B1(new_n1149), .B2(new_n1142), .ZN(new_n1150));
  AOI21_X1  g725(.A(KEYINPUT54), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n1139), .A2(new_n1068), .A3(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1147), .A2(new_n1150), .A3(KEYINPUT54), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT124), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT124), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1147), .A2(new_n1150), .A3(new_n1155), .A4(KEYINPUT54), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1131), .A2(new_n1152), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1036), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1045), .A2(new_n1049), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n801), .A2(new_n1057), .ZN(new_n1161));
  XOR2_X1   g736(.A(new_n1161), .B(KEYINPUT115), .Z(new_n1162));
  OAI21_X1  g737(.A(new_n1042), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1159), .B1(new_n1048), .B2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1095), .A2(new_n1158), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT62), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1139), .A2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1068), .A2(new_n1150), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1133), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1169));
  OAI21_X1  g744(.A(KEYINPUT62), .B1(new_n1169), .B2(new_n1134), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1167), .A2(new_n1168), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT125), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1167), .A2(new_n1168), .A3(KEYINPUT125), .A4(new_n1170), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1011), .B1(new_n1165), .B2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g751(.A1(G290), .A2(G1986), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1002), .A2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g753(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1181));
  AOI211_X1 g756(.A(new_n1180), .B(new_n1181), .C1(new_n1009), .C2(new_n1002), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1006), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1002), .B1(new_n1183), .B2(new_n722), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT46), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1185), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1186));
  NOR4_X1   g761(.A1(new_n999), .A2(new_n1001), .A3(KEYINPUT46), .A4(G1996), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1184), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  XOR2_X1   g763(.A(new_n1188), .B(KEYINPUT47), .Z(new_n1189));
  NAND2_X1  g764(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1190));
  OAI22_X1  g765(.A1(new_n1190), .A2(new_n1007), .B1(G2067), .B2(new_n766), .ZN(new_n1191));
  AOI211_X1 g766(.A(new_n1182), .B(new_n1189), .C1(new_n1002), .C2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1176), .A2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n1195));
  NOR3_X1   g769(.A1(G401), .A2(G227), .A3(new_n460), .ZN(new_n1196));
  OAI21_X1  g770(.A(new_n1196), .B1(new_n697), .B2(new_n698), .ZN(new_n1197));
  AOI21_X1  g771(.A(new_n1197), .B1(new_n896), .B2(new_n897), .ZN(new_n1198));
  NAND2_X1  g772(.A1(new_n987), .A2(new_n989), .ZN(new_n1199));
  AOI21_X1  g773(.A(new_n978), .B1(new_n992), .B2(new_n976), .ZN(new_n1200));
  OAI211_X1 g774(.A(new_n1195), .B(new_n1198), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1201));
  INV_X1    g775(.A(new_n1201), .ZN(new_n1202));
  AOI21_X1  g776(.A(new_n1195), .B1(new_n990), .B2(new_n1198), .ZN(new_n1203));
  NOR2_X1   g777(.A1(new_n1202), .A2(new_n1203), .ZN(G308));
  NAND2_X1  g778(.A1(new_n990), .A2(new_n1198), .ZN(G225));
endmodule


