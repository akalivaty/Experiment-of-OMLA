//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 0 1 1 0 0 1 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 0 1 1 0 1 1 0 0 0 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  INV_X1    g000(.A(G119), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G116), .ZN(new_n188));
  INV_X1    g002(.A(G116), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT2), .B(G113), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT66), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(G116), .B(G119), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT66), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT2), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G113), .ZN(new_n197));
  INV_X1    g011(.A(G113), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(KEYINPUT2), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n194), .B(new_n195), .C1(new_n197), .C2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n193), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n191), .A2(new_n192), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT64), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT64), .A2(G134), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(G137), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G137), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(KEYINPUT11), .A3(G134), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  AND2_X1   g026(.A1(KEYINPUT64), .A2(G134), .ZN(new_n213));
  NOR2_X1   g027(.A1(KEYINPUT64), .A2(G134), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n209), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT65), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT11), .ZN(new_n217));
  AND3_X1   g031(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n216), .B1(new_n215), .B2(new_n217), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n212), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G131), .ZN(new_n221));
  AOI21_X1  g035(.A(G137), .B1(new_n206), .B2(new_n207), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT65), .B1(new_n222), .B2(KEYINPUT11), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G131), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n226), .A3(new_n212), .ZN(new_n227));
  INV_X1    g041(.A(G146), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G143), .ZN(new_n229));
  INV_X1    g043(.A(G143), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G146), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n229), .A2(new_n231), .A3(KEYINPUT0), .A4(G128), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n229), .A2(new_n231), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT0), .B(G128), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n232), .B(new_n233), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n232), .B1(new_n234), .B2(new_n235), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT67), .ZN(new_n238));
  AOI22_X1  g052(.A1(new_n221), .A2(new_n227), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  AOI211_X1 g053(.A(G131), .B(new_n211), .C1(new_n223), .C2(new_n224), .ZN(new_n240));
  INV_X1    g054(.A(G128), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n229), .B(new_n231), .C1(KEYINPUT1), .C2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n229), .A2(new_n231), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT1), .B1(new_n230), .B2(G146), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n243), .A2(G128), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n205), .A2(G137), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n215), .A2(new_n246), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n242), .B(new_n245), .C1(new_n247), .C2(new_n226), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT30), .B1(new_n240), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n203), .B1(new_n239), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n237), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n226), .B1(new_n225), .B2(new_n212), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n251), .B1(new_n252), .B2(new_n240), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n245), .A2(new_n242), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n226), .B1(new_n215), .B2(new_n246), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n227), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(KEYINPUT30), .B1(new_n253), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT68), .B1(new_n250), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT30), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n237), .B1(new_n221), .B2(new_n227), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n211), .B1(new_n223), .B2(new_n224), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n248), .B1(new_n262), .B2(new_n226), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n203), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n238), .A2(new_n236), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n266), .B1(new_n252), .B2(new_n240), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n260), .B1(new_n227), .B2(new_n256), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n265), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT68), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n264), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n259), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n267), .A2(new_n257), .A3(new_n265), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(KEYINPUT69), .A2(G953), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(KEYINPUT69), .A2(G953), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G237), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n278), .A2(G210), .A3(new_n279), .ZN(new_n280));
  XOR2_X1   g094(.A(KEYINPUT26), .B(G101), .Z(new_n281));
  XNOR2_X1  g095(.A(new_n280), .B(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n282), .B(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n274), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n272), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n203), .B1(new_n261), .B2(new_n263), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT28), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n221), .A2(new_n227), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n263), .B1(new_n289), .B2(new_n266), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n288), .B1(new_n290), .B2(new_n265), .ZN(new_n291));
  NOR4_X1   g105(.A1(new_n239), .A2(new_n263), .A3(KEYINPUT28), .A4(new_n203), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n287), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n284), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT29), .B1(new_n286), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G902), .ZN(new_n296));
  OAI22_X1  g110(.A1(new_n291), .A2(new_n292), .B1(new_n265), .B2(new_n290), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n284), .A2(KEYINPUT29), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G472), .B1(new_n295), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n273), .A2(new_n284), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT71), .B(KEYINPUT31), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n264), .A2(new_n269), .A3(new_n270), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n270), .B1(new_n264), .B2(new_n269), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n302), .B(new_n303), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n284), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n293), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT31), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n301), .B1(new_n259), .B2(new_n271), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n306), .B(new_n308), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT32), .ZN(new_n312));
  NOR2_X1   g126(.A1(G472), .A2(G902), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n312), .B1(new_n311), .B2(new_n313), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n300), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT72), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI211_X1 g132(.A(KEYINPUT72), .B(new_n300), .C1(new_n314), .C2(new_n315), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n241), .A2(G119), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n187), .A2(G128), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT24), .B(G110), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT23), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n241), .A2(KEYINPUT23), .A3(G119), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n327), .A3(new_n321), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n324), .B1(G110), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G140), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT16), .B1(new_n330), .B2(G125), .ZN(new_n331));
  AND2_X1   g145(.A1(KEYINPUT74), .A2(G140), .ZN(new_n332));
  NOR2_X1   g146(.A1(KEYINPUT74), .A2(G140), .ZN(new_n333));
  OAI21_X1  g147(.A(G125), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT75), .ZN(new_n335));
  INV_X1    g149(.A(G125), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G140), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n338), .B(G125), .C1(new_n332), .C2(new_n333), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n335), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n331), .B1(new_n340), .B2(KEYINPUT16), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n341), .A2(new_n228), .ZN(new_n342));
  AOI211_X1 g156(.A(G146), .B(new_n331), .C1(new_n340), .C2(KEYINPUT16), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n329), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n322), .A2(new_n323), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT76), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n322), .A2(new_n323), .A3(KEYINPUT76), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n347), .B(new_n348), .C1(G110), .C2(new_n328), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n330), .A2(G125), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n337), .A2(new_n350), .A3(new_n228), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT16), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n339), .A2(new_n337), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n353), .B1(new_n354), .B2(new_n335), .ZN(new_n355));
  OAI21_X1  g169(.A(G146), .B1(new_n355), .B2(new_n331), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT77), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n352), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n357), .B1(new_n352), .B2(new_n356), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n344), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n278), .A2(G221), .A3(G234), .ZN(new_n361));
  XNOR2_X1  g175(.A(KEYINPUT22), .B(G137), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n361), .B(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n344), .B(new_n363), .C1(new_n358), .C2(new_n359), .ZN(new_n366));
  XOR2_X1   g180(.A(KEYINPUT73), .B(G217), .Z(new_n367));
  AOI21_X1  g181(.A(new_n367), .B1(G234), .B2(new_n296), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(G902), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n365), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n370), .B(KEYINPUT78), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n365), .A2(new_n366), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT25), .B1(new_n372), .B2(G902), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT25), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n365), .A2(new_n374), .A3(new_n296), .A4(new_n366), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n373), .A2(new_n375), .A3(new_n368), .ZN(new_n376));
  AND3_X1   g190(.A1(new_n371), .A2(new_n376), .A3(KEYINPUT79), .ZN(new_n377));
  AOI21_X1  g191(.A(KEYINPUT79), .B1(new_n371), .B2(new_n376), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n318), .A2(new_n319), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT80), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n318), .A2(new_n379), .A3(KEYINPUT80), .A4(new_n319), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT9), .B(G234), .ZN(new_n385));
  OAI21_X1  g199(.A(G221), .B1(new_n385), .B2(G902), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G104), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT3), .B1(new_n388), .B2(G107), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT3), .ZN(new_n390));
  INV_X1    g204(.A(G107), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n391), .A3(G104), .ZN(new_n392));
  INV_X1    g206(.A(G101), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n388), .A2(G107), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n389), .A2(new_n392), .A3(new_n393), .A4(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n388), .A2(G107), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n391), .A2(G104), .ZN(new_n397));
  OAI21_X1  g211(.A(G101), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT82), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n399), .A2(new_n400), .A3(new_n242), .A4(new_n245), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n395), .A2(new_n398), .ZN(new_n402));
  OAI21_X1  g216(.A(KEYINPUT82), .B1(new_n254), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n254), .A2(new_n402), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n401), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n289), .A2(new_n405), .ZN(new_n406));
  XOR2_X1   g220(.A(KEYINPUT83), .B(KEYINPUT12), .Z(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n252), .A2(new_n240), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT10), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n401), .A2(new_n410), .A3(new_n403), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n389), .A2(new_n392), .A3(new_n394), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT4), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(new_n413), .A3(G101), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(G101), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(KEYINPUT4), .A3(new_n395), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n266), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n399), .A2(KEYINPUT10), .A3(new_n242), .A4(new_n245), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n409), .A2(new_n411), .A3(new_n417), .A4(new_n418), .ZN(new_n419));
  NOR2_X1   g233(.A1(KEYINPUT83), .A2(KEYINPUT12), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n289), .A2(new_n405), .A3(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n408), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n278), .A2(G227), .ZN(new_n423));
  XOR2_X1   g237(.A(G110), .B(G140), .Z(new_n424));
  XOR2_X1   g238(.A(new_n423), .B(new_n424), .Z(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(KEYINPUT81), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n411), .A2(new_n417), .A3(new_n418), .ZN(new_n428));
  AOI21_X1  g242(.A(KEYINPUT84), .B1(new_n221), .B2(new_n227), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n428), .A2(new_n429), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(new_n432), .A3(new_n425), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n427), .A2(KEYINPUT85), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(KEYINPUT85), .B1(new_n433), .B2(new_n427), .ZN(new_n435));
  OAI21_X1  g249(.A(G469), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G469), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n437), .A2(new_n296), .ZN(new_n438));
  INV_X1    g252(.A(new_n425), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n428), .A2(new_n429), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n439), .B1(new_n440), .B2(new_n430), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n408), .A2(new_n419), .A3(new_n425), .A4(new_n421), .ZN(new_n442));
  AOI21_X1  g256(.A(G902), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n438), .B1(new_n443), .B2(new_n437), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n387), .B1(new_n436), .B2(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(G116), .B(G122), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n446), .B(new_n391), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n206), .A2(new_n207), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n230), .A2(G128), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n241), .A2(G143), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OR2_X1    g265(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT13), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n450), .B1(new_n449), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(KEYINPUT13), .B1(new_n230), .B2(G128), .ZN(new_n455));
  OR2_X1    g269(.A1(new_n455), .A2(KEYINPUT96), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(KEYINPUT96), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n454), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n447), .B(new_n452), .C1(new_n458), .C2(new_n205), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n451), .B(new_n448), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n446), .A2(new_n391), .ZN(new_n461));
  OR2_X1    g275(.A1(new_n461), .A2(KEYINPUT97), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(KEYINPUT97), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n189), .A2(KEYINPUT14), .A3(G122), .ZN(new_n464));
  INV_X1    g278(.A(new_n446), .ZN(new_n465));
  OAI211_X1 g279(.A(G107), .B(new_n464), .C1(new_n465), .C2(KEYINPUT14), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n460), .A2(new_n462), .A3(new_n463), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n459), .A2(new_n467), .ZN(new_n468));
  OR3_X1    g282(.A1(new_n367), .A2(G953), .A3(new_n385), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n468), .A2(new_n469), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n296), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(G478), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n473), .A2(KEYINPUT15), .ZN(new_n474));
  OR2_X1    g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n472), .A2(new_n474), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n475), .A2(KEYINPUT98), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(KEYINPUT98), .B1(new_n475), .B2(new_n476), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n341), .ZN(new_n481));
  XOR2_X1   g295(.A(KEYINPUT92), .B(G143), .Z(new_n482));
  NAND4_X1  g296(.A1(new_n482), .A2(new_n278), .A3(G214), .A4(new_n279), .ZN(new_n483));
  OR2_X1    g297(.A1(KEYINPUT69), .A2(G953), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n484), .A2(G214), .A3(new_n279), .A4(new_n275), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n485), .B1(KEYINPUT92), .B2(new_n230), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n226), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n483), .A2(new_n486), .A3(new_n226), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n481), .A2(G146), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n340), .A2(KEYINPUT19), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n337), .A2(new_n350), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n491), .B(new_n228), .C1(KEYINPUT19), .C2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n487), .A2(KEYINPUT18), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n340), .A2(G146), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n483), .A2(new_n486), .ZN(new_n496));
  NAND2_X1  g310(.A1(KEYINPUT18), .A2(G131), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n351), .A2(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AOI22_X1  g312(.A1(new_n490), .A2(new_n493), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(G113), .B(G122), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n500), .B(new_n388), .ZN(new_n501));
  OAI21_X1  g315(.A(KEYINPUT93), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(KEYINPUT94), .B1(new_n342), .B2(new_n343), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT17), .ZN(new_n504));
  AOI211_X1 g318(.A(new_n504), .B(new_n226), .C1(new_n483), .C2(new_n486), .ZN(new_n505));
  INV_X1    g319(.A(new_n489), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n506), .A2(new_n487), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n505), .B1(new_n507), .B2(new_n504), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n341), .A2(new_n228), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT94), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n356), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n503), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n498), .A2(new_n494), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n501), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n493), .ZN(new_n515));
  OAI22_X1  g329(.A1(new_n341), .A2(new_n228), .B1(new_n506), .B2(new_n487), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n513), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT93), .ZN(new_n518));
  INV_X1    g332(.A(new_n501), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n502), .A2(new_n514), .A3(new_n520), .ZN(new_n521));
  NOR2_X1   g335(.A1(G475), .A2(G902), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT20), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT20), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n521), .A2(new_n525), .A3(new_n522), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n512), .A2(new_n501), .A3(new_n513), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n501), .B1(new_n512), .B2(new_n513), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n296), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT95), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT95), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n532), .B(new_n296), .C1(new_n528), .C2(new_n529), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n531), .A2(G475), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G952), .ZN(new_n535));
  AOI211_X1 g349(.A(G953), .B(new_n535), .C1(G234), .C2(G237), .ZN(new_n536));
  AOI211_X1 g350(.A(new_n296), .B(new_n278), .C1(G234), .C2(G237), .ZN(new_n537));
  XOR2_X1   g351(.A(new_n537), .B(KEYINPUT99), .Z(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT21), .B(G898), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n480), .A2(new_n527), .A3(new_n534), .A4(new_n541), .ZN(new_n542));
  XOR2_X1   g356(.A(KEYINPUT89), .B(G224), .Z(new_n543));
  NOR2_X1   g357(.A1(new_n543), .A2(G953), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n544), .A2(KEYINPUT7), .ZN(new_n545));
  XOR2_X1   g359(.A(KEYINPUT0), .B(G128), .Z(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n243), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n336), .B1(new_n547), .B2(new_n232), .ZN(new_n548));
  AOI21_X1  g362(.A(G125), .B1(new_n245), .B2(new_n242), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n545), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT8), .ZN(new_n551));
  INV_X1    g365(.A(G122), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(G110), .ZN(new_n553));
  INV_X1    g367(.A(G110), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(G122), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT88), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n553), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n556), .B1(new_n553), .B2(new_n555), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n551), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n553), .A2(new_n555), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT88), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n553), .A2(new_n555), .A3(new_n556), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(KEYINPUT8), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n194), .A2(KEYINPUT5), .ZN(new_n564));
  OAI21_X1  g378(.A(G113), .B1(new_n188), .B2(KEYINPUT5), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  AOI22_X1  g380(.A1(new_n193), .A2(new_n200), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n559), .B(new_n563), .C1(new_n567), .C2(new_n402), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT87), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(new_n564), .A3(new_n569), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT5), .ZN(new_n571));
  OAI21_X1  g385(.A(KEYINPUT87), .B1(new_n571), .B2(new_n565), .ZN(new_n572));
  AND4_X1   g386(.A1(new_n201), .A2(new_n402), .A3(new_n570), .A4(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n550), .B1(new_n568), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n254), .A2(new_n336), .ZN(new_n575));
  INV_X1    g389(.A(new_n544), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n237), .A2(G125), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n544), .B1(new_n548), .B2(new_n549), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n545), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT90), .B1(new_n574), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n545), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n548), .A2(new_n549), .A3(new_n544), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n576), .B1(new_n575), .B2(new_n577), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT90), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n201), .A2(new_n402), .A3(new_n570), .A4(new_n572), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n559), .A2(new_n563), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n587), .B(new_n588), .C1(new_n402), .C2(new_n567), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n585), .A2(new_n586), .A3(new_n589), .A4(new_n550), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n416), .A2(new_n414), .ZN(new_n591));
  OAI21_X1  g405(.A(KEYINPUT86), .B1(new_n265), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n557), .A2(new_n558), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n201), .A2(new_n399), .A3(new_n570), .A4(new_n572), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT86), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n203), .A2(new_n596), .A3(new_n414), .A4(new_n416), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n592), .A2(new_n594), .A3(new_n595), .A4(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n581), .A2(new_n590), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n296), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(KEYINPUT91), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n592), .A2(new_n595), .A3(new_n597), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n593), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n603), .A2(KEYINPUT6), .A3(new_n598), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT6), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n602), .A2(new_n605), .A3(new_n593), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n578), .A2(new_n579), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n604), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT91), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n599), .A2(new_n609), .A3(new_n296), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n601), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(G210), .B1(G237), .B2(G902), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n601), .A2(new_n608), .A3(new_n612), .A4(new_n610), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(G214), .B1(G237), .B2(G902), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n542), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n384), .A2(new_n445), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G101), .ZN(G3));
  NAND2_X1  g436(.A1(new_n311), .A2(new_n296), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(G472), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n311), .A2(new_n313), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n445), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n628), .A2(new_n379), .ZN(new_n629));
  INV_X1    g443(.A(new_n615), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n619), .B1(new_n630), .B2(KEYINPUT100), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT100), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n614), .A2(new_n632), .A3(new_n615), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n527), .A2(new_n534), .ZN(new_n635));
  OAI21_X1  g449(.A(KEYINPUT101), .B1(new_n470), .B2(new_n471), .ZN(new_n636));
  XOR2_X1   g450(.A(new_n636), .B(KEYINPUT33), .Z(new_n637));
  NAND3_X1  g451(.A1(new_n637), .A2(G478), .A3(new_n296), .ZN(new_n638));
  INV_X1    g452(.A(new_n472), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n638), .B1(G478), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n635), .A2(new_n640), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n634), .A2(new_n641), .A3(new_n540), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n629), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT34), .B(G104), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G6));
  AND2_X1   g459(.A1(new_n527), .A2(new_n534), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n646), .A2(KEYINPUT102), .A3(new_n541), .A4(new_n479), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n631), .A2(new_n633), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n527), .A2(new_n534), .A3(new_n541), .A4(new_n479), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n647), .A2(new_n648), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n629), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT35), .B(G107), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  OR3_X1    g469(.A1(new_n360), .A2(KEYINPUT36), .A3(new_n364), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n360), .B1(KEYINPUT36), .B2(new_n364), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n656), .A2(new_n369), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n376), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n628), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n620), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT37), .B(G110), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G12));
  AND4_X1   g477(.A1(new_n445), .A2(new_n631), .A3(new_n633), .A4(new_n659), .ZN(new_n664));
  INV_X1    g478(.A(G900), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n536), .B1(new_n538), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n527), .A2(new_n534), .A3(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n668), .A2(new_n480), .ZN(new_n669));
  AND4_X1   g483(.A1(new_n318), .A2(new_n664), .A3(new_n319), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(new_n241), .ZN(G30));
  NAND2_X1  g485(.A1(new_n625), .A2(KEYINPUT32), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n307), .B1(new_n272), .B2(new_n273), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n285), .B1(new_n265), .B2(new_n290), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n296), .ZN(new_n677));
  OAI21_X1  g491(.A(G472), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n666), .B(KEYINPUT39), .Z(new_n681));
  NAND2_X1  g495(.A1(new_n445), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n682), .A2(KEYINPUT40), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n682), .A2(KEYINPUT40), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n680), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT38), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n616), .B(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n635), .A2(new_n479), .ZN(new_n688));
  NOR4_X1   g502(.A1(new_n687), .A2(new_n619), .A3(new_n659), .A4(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT103), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G143), .ZN(G45));
  AOI21_X1  g506(.A(KEYINPUT72), .B1(new_n674), .B2(new_n300), .ZN(new_n693));
  INV_X1    g507(.A(new_n319), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n641), .A2(new_n666), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n695), .A2(new_n696), .A3(new_n664), .A4(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n664), .A2(new_n318), .A3(new_n697), .A4(new_n319), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT104), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G146), .ZN(G48));
  OR2_X1    g516(.A1(new_n443), .A2(new_n437), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n443), .A2(new_n437), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n703), .A2(new_n386), .A3(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n695), .A2(new_n379), .A3(new_n642), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT41), .B(G113), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G15));
  NAND4_X1  g522(.A1(new_n318), .A2(new_n379), .A3(new_n319), .A4(new_n705), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n647), .A2(new_n648), .A3(new_n651), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(new_n189), .ZN(G18));
  INV_X1    g526(.A(new_n705), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n542), .A2(new_n713), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n631), .A2(new_n633), .A3(new_n659), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n318), .A2(new_n714), .A3(new_n715), .A4(new_n319), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  INV_X1    g531(.A(new_n313), .ZN(new_n718));
  INV_X1    g532(.A(new_n306), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n297), .A2(new_n307), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n720), .B1(new_n309), .B2(new_n310), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT105), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n719), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n720), .B(KEYINPUT105), .C1(new_n309), .C2(new_n310), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n718), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n624), .A2(KEYINPUT106), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT106), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n623), .A2(new_n727), .A3(G472), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n725), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n371), .A2(new_n376), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n688), .A2(new_n540), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n631), .A2(new_n705), .A3(new_n633), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n729), .A2(new_n730), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G122), .ZN(G24));
  NAND2_X1  g548(.A1(new_n723), .A2(new_n724), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n313), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n727), .B1(new_n623), .B2(G472), .ZN(new_n737));
  INV_X1    g551(.A(G472), .ZN(new_n738));
  AOI211_X1 g552(.A(KEYINPUT106), .B(new_n738), .C1(new_n311), .C2(new_n296), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n736), .B(new_n659), .C1(new_n737), .C2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT107), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n726), .A2(new_n728), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n743), .A2(KEYINPUT107), .A3(new_n659), .A4(new_n736), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n697), .A2(new_n732), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT108), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT108), .ZN(new_n749));
  AOI211_X1 g563(.A(new_n749), .B(new_n746), .C1(new_n742), .C2(new_n744), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(new_n336), .ZN(G27));
  AND2_X1   g566(.A1(new_n316), .A2(new_n730), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n427), .A2(KEYINPUT109), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT109), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n422), .A2(new_n755), .A3(new_n426), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n754), .A2(G469), .A3(new_n433), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n444), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT110), .B1(new_n758), .B2(new_n386), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n760));
  AOI211_X1 g574(.A(new_n760), .B(new_n387), .C1(new_n444), .C2(new_n757), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n614), .A2(new_n618), .A3(new_n615), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n759), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n753), .A2(KEYINPUT42), .A3(new_n697), .A4(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n318), .A2(new_n763), .A3(new_n319), .A4(new_n379), .ZN(new_n765));
  INV_X1    g579(.A(new_n697), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n764), .B1(new_n767), .B2(KEYINPUT42), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G131), .ZN(G33));
  INV_X1    g583(.A(new_n669), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n765), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G134), .ZN(G36));
  OR3_X1    g586(.A1(new_n434), .A2(new_n435), .A3(KEYINPUT45), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n754), .A2(KEYINPUT45), .A3(new_n433), .A4(new_n756), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(G469), .A3(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n438), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT46), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n777), .B1(new_n437), .B2(new_n443), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n775), .A2(KEYINPUT46), .A3(new_n776), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n387), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n780), .A2(new_n681), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n646), .A2(new_n640), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT43), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(new_n626), .A3(new_n659), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT44), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n762), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n781), .B(new_n787), .C1(new_n786), .C2(new_n785), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  INV_X1    g603(.A(KEYINPUT111), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n790), .A2(KEYINPUT47), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n790), .A2(KEYINPUT47), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n780), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR4_X1   g607(.A1(new_n695), .A2(new_n766), .A3(new_n379), .A4(new_n762), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n793), .B(new_n794), .C1(new_n780), .C2(new_n792), .ZN(new_n795));
  XOR2_X1   g609(.A(KEYINPUT112), .B(G140), .Z(new_n796));
  XNOR2_X1  g610(.A(new_n795), .B(new_n796), .ZN(G42));
  AOI21_X1  g611(.A(new_n670), .B1(new_n698), .B2(new_n700), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n634), .A2(new_n688), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n758), .A2(new_n386), .ZN(new_n800));
  XOR2_X1   g614(.A(new_n666), .B(KEYINPUT115), .Z(new_n801));
  NOR3_X1   g615(.A1(new_n800), .A2(new_n659), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n799), .A2(new_n679), .A3(new_n802), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n798), .B(new_n803), .C1(new_n748), .C2(new_n750), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT52), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT114), .ZN(new_n806));
  INV_X1    g620(.A(new_n641), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n648), .A2(new_n807), .A3(new_n541), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n733), .B(new_n716), .C1(new_n709), .C2(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n806), .B1(new_n809), .B2(new_n711), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n733), .A2(new_n716), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n652), .A2(new_n695), .A3(new_n379), .A4(new_n705), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n811), .A2(new_n812), .A3(new_n706), .A4(KEYINPUT114), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n803), .A2(new_n815), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n798), .B(new_n816), .C1(new_n748), .C2(new_n750), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n475), .A2(new_n476), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n445), .A2(new_n819), .A3(new_n659), .ZN(new_n820));
  OR3_X1    g634(.A1(new_n820), .A2(new_n668), .A3(new_n762), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n318), .A2(new_n319), .ZN(new_n822));
  OAI22_X1  g636(.A1(new_n765), .A2(new_n770), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n763), .A2(new_n697), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n824), .B1(new_n742), .B2(new_n744), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n641), .B1(new_n635), .B2(new_n819), .ZN(new_n827));
  AND4_X1   g641(.A1(new_n541), .A2(new_n827), .A3(new_n618), .A4(new_n616), .ZN(new_n828));
  AOI22_X1  g642(.A1(new_n828), .A2(new_n629), .B1(new_n660), .B2(new_n620), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n621), .A2(new_n826), .A3(new_n768), .A4(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n805), .A2(new_n814), .A3(new_n817), .A4(new_n830), .ZN(new_n831));
  XOR2_X1   g645(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n832));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n809), .A2(new_n711), .A3(new_n833), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n830), .A2(new_n817), .A3(new_n834), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n831), .A2(new_n832), .B1(new_n835), .B2(new_n805), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n831), .A2(new_n833), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n831), .A2(new_n832), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n838), .B1(new_n841), .B2(new_n837), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n713), .A2(new_n762), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n784), .A2(new_n536), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n753), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(KEYINPUT48), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n784), .A2(new_n536), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n729), .A2(new_n730), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n732), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n680), .A2(new_n379), .A3(new_n536), .A4(new_n843), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n851), .A2(new_n641), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n852), .A2(new_n535), .A3(G953), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n846), .A2(new_n850), .A3(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(KEYINPUT119), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n793), .B1(new_n780), .B2(new_n792), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n703), .A2(new_n704), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n856), .B1(new_n386), .B2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n859), .A2(new_n618), .A3(new_n617), .A4(new_n849), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n851), .A2(new_n635), .A3(new_n640), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n861), .B1(new_n844), .B2(new_n745), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT117), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n863), .B1(new_n713), .B2(new_n618), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n705), .A2(KEYINPUT117), .A3(new_n619), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n687), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n847), .A2(new_n848), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(KEYINPUT118), .A2(KEYINPUT50), .ZN(new_n868));
  AND2_X1   g682(.A1(KEYINPUT118), .A2(KEYINPUT50), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n870), .B1(new_n867), .B2(new_n868), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n860), .A2(KEYINPUT51), .A3(new_n862), .A4(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n860), .A2(new_n862), .A3(new_n871), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT51), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n855), .A2(new_n872), .A3(new_n875), .ZN(new_n876));
  OAI22_X1  g690(.A1(new_n842), .A2(new_n876), .B1(G952), .B2(G953), .ZN(new_n877));
  INV_X1    g691(.A(new_n782), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n878), .A2(new_n730), .A3(new_n386), .A4(new_n618), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n879), .A2(KEYINPUT113), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(KEYINPUT113), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n857), .B(KEYINPUT49), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n687), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n880), .A2(new_n680), .A3(new_n881), .A4(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n877), .A2(new_n884), .ZN(G75));
  NOR2_X1   g699(.A1(new_n278), .A2(G952), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(KEYINPUT122), .Z(new_n887));
  NAND3_X1  g701(.A1(new_n830), .A2(new_n814), .A3(new_n817), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n804), .A2(KEYINPUT52), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n832), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n805), .A2(new_n817), .A3(new_n830), .A4(new_n834), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n296), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT56), .B1(new_n892), .B2(G210), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n604), .A2(new_n606), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(new_n607), .ZN(new_n895));
  XNOR2_X1  g709(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n895), .B(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n887), .B1(new_n893), .B2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT56), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n892), .ZN(new_n902));
  INV_X1    g716(.A(G210), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT121), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT121), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n906), .B(new_n901), .C1(new_n902), .C2(new_n903), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n898), .B1(new_n905), .B2(new_n907), .ZN(G51));
  XNOR2_X1  g722(.A(new_n438), .B(KEYINPUT57), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n890), .A2(new_n891), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n910), .A2(KEYINPUT54), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n837), .B1(new_n890), .B2(new_n891), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n909), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n441), .A2(new_n442), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n902), .A2(new_n775), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n886), .B1(new_n915), .B2(new_n916), .ZN(G54));
  INV_X1    g731(.A(new_n521), .ZN(new_n918));
  NAND2_X1  g732(.A1(KEYINPUT58), .A2(G475), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n918), .B1(new_n902), .B2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n886), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n892), .A2(KEYINPUT58), .A3(G475), .A4(new_n521), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(G60));
  NAND2_X1  g737(.A1(G478), .A2(G902), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT59), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n637), .B1(new_n842), .B2(new_n925), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n637), .A2(new_n925), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n927), .B1(new_n911), .B2(new_n912), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n887), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n926), .A2(new_n929), .ZN(G63));
  NAND2_X1  g744(.A1(G217), .A2(G902), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT60), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n372), .B1(new_n836), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(KEYINPUT124), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT124), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n935), .B(new_n372), .C1(new_n836), .C2(new_n932), .ZN(new_n936));
  INV_X1    g750(.A(new_n887), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n932), .B1(new_n890), .B2(new_n891), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n656), .A2(new_n657), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT123), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n937), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n934), .A2(KEYINPUT61), .A3(new_n936), .A4(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n933), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT61), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n942), .A2(new_n945), .ZN(G66));
  NAND3_X1  g760(.A1(new_n814), .A2(new_n621), .A3(new_n829), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n278), .ZN(new_n948));
  OAI21_X1  g762(.A(G953), .B1(new_n543), .B2(new_n539), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n894), .B1(G898), .B2(new_n278), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT125), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n950), .B(new_n952), .ZN(G69));
  AOI21_X1  g767(.A(new_n258), .B1(new_n267), .B2(new_n268), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n491), .B1(KEYINPUT19), .B2(new_n492), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n954), .B(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n788), .A2(new_n795), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n682), .A2(new_n762), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n384), .A2(new_n827), .A3(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n798), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n751), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n691), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT62), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n961), .A2(KEYINPUT62), .A3(new_n691), .ZN(new_n965));
  AOI211_X1 g779(.A(new_n957), .B(new_n959), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n278), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n956), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n781), .A2(new_n753), .A3(new_n799), .ZN(new_n969));
  AND4_X1   g783(.A1(new_n788), .A2(new_n961), .A3(new_n795), .A4(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n768), .A2(new_n771), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT126), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n970), .A2(new_n278), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n956), .B1(G900), .B2(new_n967), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n278), .B1(G227), .B2(G900), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT127), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n968), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n977), .B1(new_n968), .B2(new_n975), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n978), .A2(new_n979), .ZN(G72));
  NAND2_X1  g794(.A1(new_n966), .A2(new_n675), .ZN(new_n981));
  INV_X1    g795(.A(new_n286), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n970), .A2(new_n982), .A3(new_n972), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n947), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n982), .A2(new_n675), .ZN(new_n985));
  NAND2_X1  g799(.A1(G472), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT63), .Z(new_n987));
  NAND2_X1  g801(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n841), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n921), .B1(new_n985), .B2(new_n987), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n984), .A2(new_n989), .A3(new_n990), .ZN(G57));
endmodule


