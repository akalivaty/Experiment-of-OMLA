//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1 0 0 0 1 0 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0 0 1 1 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT65), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  XNOR2_X1  g0008(.A(KEYINPUT68), .B(G244), .ZN(new_n209));
  XNOR2_X1  g0009(.A(KEYINPUT67), .B(G68), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G77), .A2(new_n209), .B1(new_n210), .B2(G238), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G97), .A2(G257), .ZN(new_n214));
  AND3_X1   g0014(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n211), .B(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G20), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT69), .Z(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT1), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n219), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  INV_X1    g0024(.A(KEYINPUT0), .ZN(new_n225));
  OR2_X1    g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(G50), .B1(G58), .B2(G68), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n228), .A2(G20), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n224), .A2(new_n225), .ZN(new_n232));
  NAND3_X1  g0032(.A1(new_n226), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT66), .Z(new_n234));
  NOR2_X1   g0034(.A1(new_n222), .A2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(new_n217), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT2), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n238), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G264), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n241), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT70), .ZN(new_n245));
  INV_X1    g0045(.A(G107), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G68), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(G58), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(new_n205), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  XNOR2_X1  g0053(.A(KEYINPUT3), .B(G33), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G223), .A3(G1698), .ZN(new_n255));
  INV_X1    g0055(.A(G1698), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n254), .A2(G222), .A3(new_n256), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n255), .B(new_n257), .C1(new_n205), .C2(new_n254), .ZN(new_n258));
  OR2_X1    g0058(.A1(new_n258), .A2(KEYINPUT71), .ZN(new_n259));
  AND2_X1   g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(new_n229), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n258), .A2(KEYINPUT71), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n259), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  INV_X1    g0064(.A(G45), .ZN(new_n265));
  AOI21_X1  g0065(.A(G1), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G274), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n261), .A2(new_n266), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n268), .B1(new_n269), .B2(G226), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n263), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G200), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n229), .B1(new_n219), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G20), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT8), .B(G58), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT72), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT72), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(new_n216), .A3(KEYINPUT8), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT73), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n281), .B1(new_n273), .B2(G20), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n275), .A2(KEYINPUT73), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI22_X1  g0084(.A1(new_n204), .A2(new_n275), .B1(new_n280), .B2(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G20), .A2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G150), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n274), .B1(new_n285), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G1), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(G13), .A3(G20), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT74), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n291), .A2(KEYINPUT74), .A3(G13), .A4(G20), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n202), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(new_n274), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n275), .A2(G1), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n298), .A2(G50), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n290), .A2(new_n297), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT9), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n272), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT10), .ZN(new_n306));
  INV_X1    g0106(.A(new_n302), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT9), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n263), .A2(G190), .A3(new_n270), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n305), .A2(new_n306), .A3(new_n308), .A4(new_n309), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n308), .A2(new_n309), .A3(new_n272), .A4(new_n304), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT10), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G179), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n263), .A2(new_n314), .A3(new_n270), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT75), .ZN(new_n316));
  OR2_X1    g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n315), .A2(new_n316), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n307), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G169), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n271), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n313), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n294), .A2(new_n295), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT76), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n274), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n294), .A2(KEYINPUT76), .A3(new_n295), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n327), .A2(new_n300), .A3(new_n328), .A4(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(new_n205), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G20), .A2(G77), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT15), .B(G87), .ZN(new_n333));
  OAI221_X1 g0133(.A(new_n332), .B1(new_n276), .B2(new_n287), .C1(new_n284), .C2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n331), .B1(new_n274), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n327), .A2(new_n329), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n335), .B1(G77), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n254), .A2(G238), .A3(G1698), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(new_n246), .B2(new_n254), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n273), .A2(KEYINPUT3), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT3), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G33), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NOR3_X1   g0145(.A1(new_n345), .A2(new_n217), .A3(G1698), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n261), .B1(new_n341), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n269), .A2(new_n209), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n347), .A2(new_n267), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G200), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n339), .A2(KEYINPUT77), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G190), .ZN(new_n352));
  OR2_X1    g0152(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT77), .ZN(new_n354));
  INV_X1    g0154(.A(new_n350), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n354), .B1(new_n338), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n351), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n254), .A2(G226), .A3(new_n256), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n254), .A2(G232), .A3(G1698), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G33), .A2(G97), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n261), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n269), .A2(G238), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(new_n267), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT13), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n362), .A2(KEYINPUT13), .A3(new_n267), .A4(new_n363), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(G169), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT14), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n364), .A2(KEYINPUT79), .A3(KEYINPUT13), .ZN(new_n370));
  NAND2_X1  g0170(.A1(KEYINPUT79), .A2(KEYINPUT13), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n362), .A2(new_n371), .A3(new_n267), .A4(new_n363), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n370), .A2(G179), .A3(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT14), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n366), .A2(new_n374), .A3(G169), .A4(new_n367), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n369), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  OAI22_X1  g0176(.A1(new_n284), .A2(new_n205), .B1(new_n210), .B2(new_n275), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT80), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n286), .A2(G50), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT80), .ZN(new_n380));
  OAI221_X1 g0180(.A(new_n380), .B1(new_n210), .B2(new_n275), .C1(new_n284), .C2(new_n205), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n378), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n274), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT11), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT11), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n382), .A2(new_n385), .A3(new_n274), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT12), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n325), .A2(new_n388), .ZN(new_n389));
  NOR3_X1   g0189(.A1(new_n337), .A2(new_n388), .A3(new_n210), .ZN(new_n390));
  INV_X1    g0190(.A(G68), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n391), .B1(new_n330), .B2(KEYINPUT12), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n387), .A2(new_n389), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n376), .A2(new_n394), .ZN(new_n395));
  AND2_X1   g0195(.A1(new_n387), .A2(new_n393), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n370), .A2(G190), .A3(new_n372), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n366), .A2(G200), .A3(new_n367), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n396), .A2(new_n397), .A3(new_n389), .A4(new_n398), .ZN(new_n399));
  AND3_X1   g0199(.A1(new_n357), .A2(new_n395), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n254), .A2(G226), .A3(G1698), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n254), .A2(G223), .A3(new_n256), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G33), .A2(G87), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n268), .B1(new_n404), .B2(new_n261), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n269), .A2(G232), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n320), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n404), .A2(new_n261), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n409), .A2(new_n314), .A3(new_n267), .A4(new_n406), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT83), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT83), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n405), .A2(new_n412), .A3(new_n314), .A4(new_n406), .ZN(new_n413));
  AND3_X1   g0213(.A1(new_n408), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  XNOR2_X1  g0214(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n210), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT82), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n273), .B2(KEYINPUT3), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n343), .A2(KEYINPUT82), .A3(G33), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(new_n342), .A3(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n421), .A2(KEYINPUT7), .A3(new_n275), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT7), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(new_n254), .B2(G20), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n417), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n201), .B1(new_n210), .B2(G58), .ZN(new_n426));
  INV_X1    g0226(.A(G159), .ZN(new_n427));
  OAI22_X1  g0227(.A1(new_n426), .A2(new_n275), .B1(new_n427), .B2(new_n287), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n416), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n345), .A2(KEYINPUT7), .A3(new_n275), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n391), .B1(new_n424), .B2(new_n430), .ZN(new_n431));
  OR2_X1    g0231(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT16), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n274), .B(new_n429), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n280), .A2(new_n299), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n435), .A2(new_n298), .B1(new_n296), .B2(new_n280), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n414), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT18), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n414), .A2(KEYINPUT18), .A3(new_n437), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n407), .A2(G200), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n405), .A2(G190), .A3(new_n406), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n434), .A2(new_n436), .A3(new_n443), .A4(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT17), .ZN(new_n446));
  INV_X1    g0246(.A(new_n436), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n428), .A2(new_n431), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n328), .B1(new_n448), .B2(KEYINPUT16), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n447), .B1(new_n449), .B2(new_n429), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT17), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n450), .A2(new_n451), .A3(new_n443), .A4(new_n444), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n446), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n442), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n349), .A2(G179), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n456), .B(KEYINPUT78), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n349), .A2(new_n320), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n457), .A2(new_n338), .A3(new_n458), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n324), .A2(new_n400), .A3(new_n455), .A4(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT21), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G283), .ZN(new_n462));
  INV_X1    g0262(.A(G97), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n462), .B(new_n275), .C1(G33), .C2(new_n463), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n464), .B(new_n274), .C1(new_n275), .C2(G116), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT20), .ZN(new_n466));
  XNOR2_X1  g0266(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n336), .A2(new_n248), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n327), .A2(G116), .A3(new_n328), .A4(new_n329), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n291), .A2(G33), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(KEYINPUT87), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  AND3_X1   g0273(.A1(new_n294), .A2(KEYINPUT76), .A3(new_n295), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT76), .B1(new_n294), .B2(new_n295), .ZN(new_n475));
  NOR3_X1   g0275(.A1(new_n474), .A2(new_n475), .A3(new_n274), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT87), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n476), .A2(new_n477), .A3(G116), .A4(new_n471), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n469), .B1(new_n473), .B2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n342), .A2(new_n344), .A3(G257), .A4(new_n256), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n342), .A2(new_n344), .A3(G264), .A4(G1698), .ZN(new_n481));
  INV_X1    g0281(.A(G303), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n480), .B(new_n481), .C1(new_n482), .C2(new_n254), .ZN(new_n483));
  XNOR2_X1  g0283(.A(KEYINPUT5), .B(G41), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n291), .A2(G45), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n261), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n483), .A2(new_n261), .B1(new_n487), .B2(G270), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n484), .A2(G274), .A3(new_n486), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G169), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n461), .B1(new_n479), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n478), .A2(new_n473), .ZN(new_n493));
  INV_X1    g0293(.A(new_n469), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n491), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(KEYINPUT21), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n483), .A2(new_n261), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n487), .A2(G270), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n498), .A2(G179), .A3(new_n489), .A4(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n490), .A2(G200), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n488), .A2(G190), .A3(new_n489), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n479), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n492), .A2(new_n497), .A3(new_n502), .A4(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n342), .A2(new_n344), .A3(G244), .A4(new_n256), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT4), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n254), .A2(KEYINPUT4), .A3(G244), .A4(new_n256), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n254), .A2(G250), .A3(G1698), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n509), .A2(new_n510), .A3(new_n462), .A4(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n261), .ZN(new_n513));
  INV_X1    g0313(.A(new_n489), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n514), .B1(G257), .B2(new_n487), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n320), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n246), .B1(new_n422), .B2(new_n424), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT6), .ZN(new_n519));
  NOR3_X1   g0319(.A1(new_n519), .A2(new_n463), .A3(G107), .ZN(new_n520));
  XNOR2_X1  g0320(.A(G97), .B(G107), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n520), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  OAI22_X1  g0322(.A1(new_n522), .A2(new_n275), .B1(new_n205), .B2(new_n287), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n274), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n325), .A2(G97), .ZN(new_n525));
  NOR3_X1   g0325(.A1(new_n296), .A2(new_n274), .A3(new_n472), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n525), .B1(new_n526), .B2(G97), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n484), .A2(new_n486), .ZN(new_n529));
  INV_X1    g0329(.A(new_n261), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n529), .A2(new_n530), .A3(G257), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n489), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(new_n261), .B2(new_n512), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n314), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n517), .A2(new_n528), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n513), .A2(G190), .A3(new_n515), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(KEYINPUT84), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT84), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n533), .A2(new_n538), .A3(G190), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(G200), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n524), .B(new_n527), .C1(new_n533), .C2(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n535), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n342), .A2(new_n344), .A3(G238), .A4(new_n256), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n342), .A2(new_n344), .A3(G244), .A4(G1698), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G116), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n261), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n486), .A2(G274), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n485), .B(G250), .C1(new_n260), .C2(new_n229), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(G200), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n282), .A2(G97), .A3(new_n283), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT19), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n342), .A2(new_n344), .A3(new_n275), .A4(G68), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n275), .B1(new_n360), .B2(new_n557), .ZN(new_n560));
  INV_X1    g0360(.A(G87), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n561), .A2(new_n463), .A3(new_n246), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n558), .A2(new_n559), .A3(new_n563), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n336), .A2(new_n333), .B1(new_n564), .B2(new_n274), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT85), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n325), .A2(new_n328), .A3(G87), .A4(new_n471), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n555), .A2(new_n565), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n556), .A2(new_n557), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n563), .A2(new_n559), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n274), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n333), .B1(new_n474), .B2(new_n475), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(new_n567), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n552), .B1(new_n548), .B2(new_n261), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n574), .A2(new_n541), .ZN(new_n575));
  OAI21_X1  g0375(.A(KEYINPUT85), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n549), .A2(new_n553), .A3(G190), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT86), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n574), .A2(KEYINPUT86), .A3(G190), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n568), .A2(new_n576), .A3(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n526), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n565), .B1(new_n333), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n554), .A2(new_n320), .ZN(new_n585));
  AOI211_X1 g0385(.A(G179), .B(new_n552), .C1(new_n261), .C2(new_n548), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n584), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n582), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n342), .A2(new_n344), .A3(G257), .A4(G1698), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n342), .A2(new_n344), .A3(G250), .A4(new_n256), .ZN(new_n591));
  NAND2_X1  g0391(.A1(G33), .A2(G294), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n261), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n487), .A2(G264), .ZN(new_n595));
  AOI21_X1  g0395(.A(KEYINPUT88), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n594), .A2(new_n595), .A3(KEYINPUT88), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n514), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n594), .A2(new_n595), .A3(new_n489), .ZN(new_n600));
  OAI22_X1  g0400(.A1(new_n599), .A2(G200), .B1(G190), .B2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n342), .A2(new_n344), .A3(new_n275), .A4(G87), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT22), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT22), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n254), .A2(new_n604), .A3(new_n275), .A4(G87), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n275), .A2(G33), .A3(G116), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n246), .A2(G20), .ZN(new_n608));
  XNOR2_X1  g0408(.A(new_n608), .B(KEYINPUT23), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n606), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT24), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n609), .B1(new_n603), .B2(new_n605), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT24), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(new_n614), .A3(new_n607), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n328), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n583), .A2(new_n246), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n296), .A2(new_n246), .ZN(new_n618));
  XNOR2_X1  g0418(.A(new_n618), .B(KEYINPUT25), .ZN(new_n619));
  NOR3_X1   g0419(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n601), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n612), .A2(new_n615), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n274), .ZN(new_n623));
  INV_X1    g0423(.A(new_n617), .ZN(new_n624));
  INV_X1    g0424(.A(new_n619), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n594), .A2(KEYINPUT88), .A3(new_n595), .ZN(new_n627));
  OAI211_X1 g0427(.A(G179), .B(new_n489), .C1(new_n627), .C2(new_n596), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n600), .A2(G169), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n544), .A2(new_n589), .A3(new_n621), .A4(new_n631), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n460), .A2(new_n506), .A3(new_n632), .ZN(G372));
  NAND2_X1  g0433(.A1(new_n440), .A2(new_n441), .ZN(new_n634));
  INV_X1    g0434(.A(new_n459), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n635), .A2(new_n399), .B1(new_n394), .B2(new_n376), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n634), .B1(new_n636), .B2(new_n454), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n637), .A2(new_n313), .B1(new_n321), .B2(new_n319), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n517), .A2(new_n528), .A3(new_n534), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n639), .A2(new_n582), .A3(new_n588), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(KEYINPUT26), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT90), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT89), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n548), .A2(new_n643), .A3(new_n261), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n643), .B1(new_n548), .B2(new_n261), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n553), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n320), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n642), .B1(new_n647), .B2(new_n587), .ZN(new_n648));
  AOI211_X1 g0448(.A(KEYINPUT90), .B(new_n586), .C1(new_n646), .C2(new_n320), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n584), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n641), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT26), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n646), .A2(G200), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n653), .A2(new_n577), .A3(new_n567), .A4(new_n565), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n650), .A2(new_n652), .A3(new_n654), .A4(new_n639), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n492), .A2(new_n497), .A3(new_n502), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n617), .B1(new_n622), .B2(new_n274), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n657), .A2(new_n625), .B1(new_n629), .B2(new_n628), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n544), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n650), .A2(new_n621), .A3(new_n654), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n651), .B(new_n655), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n638), .B1(new_n460), .B2(new_n662), .ZN(G369));
  INV_X1    g0463(.A(G13), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(G20), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n291), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G213), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(G343), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n479), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n656), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n506), .B2(new_n673), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G330), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n600), .A2(G190), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n489), .B1(new_n627), .B2(new_n596), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n678), .B1(new_n679), .B2(new_n541), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n626), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(new_n658), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n620), .B2(new_n672), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n631), .B2(new_n672), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n677), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n656), .A2(new_n672), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n682), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n658), .A2(new_n672), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n685), .A2(new_n690), .ZN(G399));
  INV_X1    g0491(.A(new_n223), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n562), .A2(G116), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G1), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n227), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT95), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT29), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n640), .A2(new_n652), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT93), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n650), .A2(KEYINPUT26), .A3(new_n654), .A4(new_n639), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT93), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n640), .A2(new_n704), .A3(new_n652), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n650), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(KEYINPUT94), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n659), .A2(new_n660), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT94), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n706), .A2(new_n710), .A3(new_n650), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n708), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n700), .B1(new_n712), .B2(new_n672), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n661), .A2(new_n672), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(KEYINPUT29), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n500), .A2(KEYINPUT91), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT91), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n488), .A2(new_n718), .A3(G179), .A4(new_n489), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n597), .A2(new_n598), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n513), .A2(new_n574), .A3(new_n515), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n720), .A2(KEYINPUT30), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n721), .A2(new_n722), .A3(new_n717), .A4(new_n719), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT30), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n646), .A2(new_n314), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n727), .A2(new_n490), .A3(new_n679), .A4(new_n516), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n723), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n671), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n730), .A2(KEYINPUT31), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(KEYINPUT31), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n632), .A2(new_n506), .ZN(new_n734));
  AOI21_X1  g0534(.A(KEYINPUT92), .B1(new_n734), .B2(new_n672), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT92), .ZN(new_n736));
  NOR4_X1   g0536(.A1(new_n632), .A2(new_n736), .A3(new_n506), .A4(new_n671), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n733), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G330), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n699), .B1(new_n716), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n716), .A2(new_n699), .A3(new_n739), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n698), .B1(new_n743), .B2(G1), .ZN(G364));
  AOI21_X1  g0544(.A(new_n291), .B1(new_n665), .B2(G45), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n693), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n692), .A2(new_n254), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n228), .A2(new_n265), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n749), .B(new_n750), .C1(new_n252), .C2(new_n265), .ZN(new_n751));
  INV_X1    g0551(.A(G355), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n254), .A2(new_n223), .ZN(new_n753));
  OAI221_X1 g0553(.A(new_n751), .B1(G116), .B2(new_n223), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G13), .A2(G33), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G20), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n229), .B1(G20), .B2(new_n320), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n748), .B1(new_n754), .B2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n757), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n760), .B1(new_n675), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n275), .A2(G179), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G190), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n254), .B1(new_n766), .B2(G329), .ZN(new_n767));
  INV_X1    g0567(.A(G294), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n352), .A2(G179), .A3(G200), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n275), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n767), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n352), .A2(new_n541), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n275), .A2(new_n314), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(KEYINPUT97), .B(G326), .Z(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n773), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n778), .A2(new_n352), .A3(G200), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G322), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n777), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n778), .A2(new_n541), .A3(G190), .ZN(new_n783));
  XNOR2_X1  g0583(.A(KEYINPUT33), .B(G317), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G311), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n773), .A2(new_n764), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n785), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n763), .A2(new_n352), .A3(G200), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT96), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n771), .B(new_n788), .C1(G283), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n772), .A2(new_n763), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n795), .B1(new_n482), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n770), .A2(new_n463), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n796), .A2(new_n561), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n799), .B1(G50), .B2(new_n775), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(new_n205), .B2(new_n787), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n798), .B(new_n801), .C1(G68), .C2(new_n783), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n345), .B1(new_n779), .B2(G58), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n802), .B(new_n803), .C1(new_n246), .C2(new_n793), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n766), .A2(G159), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT32), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n797), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT98), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n762), .B1(new_n808), .B2(new_n758), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT99), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n677), .A2(new_n747), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(G330), .B2(new_n675), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n810), .A2(new_n812), .ZN(G396));
  OAI22_X1  g0613(.A1(new_n246), .A2(new_n796), .B1(new_n787), .B2(new_n248), .ZN(new_n814));
  INV_X1    g0614(.A(new_n783), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n815), .A2(KEYINPUT100), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(KEYINPUT100), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n814), .B1(new_n819), .B2(G283), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n775), .A2(G303), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n794), .A2(G87), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n345), .B1(new_n780), .B2(new_n768), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n798), .B(new_n823), .C1(G311), .C2(new_n766), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n820), .A2(new_n821), .A3(new_n822), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n794), .A2(G68), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n254), .B1(new_n770), .B2(new_n216), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(G132), .B2(new_n766), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n826), .B(new_n828), .C1(new_n202), .C2(new_n796), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT101), .ZN(new_n830));
  INV_X1    g0630(.A(new_n787), .ZN(new_n831));
  AOI22_X1  g0631(.A1(G137), .A2(new_n775), .B1(new_n831), .B2(G159), .ZN(new_n832));
  INV_X1    g0632(.A(G143), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n832), .B1(new_n780), .B2(new_n833), .C1(new_n288), .C2(new_n815), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT34), .Z(new_n835));
  OAI21_X1  g0635(.A(new_n825), .B1(new_n830), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n758), .A2(new_n755), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n836), .A2(new_n758), .B1(new_n205), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n459), .A2(new_n671), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n338), .A2(new_n671), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n357), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n839), .B1(new_n841), .B2(new_n459), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n747), .B(new_n838), .C1(new_n842), .C2(new_n756), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n841), .A2(new_n459), .ZN(new_n844));
  INV_X1    g0644(.A(new_n839), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n714), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n842), .A2(new_n661), .A3(new_n672), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(new_n739), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n843), .B1(new_n850), .B2(new_n747), .ZN(G384));
  INV_X1    g0651(.A(KEYINPUT105), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n408), .A2(new_n411), .A3(new_n413), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n450), .B1(new_n853), .B2(new_n669), .ZN(new_n854));
  INV_X1    g0654(.A(new_n445), .ZN(new_n855));
  OAI21_X1  g0655(.A(KEYINPUT37), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT37), .ZN(new_n857));
  INV_X1    g0657(.A(new_n669), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n437), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n438), .A2(new_n857), .A3(new_n859), .A4(new_n445), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n453), .A2(KEYINPUT104), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT104), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n446), .A2(new_n863), .A3(new_n452), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n862), .A2(new_n634), .A3(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n859), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n861), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n852), .B1(new_n867), .B2(KEYINPUT38), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT38), .ZN(new_n869));
  AOI22_X1  g0669(.A1(KEYINPUT104), .A2(new_n453), .B1(new_n440), .B2(new_n441), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n859), .B1(new_n870), .B2(new_n864), .ZN(new_n871));
  OAI211_X1 g0671(.A(KEYINPUT105), .B(new_n869), .C1(new_n871), .C2(new_n861), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT39), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT103), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n432), .A2(new_n416), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n447), .B1(new_n449), .B2(new_n875), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n445), .B(new_n874), .C1(new_n853), .C2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n876), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n858), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n878), .A2(new_n414), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n874), .B1(new_n881), .B2(new_n445), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT37), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n860), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n879), .B1(new_n634), .B2(new_n453), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n884), .A2(new_n886), .A3(KEYINPUT38), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n868), .A2(new_n872), .A3(new_n873), .A4(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n860), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n876), .A2(new_n853), .ZN(new_n890));
  OAI21_X1  g0690(.A(KEYINPUT103), .B1(new_n890), .B2(new_n855), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n891), .A2(new_n879), .A3(new_n877), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n889), .B1(new_n892), .B2(KEYINPUT37), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n869), .B1(new_n893), .B2(new_n885), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n887), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT39), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n888), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n395), .A2(new_n671), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n395), .A2(new_n672), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n394), .A2(new_n671), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n395), .A2(new_n399), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT102), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT102), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n395), .A2(new_n399), .A3(new_n904), .A4(new_n901), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n900), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(new_n848), .B2(new_n845), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n895), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n442), .A2(new_n669), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n899), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n460), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n713), .B2(new_n715), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n638), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n910), .B(new_n913), .Z(new_n914));
  NOR3_X1   g0714(.A1(new_n681), .A2(new_n658), .A3(new_n543), .ZN(new_n915));
  AND4_X1   g0715(.A1(new_n492), .A2(new_n497), .A3(new_n502), .A4(new_n505), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n915), .A2(new_n916), .A3(new_n589), .A4(new_n672), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n736), .ZN(new_n918));
  INV_X1    g0718(.A(new_n632), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n919), .A2(KEYINPUT92), .A3(new_n916), .A4(new_n672), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n846), .B1(new_n921), .B2(new_n733), .ZN(new_n922));
  INV_X1    g0722(.A(new_n906), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n922), .A2(new_n895), .A3(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT40), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n868), .A2(new_n872), .A3(new_n887), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n927), .A2(KEYINPUT40), .A3(new_n923), .A4(new_n922), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n918), .A2(new_n920), .B1(new_n732), .B2(new_n731), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n460), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n929), .B(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(G330), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n914), .B(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n291), .B2(new_n665), .ZN(new_n935));
  INV_X1    g0735(.A(new_n522), .ZN(new_n936));
  OAI211_X1 g0736(.A(G20), .B(new_n230), .C1(new_n936), .C2(KEYINPUT35), .ZN(new_n937));
  AOI211_X1 g0737(.A(new_n248), .B(new_n937), .C1(KEYINPUT35), .C2(new_n936), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n938), .B(KEYINPUT36), .Z(new_n939));
  OAI211_X1 g0739(.A(G77), .B(new_n228), .C1(new_n417), .C2(new_n216), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(G50), .B2(new_n391), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(G1), .A3(new_n664), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n935), .A2(new_n939), .A3(new_n942), .ZN(G367));
  NOR2_X1   g0743(.A1(new_n818), .A2(new_n427), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n779), .A2(G150), .B1(G50), .B2(new_n831), .ZN(new_n945));
  INV_X1    g0745(.A(new_n770), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n946), .A2(G68), .B1(G137), .B2(new_n766), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n945), .B(new_n947), .C1(new_n833), .C2(new_n774), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n345), .B1(new_n794), .B2(G77), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n944), .B(new_n948), .C1(KEYINPUT110), .C2(new_n949), .ZN(new_n950));
  OAI221_X1 g0750(.A(new_n950), .B1(KEYINPUT110), .B2(new_n949), .C1(new_n216), .C2(new_n796), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n780), .A2(new_n482), .ZN(new_n952));
  INV_X1    g0752(.A(G283), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n345), .B1(new_n787), .B2(new_n953), .C1(new_n786), .C2(new_n774), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n819), .B2(G294), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n794), .A2(G97), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT46), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n796), .A2(new_n957), .A3(new_n248), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n957), .B1(new_n796), .B2(new_n248), .ZN(new_n959));
  INV_X1    g0759(.A(G317), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n959), .B1(new_n960), .B2(new_n765), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n958), .B(new_n961), .C1(G107), .C2(new_n946), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n955), .A2(new_n956), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n951), .B1(new_n952), .B2(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT47), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n748), .B1(new_n965), .B2(new_n758), .ZN(new_n966));
  INV_X1    g0766(.A(new_n749), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n759), .B1(new_n223), .B2(new_n333), .C1(new_n242), .C2(new_n967), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n650), .A2(new_n654), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n573), .A2(new_n671), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT106), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n650), .A2(new_n970), .ZN(new_n972));
  MUX2_X1   g0772(.A(new_n971), .B(KEYINPUT106), .S(new_n972), .Z(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n757), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n966), .A2(new_n968), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n528), .A2(new_n671), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n544), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n639), .A2(new_n671), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n689), .A2(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT45), .ZN(new_n982));
  XOR2_X1   g0782(.A(KEYINPUT108), .B(KEYINPUT44), .Z(new_n983));
  NAND3_X1  g0783(.A1(new_n689), .A2(new_n980), .A3(new_n983), .ZN(new_n984));
  OAI211_X1 g0784(.A(KEYINPUT108), .B(KEYINPUT44), .C1(new_n690), .C2(new_n979), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n982), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n685), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n986), .A2(new_n987), .ZN(new_n990));
  OAI21_X1  g0790(.A(KEYINPUT109), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT109), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n988), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n687), .B1(new_n684), .B2(new_n686), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(new_n676), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n742), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n994), .B(new_n997), .C1(new_n998), .C2(new_n740), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n743), .B1(new_n992), .B2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n693), .B(KEYINPUT41), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n746), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n687), .A2(new_n977), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT42), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n535), .B1(new_n977), .B2(new_n631), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n672), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT43), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n973), .A2(new_n1008), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n973), .A2(new_n1008), .ZN(new_n1010));
  AND3_X1   g0810(.A1(new_n1007), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT107), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1013), .B(new_n1014), .C1(new_n1009), .C2(new_n1007), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n685), .A2(new_n980), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1015), .B(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n975), .B1(new_n1002), .B2(new_n1018), .ZN(G387));
  NAND3_X1  g0819(.A1(new_n741), .A2(new_n742), .A3(new_n996), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(KEYINPUT112), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n743), .A2(new_n997), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n693), .B1(new_n1020), .B2(KEYINPUT112), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n997), .A2(new_n746), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n779), .A2(G317), .B1(new_n775), .B2(G322), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n482), .B2(new_n787), .C1(new_n818), .C2(new_n786), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT48), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n953), .B2(new_n770), .C1(new_n768), .C2(new_n796), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT49), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n766), .A2(new_n776), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n254), .B1(new_n794), .B2(G116), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n774), .A2(new_n427), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n780), .A2(new_n202), .B1(new_n787), .B2(new_n391), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n280), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1038), .B1(new_n1039), .B2(new_n783), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n254), .B1(new_n796), .B2(new_n205), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n770), .A2(new_n333), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1041), .B(new_n1042), .C1(G150), .C2(new_n766), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1040), .A2(new_n956), .A3(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1036), .B1(new_n1037), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n758), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n749), .B1(new_n239), .B2(new_n265), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n695), .B2(new_n753), .ZN(new_n1048));
  AOI211_X1 g0848(.A(G116), .B(new_n562), .C1(G68), .C2(G77), .ZN(new_n1049));
  OR3_X1    g0849(.A1(new_n276), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1050));
  OAI21_X1  g0850(.A(KEYINPUT50), .B1(new_n276), .B2(G50), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n265), .A4(new_n1051), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n1048), .A2(new_n1052), .B1(new_n246), .B2(new_n692), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n759), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n747), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT111), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1046), .B(new_n1056), .C1(new_n684), .C2(new_n761), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1025), .A2(new_n1026), .A3(new_n1057), .ZN(G393));
  OAI21_X1  g0858(.A(new_n693), .B1(new_n999), .B2(new_n992), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n989), .A2(new_n990), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n743), .B2(new_n997), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n746), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n796), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n345), .B1(new_n1064), .B2(new_n210), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n205), .B2(new_n770), .C1(new_n833), .C2(new_n765), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n819), .B2(G50), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n787), .A2(new_n276), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n779), .A2(G159), .B1(new_n775), .B2(G150), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT51), .Z(new_n1070));
  NAND4_X1  g0870(.A1(new_n1067), .A2(new_n822), .A3(new_n1068), .A4(new_n1070), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n345), .B1(new_n248), .B2(new_n770), .C1(new_n818), .C2(new_n482), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(G107), .B2(new_n794), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n779), .A2(G311), .B1(new_n775), .B2(G317), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT52), .Z(new_n1075));
  OAI211_X1 g0875(.A(new_n1073), .B(new_n1075), .C1(new_n768), .C2(new_n787), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n796), .A2(new_n953), .B1(new_n765), .B2(new_n781), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT113), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1071), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n748), .B1(new_n1079), .B2(new_n758), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n249), .A2(new_n749), .B1(G97), .B2(new_n692), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n759), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1080), .B(new_n1082), .C1(new_n761), .C2(new_n979), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1063), .A2(new_n1083), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1062), .A2(new_n1084), .ZN(G390));
  OAI211_X1 g0885(.A(new_n888), .B(new_n896), .C1(new_n898), .C2(new_n907), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n712), .A2(new_n672), .A3(new_n844), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n906), .B1(new_n1087), .B2(new_n845), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n927), .B1(new_n395), .B2(new_n671), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1086), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(G330), .ZN(new_n1091));
  NOR4_X1   g0891(.A1(new_n930), .A2(new_n846), .A3(new_n906), .A4(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n922), .A2(G330), .A3(new_n923), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1086), .B(new_n1094), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1093), .A2(new_n746), .A3(new_n1095), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n770), .A2(new_n427), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1064), .A2(G150), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT53), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1097), .B(new_n1099), .C1(G125), .C2(new_n766), .ZN(new_n1100));
  XOR2_X1   g0900(.A(KEYINPUT54), .B(G143), .Z(new_n1101));
  AOI21_X1  g0901(.A(new_n345), .B1(new_n831), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(G128), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1102), .B1(new_n1103), .B2(new_n774), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n819), .B2(G137), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1100), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(G132), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1106), .B1(new_n202), .B2(new_n793), .C1(new_n1107), .C2(new_n780), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n787), .A2(new_n463), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n780), .A2(new_n248), .B1(new_n774), .B2(new_n953), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n819), .B2(G107), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n345), .B1(new_n765), .B2(new_n768), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n799), .B(new_n1112), .C1(G77), .C2(new_n946), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1111), .A2(new_n826), .A3(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1108), .B1(new_n1109), .B2(new_n1114), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1115), .A2(new_n758), .B1(new_n280), .B2(new_n837), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n747), .B(new_n1116), .C1(new_n897), .C2(new_n756), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1096), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n931), .A2(G330), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n912), .A2(new_n638), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n848), .A2(new_n845), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n923), .B1(new_n922), .B2(G330), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1122), .B1(new_n1123), .B2(new_n1092), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT114), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1123), .A2(new_n1092), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n706), .A2(new_n710), .A3(new_n650), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n710), .B1(new_n706), .B2(new_n650), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n671), .B1(new_n1129), .B2(new_n709), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n839), .B1(new_n1130), .B2(new_n844), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1124), .A2(new_n1125), .B1(new_n1126), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n738), .A2(G330), .A3(new_n842), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n906), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1134), .A2(new_n845), .A3(new_n1087), .A4(new_n1094), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1135), .A2(KEYINPUT114), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1121), .B1(new_n1132), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1138));
  OAI21_X1  g0938(.A(KEYINPUT115), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1122), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n1134), .B2(new_n1094), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1135), .B1(new_n1141), .B2(KEYINPUT114), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1126), .A2(new_n1131), .A3(new_n1125), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1120), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT115), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1144), .A2(new_n1145), .A3(new_n1093), .A4(new_n1095), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1139), .A2(new_n1146), .B1(new_n1138), .B2(new_n1137), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1118), .B1(new_n1147), .B2(new_n693), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(G378));
  NOR2_X1   g0949(.A1(new_n307), .A2(new_n669), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n313), .A2(new_n322), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1151), .B1(new_n313), .B2(new_n322), .ZN(new_n1154));
  OAI21_X1  g0954(.A(KEYINPUT55), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n323), .A2(new_n1150), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT55), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1156), .A2(new_n1157), .A3(new_n1152), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n1155), .A2(KEYINPUT56), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT56), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n755), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n779), .A2(G107), .B1(new_n775), .B2(G116), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1163), .B1(new_n463), .B2(new_n815), .C1(new_n333), .C2(new_n787), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G68), .B2(new_n946), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n794), .A2(G58), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n264), .B1(new_n796), .B2(new_n205), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G283), .B2(new_n766), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1165), .A2(new_n345), .A3(new_n1166), .A4(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT116), .ZN(new_n1170));
  AOI21_X1  g0970(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n1170), .A2(KEYINPUT58), .B1(G50), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT117), .ZN(new_n1173));
  OR2_X1    g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1170), .A2(KEYINPUT58), .ZN(new_n1176));
  AOI21_X1  g0976(.A(G33), .B1(new_n766), .B2(G124), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n264), .B(new_n1177), .C1(new_n793), .C2(new_n427), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT118), .ZN(new_n1179));
  OR2_X1    g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n779), .A2(G128), .B1(new_n1064), .B2(new_n1101), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n946), .A2(G150), .B1(new_n831), .B2(G137), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n783), .A2(G132), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n775), .A2(G125), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  OR2_X1    g0985(.A1(new_n1185), .A2(KEYINPUT59), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(KEYINPUT59), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1180), .A2(new_n1186), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .A4(new_n1189), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1190), .A2(new_n758), .B1(new_n202), .B2(new_n837), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1162), .A2(new_n747), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1161), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n929), .B2(new_n1091), .ZN(new_n1194));
  NOR4_X1   g0994(.A1(new_n930), .A2(new_n846), .A3(new_n906), .A4(new_n925), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n1195), .A2(new_n927), .B1(new_n924), .B2(new_n925), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1196), .A2(G330), .A3(new_n1161), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n1194), .A2(new_n910), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n910), .B1(new_n1194), .B2(new_n1197), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1192), .B1(new_n1200), .B2(new_n745), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1139), .A2(new_n1146), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n1121), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1200), .ZN(new_n1205));
  AOI21_X1  g1005(.A(KEYINPUT57), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n910), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1196), .A2(G330), .A3(new_n1161), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1161), .B1(new_n1196), .B2(G330), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1207), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1194), .A2(new_n910), .A3(new_n1197), .ZN(new_n1211));
  AOI21_X1  g1011(.A(KEYINPUT119), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(KEYINPUT119), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(KEYINPUT57), .B1(new_n1212), .B2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1120), .B1(new_n1139), .B2(new_n1146), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n693), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1202), .B1(new_n1206), .B2(new_n1217), .ZN(G375));
  OAI21_X1  g1018(.A(new_n746), .B1(new_n1132), .B2(new_n1136), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n770), .A2(new_n202), .B1(new_n1103), .B2(new_n765), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n345), .B(new_n1220), .C1(G159), .C2(new_n1064), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1221), .B(new_n1166), .C1(new_n288), .C2(new_n787), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT121), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n819), .A2(new_n1101), .B1(G137), .B2(new_n779), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(new_n1107), .C2(new_n774), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n774), .A2(new_n768), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n345), .B1(new_n246), .B2(new_n787), .C1(new_n780), .C2(new_n953), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n1042), .B(new_n1227), .C1(new_n819), .C2(G116), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n796), .A2(new_n463), .B1(new_n765), .B2(new_n482), .ZN(new_n1229));
  XOR2_X1   g1029(.A(new_n1229), .B(KEYINPUT120), .Z(new_n1230));
  OAI211_X1 g1030(.A(new_n1228), .B(new_n1230), .C1(new_n205), .C2(new_n793), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1225), .B1(new_n1226), .B2(new_n1231), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1232), .A2(new_n758), .B1(new_n391), .B2(new_n837), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n747), .B(new_n1233), .C1(new_n923), .C2(new_n756), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1219), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1142), .A2(new_n1120), .A3(new_n1143), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1137), .A2(new_n1001), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1236), .A2(new_n1238), .ZN(G381));
  INV_X1    g1039(.A(G396), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1025), .A2(new_n1240), .A3(new_n1026), .A4(new_n1057), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(G390), .A2(new_n1241), .A3(G387), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1148), .B(new_n1202), .C1(new_n1206), .C2(new_n1217), .ZN(new_n1244));
  OR4_X1    g1044(.A1(G384), .A2(new_n1243), .A3(G381), .A4(new_n1244), .ZN(G407));
  OAI211_X1 g1045(.A(G407), .B(G213), .C1(G343), .C2(new_n1244), .ZN(G409));
  NOR2_X1   g1046(.A1(new_n1062), .A2(new_n1084), .ZN(new_n1247));
  OR2_X1    g1047(.A1(G387), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(G387), .A2(new_n1247), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(G393), .A2(G396), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n1241), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1250), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT61), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1248), .A2(new_n1241), .A3(new_n1251), .A4(new_n1249), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT124), .ZN(new_n1257));
  OR2_X1    g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1204), .A2(new_n1205), .A3(new_n1001), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n746), .B1(new_n1212), .B2(new_n1214), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1259), .A2(new_n1148), .A3(new_n1192), .A4(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n670), .A2(G213), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT57), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT119), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1263), .B1(new_n1265), .B2(new_n1213), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n694), .B1(new_n1204), .B2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1263), .B1(new_n1216), .B2(new_n1200), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1201), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1261), .B(new_n1262), .C1(new_n1269), .C2(new_n1148), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT60), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1237), .A2(new_n1271), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1272), .A2(new_n1144), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n694), .B1(new_n1237), .B2(new_n1271), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(G384), .B(KEYINPUT122), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1275), .A2(new_n1236), .A3(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1235), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G384), .A2(KEYINPUT122), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1277), .B1(new_n1278), .B2(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1270), .A2(new_n1281), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n1256), .A2(new_n1257), .B1(new_n1282), .B2(KEYINPUT63), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1262), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1284), .A2(KEYINPUT123), .A3(G2897), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1277), .B(new_n1285), .C1(new_n1278), .C2(new_n1280), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT123), .B1(new_n1284), .B2(G2897), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(new_n1286), .B(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1270), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1289), .A2(KEYINPUT63), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1258), .B(new_n1283), .C1(new_n1282), .C2(new_n1290), .ZN(new_n1291));
  OR3_X1    g1091(.A1(new_n1270), .A2(KEYINPUT62), .A3(new_n1281), .ZN(new_n1292));
  OAI21_X1  g1092(.A(KEYINPUT62), .B1(new_n1270), .B2(new_n1281), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT125), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1295), .B1(new_n1289), .B2(new_n1254), .ZN(new_n1296));
  AOI211_X1 g1096(.A(KEYINPUT125), .B(KEYINPUT61), .C1(new_n1288), .C2(new_n1270), .ZN(new_n1297));
  NOR3_X1   g1097(.A1(new_n1294), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1253), .A2(new_n1255), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1291), .B1(new_n1298), .B2(new_n1300), .ZN(G405));
  INV_X1    g1101(.A(new_n1281), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1244), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1204), .A2(new_n1266), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1304), .A2(new_n1268), .A3(new_n693), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1148), .B1(new_n1305), .B2(new_n1202), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1302), .B1(new_n1303), .B2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(G375), .A2(G378), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1308), .A2(new_n1244), .A3(new_n1281), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1307), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT126), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1299), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1307), .A2(KEYINPUT126), .A3(new_n1309), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(KEYINPUT127), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT127), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1307), .A2(KEYINPUT126), .A3(new_n1309), .A4(new_n1315), .ZN(new_n1316));
  AND3_X1   g1116(.A1(new_n1312), .A2(new_n1314), .A3(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1318));
  AOI22_X1  g1118(.A1(new_n1314), .A2(new_n1316), .B1(new_n1318), .B2(new_n1300), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1317), .A2(new_n1319), .ZN(G402));
endmodule


