

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595;

  XNOR2_X1 U324 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U325 ( .A(n487), .B(KEYINPUT65), .ZN(n582) );
  XNOR2_X1 U326 ( .A(n356), .B(n327), .ZN(n331) );
  XOR2_X1 U327 ( .A(n438), .B(n437), .Z(n572) );
  XNOR2_X1 U328 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U329 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U330 ( .A(n461), .B(KEYINPUT109), .ZN(n527) );
  XOR2_X1 U331 ( .A(n488), .B(KEYINPUT28), .Z(n545) );
  XNOR2_X1 U332 ( .A(n342), .B(n334), .ZN(n534) );
  XOR2_X1 U333 ( .A(n485), .B(n484), .Z(n292) );
  AND2_X1 U334 ( .A1(n572), .A2(n561), .ZN(n472) );
  INV_X1 U335 ( .A(KEYINPUT90), .ZN(n351) );
  XNOR2_X1 U336 ( .A(n352), .B(n351), .ZN(n353) );
  AND2_X1 U337 ( .A1(n479), .A2(n478), .ZN(n480) );
  XNOR2_X1 U338 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U339 ( .A(G92GAT), .B(G85GAT), .Z(n440) );
  INV_X1 U340 ( .A(n385), .ZN(n360) );
  XNOR2_X1 U341 ( .A(n326), .B(KEYINPUT95), .ZN(n327) );
  INV_X1 U342 ( .A(n532), .ZN(n486) );
  XNOR2_X1 U343 ( .A(n489), .B(KEYINPUT55), .ZN(n490) );
  XNOR2_X1 U344 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U345 ( .A(KEYINPUT106), .B(KEYINPUT36), .ZN(n466) );
  XNOR2_X1 U346 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U347 ( .A(n363), .B(n362), .ZN(n367) );
  XNOR2_X1 U348 ( .A(n504), .B(n466), .ZN(n593) );
  XNOR2_X1 U349 ( .A(n415), .B(n414), .ZN(n420) );
  XOR2_X1 U350 ( .A(n460), .B(KEYINPUT41), .Z(n561) );
  INV_X1 U351 ( .A(G57GAT), .ZN(n462) );
  XOR2_X1 U352 ( .A(KEYINPUT38), .B(n499), .Z(n522) );
  XNOR2_X1 U353 ( .A(n505), .B(KEYINPUT58), .ZN(n506) );
  XNOR2_X1 U354 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U355 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U356 ( .A(n507), .B(n506), .ZN(G1351GAT) );
  XNOR2_X1 U357 ( .A(n465), .B(n464), .ZN(G1332GAT) );
  XOR2_X1 U358 ( .A(G127GAT), .B(KEYINPUT81), .Z(n294) );
  XNOR2_X1 U359 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n293) );
  XNOR2_X1 U360 ( .A(n294), .B(n293), .ZN(n339) );
  XOR2_X1 U361 ( .A(n339), .B(G134GAT), .Z(n296) );
  NAND2_X1 U362 ( .A1(G225GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U363 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U364 ( .A(G29GAT), .B(n297), .ZN(n314) );
  XOR2_X1 U365 ( .A(KEYINPUT4), .B(KEYINPUT92), .Z(n299) );
  XNOR2_X1 U366 ( .A(KEYINPUT93), .B(KEYINPUT5), .ZN(n298) );
  XNOR2_X1 U367 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U368 ( .A(G57GAT), .B(G155GAT), .Z(n301) );
  XNOR2_X1 U369 ( .A(G1GAT), .B(G120GAT), .ZN(n300) );
  XNOR2_X1 U370 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U371 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U372 ( .A(G85GAT), .B(KEYINPUT76), .Z(n305) );
  XNOR2_X1 U373 ( .A(G148GAT), .B(G162GAT), .ZN(n304) );
  XNOR2_X1 U374 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U375 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U376 ( .A(n308), .B(KEYINPUT1), .Z(n312) );
  XOR2_X1 U377 ( .A(KEYINPUT2), .B(KEYINPUT89), .Z(n310) );
  XNOR2_X1 U378 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n309) );
  XNOR2_X1 U379 ( .A(n310), .B(n309), .ZN(n359) );
  XNOR2_X1 U380 ( .A(n359), .B(KEYINPUT6), .ZN(n311) );
  XNOR2_X1 U381 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U382 ( .A(n314), .B(n313), .ZN(n532) );
  XNOR2_X1 U383 ( .A(KEYINPUT27), .B(KEYINPUT98), .ZN(n335) );
  XOR2_X1 U384 ( .A(G183GAT), .B(KEYINPUT19), .Z(n316) );
  XNOR2_X1 U385 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n315) );
  XNOR2_X1 U386 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U387 ( .A(KEYINPUT18), .B(KEYINPUT83), .Z(n318) );
  XNOR2_X1 U388 ( .A(G190GAT), .B(KEYINPUT84), .ZN(n317) );
  XNOR2_X1 U389 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U390 ( .A(n320), .B(n319), .Z(n342) );
  XOR2_X1 U391 ( .A(KEYINPUT88), .B(G218GAT), .Z(n322) );
  XNOR2_X1 U392 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n321) );
  XNOR2_X1 U393 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U394 ( .A(G197GAT), .B(n323), .Z(n356) );
  XOR2_X1 U395 ( .A(KEYINPUT94), .B(KEYINPUT97), .Z(n325) );
  NAND2_X1 U396 ( .A1(G226GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U397 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U398 ( .A(G176GAT), .B(G64GAT), .Z(n449) );
  XOR2_X1 U399 ( .A(G92GAT), .B(n449), .Z(n329) );
  XOR2_X1 U400 ( .A(G36GAT), .B(KEYINPUT77), .Z(n412) );
  XNOR2_X1 U401 ( .A(G204GAT), .B(n412), .ZN(n328) );
  XNOR2_X1 U402 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U403 ( .A(n331), .B(n330), .Z(n333) );
  XNOR2_X1 U404 ( .A(G8GAT), .B(KEYINPUT96), .ZN(n332) );
  XNOR2_X1 U405 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U406 ( .A(n335), .B(n534), .Z(n376) );
  INV_X1 U407 ( .A(n376), .ZN(n336) );
  NAND2_X1 U408 ( .A1(n532), .A2(n336), .ZN(n541) );
  XOR2_X1 U409 ( .A(G43GAT), .B(G134GAT), .Z(n411) );
  XOR2_X1 U410 ( .A(G176GAT), .B(KEYINPUT20), .Z(n338) );
  XNOR2_X1 U411 ( .A(G15GAT), .B(KEYINPUT82), .ZN(n337) );
  XNOR2_X1 U412 ( .A(n338), .B(n337), .ZN(n340) );
  XOR2_X1 U413 ( .A(n340), .B(n339), .Z(n344) );
  XNOR2_X1 U414 ( .A(G99GAT), .B(G71GAT), .ZN(n341) );
  XNOR2_X1 U415 ( .A(n341), .B(G120GAT), .ZN(n452) );
  XNOR2_X1 U416 ( .A(n342), .B(n452), .ZN(n343) );
  XNOR2_X1 U417 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U418 ( .A(n411), .B(n345), .Z(n347) );
  NAND2_X1 U419 ( .A1(G227GAT), .A2(G233GAT), .ZN(n346) );
  XOR2_X2 U420 ( .A(n347), .B(n346), .Z(n546) );
  XOR2_X1 U421 ( .A(KEYINPUT85), .B(n546), .Z(n348) );
  NOR2_X1 U422 ( .A1(n541), .A2(n348), .ZN(n369) );
  XOR2_X1 U423 ( .A(KEYINPUT91), .B(KEYINPUT24), .Z(n350) );
  XNOR2_X1 U424 ( .A(KEYINPUT22), .B(KEYINPUT87), .ZN(n349) );
  XNOR2_X1 U425 ( .A(n350), .B(n349), .ZN(n354) );
  NAND2_X1 U426 ( .A1(G228GAT), .A2(G233GAT), .ZN(n352) );
  XOR2_X1 U427 ( .A(n355), .B(KEYINPUT23), .Z(n358) );
  XNOR2_X1 U428 ( .A(n356), .B(KEYINPUT86), .ZN(n357) );
  XNOR2_X1 U429 ( .A(n358), .B(n357), .ZN(n363) );
  XOR2_X1 U430 ( .A(G50GAT), .B(G162GAT), .Z(n401) );
  XNOR2_X1 U431 ( .A(n401), .B(n359), .ZN(n361) );
  XOR2_X1 U432 ( .A(G22GAT), .B(G155GAT), .Z(n385) );
  XOR2_X1 U433 ( .A(G148GAT), .B(G106GAT), .Z(n365) );
  XNOR2_X1 U434 ( .A(G204GAT), .B(G78GAT), .ZN(n364) );
  XNOR2_X1 U435 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U436 ( .A(KEYINPUT70), .B(n366), .Z(n439) );
  XOR2_X1 U437 ( .A(n367), .B(n439), .Z(n488) );
  INV_X1 U438 ( .A(n545), .ZN(n368) );
  NAND2_X1 U439 ( .A1(n369), .A2(n368), .ZN(n370) );
  XNOR2_X1 U440 ( .A(n370), .B(KEYINPUT99), .ZN(n382) );
  NAND2_X1 U441 ( .A1(n546), .A2(n534), .ZN(n371) );
  XNOR2_X1 U442 ( .A(KEYINPUT100), .B(n371), .ZN(n372) );
  NAND2_X1 U443 ( .A1(n372), .A2(n488), .ZN(n374) );
  XOR2_X1 U444 ( .A(KEYINPUT25), .B(KEYINPUT101), .Z(n373) );
  XNOR2_X1 U445 ( .A(n374), .B(n373), .ZN(n378) );
  NOR2_X1 U446 ( .A1(n488), .A2(n546), .ZN(n375) );
  XNOR2_X1 U447 ( .A(KEYINPUT26), .B(n375), .ZN(n581) );
  INV_X1 U448 ( .A(n581), .ZN(n559) );
  NOR2_X1 U449 ( .A1(n559), .A2(n376), .ZN(n377) );
  NOR2_X1 U450 ( .A1(n378), .A2(n377), .ZN(n379) );
  XNOR2_X1 U451 ( .A(KEYINPUT102), .B(n379), .ZN(n380) );
  NOR2_X1 U452 ( .A1(n380), .A2(n532), .ZN(n381) );
  NOR2_X1 U453 ( .A1(n382), .A2(n381), .ZN(n383) );
  XOR2_X1 U454 ( .A(KEYINPUT103), .B(n383), .Z(n496) );
  XNOR2_X1 U455 ( .A(G57GAT), .B(KEYINPUT67), .ZN(n384) );
  XNOR2_X1 U456 ( .A(n384), .B(KEYINPUT13), .ZN(n441) );
  XOR2_X1 U457 ( .A(n441), .B(n385), .Z(n387) );
  XNOR2_X1 U458 ( .A(G78GAT), .B(G211GAT), .ZN(n386) );
  XNOR2_X1 U459 ( .A(n387), .B(n386), .ZN(n392) );
  XNOR2_X1 U460 ( .A(G15GAT), .B(G8GAT), .ZN(n388) );
  XNOR2_X1 U461 ( .A(n388), .B(G1GAT), .ZN(n433) );
  XOR2_X1 U462 ( .A(n433), .B(KEYINPUT78), .Z(n390) );
  NAND2_X1 U463 ( .A1(G231GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U464 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U465 ( .A(n392), .B(n391), .Z(n400) );
  XOR2_X1 U466 ( .A(G64GAT), .B(G127GAT), .Z(n394) );
  XNOR2_X1 U467 ( .A(G183GAT), .B(G71GAT), .ZN(n393) );
  XNOR2_X1 U468 ( .A(n394), .B(n393), .ZN(n398) );
  XOR2_X1 U469 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n396) );
  XNOR2_X1 U470 ( .A(KEYINPUT15), .B(KEYINPUT79), .ZN(n395) );
  XNOR2_X1 U471 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U472 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U473 ( .A(n400), .B(n399), .Z(n566) );
  INV_X1 U474 ( .A(n566), .ZN(n590) );
  XNOR2_X1 U475 ( .A(n440), .B(n401), .ZN(n403) );
  XOR2_X1 U476 ( .A(G106GAT), .B(G218GAT), .Z(n402) );
  XNOR2_X1 U477 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U478 ( .A(n404), .B(KEYINPUT66), .Z(n409) );
  XOR2_X1 U479 ( .A(KEYINPUT74), .B(KEYINPUT9), .Z(n406) );
  XNOR2_X1 U480 ( .A(G99GAT), .B(KEYINPUT75), .ZN(n405) );
  XNOR2_X1 U481 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U482 ( .A(G190GAT), .B(n407), .ZN(n408) );
  XNOR2_X1 U483 ( .A(n409), .B(n408), .ZN(n415) );
  XNOR2_X1 U484 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n410) );
  XNOR2_X1 U485 ( .A(n410), .B(KEYINPUT8), .ZN(n434) );
  XOR2_X1 U486 ( .A(n434), .B(n411), .Z(n413) );
  XOR2_X1 U487 ( .A(KEYINPUT10), .B(KEYINPUT76), .Z(n417) );
  NAND2_X1 U488 ( .A1(G232GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U489 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U490 ( .A(KEYINPUT11), .B(n418), .Z(n419) );
  XNOR2_X1 U491 ( .A(n420), .B(n419), .ZN(n570) );
  NOR2_X1 U492 ( .A1(n590), .A2(n570), .ZN(n421) );
  XOR2_X1 U493 ( .A(KEYINPUT80), .B(n421), .Z(n422) );
  XNOR2_X1 U494 ( .A(n422), .B(KEYINPUT16), .ZN(n423) );
  NOR2_X1 U495 ( .A1(n496), .A2(n423), .ZN(n424) );
  XNOR2_X1 U496 ( .A(KEYINPUT104), .B(n424), .ZN(n508) );
  XOR2_X1 U497 ( .A(G43GAT), .B(G36GAT), .Z(n426) );
  NAND2_X1 U498 ( .A1(G229GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U499 ( .A(n426), .B(n425), .ZN(n438) );
  XOR2_X1 U500 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n428) );
  XNOR2_X1 U501 ( .A(G169GAT), .B(G113GAT), .ZN(n427) );
  XNOR2_X1 U502 ( .A(n428), .B(n427), .ZN(n432) );
  XOR2_X1 U503 ( .A(G197GAT), .B(G22GAT), .Z(n430) );
  XNOR2_X1 U504 ( .A(G50GAT), .B(G141GAT), .ZN(n429) );
  XNOR2_X1 U505 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U506 ( .A(n432), .B(n431), .Z(n436) );
  XNOR2_X1 U507 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U508 ( .A(n436), .B(n435), .ZN(n437) );
  INV_X1 U509 ( .A(n439), .ZN(n445) );
  XOR2_X1 U510 ( .A(n441), .B(n440), .Z(n443) );
  NAND2_X1 U511 ( .A1(G230GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U512 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U513 ( .A(n445), .B(n444), .ZN(n458) );
  XOR2_X1 U514 ( .A(KEYINPUT31), .B(KEYINPUT72), .Z(n447) );
  XNOR2_X1 U515 ( .A(KEYINPUT68), .B(KEYINPUT71), .ZN(n446) );
  XNOR2_X1 U516 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U517 ( .A(n448), .B(KEYINPUT69), .ZN(n451) );
  XOR2_X1 U518 ( .A(n449), .B(KEYINPUT73), .Z(n450) );
  XNOR2_X1 U519 ( .A(n451), .B(n450), .ZN(n456) );
  XNOR2_X1 U520 ( .A(n452), .B(KEYINPUT33), .ZN(n454) );
  INV_X1 U521 ( .A(KEYINPUT32), .ZN(n453) );
  XNOR2_X1 U522 ( .A(n458), .B(n457), .ZN(n587) );
  INV_X1 U523 ( .A(KEYINPUT64), .ZN(n459) );
  XNOR2_X1 U524 ( .A(n587), .B(n459), .ZN(n460) );
  INV_X1 U525 ( .A(n561), .ZN(n578) );
  NOR2_X1 U526 ( .A1(n572), .A2(n578), .ZN(n530) );
  NAND2_X1 U527 ( .A1(n508), .A2(n530), .ZN(n461) );
  NAND2_X1 U528 ( .A1(n527), .A2(n532), .ZN(n465) );
  XOR2_X1 U529 ( .A(KEYINPUT42), .B(KEYINPUT110), .Z(n463) );
  XOR2_X1 U530 ( .A(KEYINPUT121), .B(KEYINPUT54), .Z(n485) );
  XNOR2_X1 U531 ( .A(KEYINPUT45), .B(KEYINPUT115), .ZN(n468) );
  INV_X1 U532 ( .A(n570), .ZN(n504) );
  NOR2_X1 U533 ( .A1(n593), .A2(n590), .ZN(n467) );
  XNOR2_X1 U534 ( .A(n468), .B(n467), .ZN(n469) );
  NOR2_X1 U535 ( .A1(n469), .A2(n572), .ZN(n470) );
  NAND2_X1 U536 ( .A1(n587), .A2(n470), .ZN(n479) );
  XOR2_X1 U537 ( .A(KEYINPUT113), .B(KEYINPUT46), .Z(n471) );
  XNOR2_X1 U538 ( .A(n472), .B(n471), .ZN(n474) );
  OR2_X1 U539 ( .A1(n570), .A2(n566), .ZN(n473) );
  NOR2_X1 U540 ( .A1(n474), .A2(n473), .ZN(n476) );
  XNOR2_X1 U541 ( .A(KEYINPUT47), .B(KEYINPUT114), .ZN(n475) );
  XNOR2_X1 U542 ( .A(n476), .B(n475), .ZN(n481) );
  NAND2_X1 U543 ( .A1(n479), .A2(n481), .ZN(n477) );
  NAND2_X1 U544 ( .A1(n477), .A2(KEYINPUT48), .ZN(n483) );
  INV_X1 U545 ( .A(KEYINPUT48), .ZN(n478) );
  NAND2_X1 U546 ( .A1(n481), .A2(n480), .ZN(n482) );
  NAND2_X1 U547 ( .A1(n483), .A2(n482), .ZN(n543) );
  NAND2_X1 U548 ( .A1(n543), .A2(n534), .ZN(n484) );
  NAND2_X1 U549 ( .A1(n292), .A2(n486), .ZN(n487) );
  NAND2_X1 U550 ( .A1(n582), .A2(n488), .ZN(n491) );
  XOR2_X1 U551 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n489) );
  AND2_X1 U552 ( .A1(n546), .A2(n492), .ZN(n493) );
  XOR2_X1 U553 ( .A(n493), .B(KEYINPUT124), .Z(n577) );
  NOR2_X1 U554 ( .A1(n577), .A2(n590), .ZN(n495) );
  INV_X1 U555 ( .A(G183GAT), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n495), .B(n494), .ZN(G1350GAT) );
  NOR2_X1 U557 ( .A1(n593), .A2(n496), .ZN(n497) );
  NAND2_X1 U558 ( .A1(n497), .A2(n590), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n498), .B(KEYINPUT37), .ZN(n531) );
  AND2_X1 U560 ( .A1(n587), .A2(n572), .ZN(n509) );
  NAND2_X1 U561 ( .A1(n531), .A2(n509), .ZN(n499) );
  NAND2_X1 U562 ( .A1(n522), .A2(n546), .ZN(n503) );
  XOR2_X1 U563 ( .A(KEYINPUT108), .B(KEYINPUT40), .Z(n501) );
  INV_X1 U564 ( .A(G43GAT), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n503), .B(n502), .ZN(G1330GAT) );
  NOR2_X1 U566 ( .A1(n577), .A2(n504), .ZN(n507) );
  INV_X1 U567 ( .A(G190GAT), .ZN(n505) );
  AND2_X1 U568 ( .A1(n509), .A2(n508), .ZN(n515) );
  NAND2_X1 U569 ( .A1(n532), .A2(n515), .ZN(n510) );
  XNOR2_X1 U570 ( .A(KEYINPUT34), .B(n510), .ZN(n511) );
  XNOR2_X1 U571 ( .A(G1GAT), .B(n511), .ZN(G1324GAT) );
  NAND2_X1 U572 ( .A1(n534), .A2(n515), .ZN(n512) );
  XNOR2_X1 U573 ( .A(n512), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U574 ( .A(G15GAT), .B(KEYINPUT35), .Z(n514) );
  NAND2_X1 U575 ( .A1(n515), .A2(n546), .ZN(n513) );
  XNOR2_X1 U576 ( .A(n514), .B(n513), .ZN(G1326GAT) );
  XOR2_X1 U577 ( .A(G22GAT), .B(KEYINPUT105), .Z(n517) );
  NAND2_X1 U578 ( .A1(n515), .A2(n545), .ZN(n516) );
  XNOR2_X1 U579 ( .A(n517), .B(n516), .ZN(G1327GAT) );
  XOR2_X1 U580 ( .A(G29GAT), .B(KEYINPUT39), .Z(n519) );
  NAND2_X1 U581 ( .A1(n532), .A2(n522), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n519), .B(n518), .ZN(G1328GAT) );
  XOR2_X1 U583 ( .A(G36GAT), .B(KEYINPUT107), .Z(n521) );
  NAND2_X1 U584 ( .A1(n522), .A2(n534), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n521), .B(n520), .ZN(G1329GAT) );
  NAND2_X1 U586 ( .A1(n545), .A2(n522), .ZN(n523) );
  XNOR2_X1 U587 ( .A(G50GAT), .B(n523), .ZN(G1331GAT) );
  XOR2_X1 U588 ( .A(G64GAT), .B(KEYINPUT111), .Z(n525) );
  NAND2_X1 U589 ( .A1(n527), .A2(n534), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(G1333GAT) );
  NAND2_X1 U591 ( .A1(n546), .A2(n527), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n526), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U593 ( .A(G78GAT), .B(KEYINPUT43), .Z(n529) );
  NAND2_X1 U594 ( .A1(n527), .A2(n545), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n529), .B(n528), .ZN(G1335GAT) );
  AND2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n537) );
  NAND2_X1 U597 ( .A1(n532), .A2(n537), .ZN(n533) );
  XNOR2_X1 U598 ( .A(G85GAT), .B(n533), .ZN(G1336GAT) );
  NAND2_X1 U599 ( .A1(n534), .A2(n537), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n535), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U601 ( .A1(n546), .A2(n537), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n536), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT44), .B(KEYINPUT112), .Z(n539) );
  NAND2_X1 U604 ( .A1(n537), .A2(n545), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U606 ( .A(G106GAT), .B(n540), .Z(G1339GAT) );
  INV_X1 U607 ( .A(n541), .ZN(n542) );
  NAND2_X1 U608 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U609 ( .A(KEYINPUT116), .B(n544), .ZN(n558) );
  NOR2_X1 U610 ( .A1(n545), .A2(n558), .ZN(n547) );
  NAND2_X1 U611 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U612 ( .A(KEYINPUT117), .B(n548), .ZN(n555) );
  NAND2_X1 U613 ( .A1(n555), .A2(n572), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n549), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U615 ( .A(G120GAT), .B(KEYINPUT49), .Z(n551) );
  NAND2_X1 U616 ( .A1(n555), .A2(n561), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(G1341GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n553) );
  NAND2_X1 U619 ( .A1(n555), .A2(n566), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U621 ( .A(G127GAT), .B(n554), .Z(G1342GAT) );
  XOR2_X1 U622 ( .A(G134GAT), .B(KEYINPUT51), .Z(n557) );
  NAND2_X1 U623 ( .A1(n555), .A2(n570), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1343GAT) );
  NOR2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n569) );
  NAND2_X1 U626 ( .A1(n572), .A2(n569), .ZN(n560) );
  XNOR2_X1 U627 ( .A(G141GAT), .B(n560), .ZN(G1344GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n563) );
  NAND2_X1 U629 ( .A1(n569), .A2(n561), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n565) );
  XOR2_X1 U631 ( .A(G148GAT), .B(KEYINPUT52), .Z(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(G1345GAT) );
  NAND2_X1 U633 ( .A1(n566), .A2(n569), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(KEYINPUT120), .ZN(n568) );
  XNOR2_X1 U635 ( .A(G155GAT), .B(n568), .ZN(G1346GAT) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(G162GAT), .ZN(G1347GAT) );
  INV_X1 U638 ( .A(n572), .ZN(n583) );
  NOR2_X1 U639 ( .A1(n577), .A2(n583), .ZN(n573) );
  XOR2_X1 U640 ( .A(G169GAT), .B(n573), .Z(G1348GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT57), .B(KEYINPUT126), .Z(n575) );
  XNOR2_X1 U642 ( .A(G176GAT), .B(KEYINPUT125), .ZN(n574) );
  XNOR2_X1 U643 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U644 ( .A(KEYINPUT56), .B(n576), .ZN(n580) );
  NOR2_X1 U645 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(G1349GAT) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n592) );
  NOR2_X1 U648 ( .A1(n583), .A2(n592), .ZN(n585) );
  XNOR2_X1 U649 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(G197GAT), .B(n586), .ZN(G1352GAT) );
  NOR2_X1 U652 ( .A1(n587), .A2(n592), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(G1353GAT) );
  NOR2_X1 U655 ( .A1(n590), .A2(n592), .ZN(n591) );
  XOR2_X1 U656 ( .A(G211GAT), .B(n591), .Z(G1354GAT) );
  NOR2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U658 ( .A(KEYINPUT62), .B(n594), .Z(n595) );
  XNOR2_X1 U659 ( .A(G218GAT), .B(n595), .ZN(G1355GAT) );
endmodule

