//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0 1 0 0 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n872, new_n873, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n988,
    new_n989;
  INV_X1    g000(.A(KEYINPUT3), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT74), .ZN(new_n203));
  INV_X1    g002(.A(G155gat), .ZN(new_n204));
  INV_X1    g003(.A(G162gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT73), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G141gat), .ZN(new_n207));
  INV_X1    g006(.A(G148gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n212), .B1(G155gat), .B2(G162gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n206), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G155gat), .B(G162gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT2), .B1(new_n204), .B2(new_n205), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(new_n209), .A3(new_n210), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n215), .B1(new_n219), .B2(new_n206), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n203), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n214), .A2(new_n216), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n219), .A2(new_n215), .A3(new_n206), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(new_n223), .A3(KEYINPUT74), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n202), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G127gat), .ZN(new_n226));
  INV_X1    g025(.A(G134gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G113gat), .B(G120gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT65), .B(G134gat), .ZN(new_n230));
  OAI221_X1 g029(.A(new_n228), .B1(new_n229), .B2(KEYINPUT1), .C1(new_n226), .C2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT1), .ZN(new_n234));
  XNOR2_X1  g033(.A(G127gat), .B(G134gat), .ZN(new_n235));
  INV_X1    g034(.A(G120gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n236), .A2(KEYINPUT66), .A3(G113gat), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n233), .A2(new_n234), .A3(new_n235), .A4(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n231), .A2(new_n238), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n217), .A2(new_n220), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n239), .B1(new_n240), .B2(KEYINPUT3), .ZN(new_n241));
  OR2_X1    g040(.A1(new_n225), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G225gat), .A2(G233gat), .ZN(new_n243));
  XOR2_X1   g042(.A(new_n243), .B(KEYINPUT75), .Z(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  AND2_X1   g044(.A1(new_n231), .A2(new_n238), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n222), .A2(new_n223), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(KEYINPUT4), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT4), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n249), .B1(new_n240), .B2(new_n239), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n242), .A2(new_n245), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n246), .B1(new_n224), .B2(new_n221), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n240), .A2(new_n239), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n244), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT76), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI211_X1 g056(.A(KEYINPUT76), .B(new_n244), .C1(new_n253), .C2(new_n254), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n252), .A2(new_n257), .A3(KEYINPUT5), .A4(new_n258), .ZN(new_n259));
  XOR2_X1   g058(.A(G1gat), .B(G29gat), .Z(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(G57gat), .B(G85gat), .Z(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n250), .B(new_n248), .C1(new_n225), .C2(new_n241), .ZN(new_n265));
  OR3_X1    g064(.A1(new_n265), .A2(KEYINPUT5), .A3(new_n244), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n259), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT6), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT80), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n259), .A2(new_n266), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n264), .B(KEYINPUT79), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n272), .ZN(new_n274));
  AOI211_X1 g073(.A(KEYINPUT80), .B(new_n274), .C1(new_n259), .C2(new_n266), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n269), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT81), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n264), .B1(new_n259), .B2(new_n266), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT6), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n269), .B(KEYINPUT81), .C1(new_n273), .C2(new_n275), .ZN(new_n281));
  INV_X1    g080(.A(G226gat), .ZN(new_n282));
  INV_X1    g081(.A(G233gat), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n286));
  MUX2_X1   g085(.A(G183gat), .B(new_n286), .S(G190gat), .Z(new_n287));
  NAND2_X1  g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT24), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT23), .ZN(new_n293));
  NAND2_X1  g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT23), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(G169gat), .B2(G176gat), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n293), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT25), .B1(new_n291), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n293), .A2(KEYINPUT25), .A3(new_n296), .A4(new_n294), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT24), .B1(new_n288), .B2(KEYINPUT64), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n301), .B1(KEYINPUT64), .B2(new_n288), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n300), .B1(new_n287), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT27), .B(G183gat), .ZN(new_n305));
  INV_X1    g104(.A(G190gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT28), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n305), .A2(KEYINPUT28), .A3(new_n306), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n292), .A2(KEYINPUT26), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(new_n288), .ZN(new_n313));
  INV_X1    g112(.A(G169gat), .ZN(new_n314));
  INV_X1    g113(.A(G176gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n313), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n299), .A2(new_n304), .B1(new_n311), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n285), .B1(new_n319), .B2(KEYINPUT29), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n299), .A2(new_n304), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n311), .A2(new_n318), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(new_n284), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT70), .B(G197gat), .ZN(new_n325));
  INV_X1    g124(.A(G204gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n325), .B(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT22), .ZN(new_n328));
  INV_X1    g127(.A(G211gat), .ZN(new_n329));
  INV_X1    g128(.A(G218gat), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G211gat), .B(G218gat), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n327), .A2(new_n333), .A3(new_n331), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n320), .A2(new_n324), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n337), .B1(new_n320), .B2(new_n324), .ZN(new_n340));
  OAI21_X1  g139(.A(KEYINPUT37), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  XOR2_X1   g140(.A(KEYINPUT82), .B(KEYINPUT38), .Z(new_n342));
  XNOR2_X1  g141(.A(G8gat), .B(G36gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(G64gat), .B(G92gat), .ZN(new_n344));
  XOR2_X1   g143(.A(new_n343), .B(new_n344), .Z(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n335), .A2(new_n336), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT29), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n284), .B1(new_n323), .B2(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n319), .A2(new_n285), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n347), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT37), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(new_n352), .A3(new_n338), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n341), .A2(new_n342), .A3(new_n346), .A4(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n351), .A2(new_n338), .A3(new_n345), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT72), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT72), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n351), .A2(new_n338), .A3(new_n357), .A4(new_n345), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n354), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n342), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT83), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n352), .B1(new_n351), .B2(new_n338), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n361), .B1(new_n362), .B2(new_n345), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n341), .A2(KEYINPUT83), .A3(new_n346), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n363), .A2(new_n364), .A3(new_n353), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n359), .B1(new_n360), .B2(new_n365), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n278), .A2(new_n280), .A3(new_n281), .A4(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n221), .A2(new_n224), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT29), .B1(new_n335), .B2(new_n336), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n368), .B1(new_n369), .B2(KEYINPUT3), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n240), .A2(KEYINPUT3), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n347), .B1(KEYINPUT29), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G228gat), .A2(G233gat), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT78), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n335), .A2(new_n377), .A3(new_n336), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n333), .B1(new_n327), .B2(new_n331), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT29), .B1(new_n379), .B2(KEYINPUT78), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT3), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n372), .B(new_n374), .C1(new_n381), .C2(new_n247), .ZN(new_n382));
  XNOR2_X1  g181(.A(KEYINPUT31), .B(G50gat), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n376), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n384), .B1(new_n376), .B2(new_n382), .ZN(new_n386));
  XNOR2_X1  g185(.A(G78gat), .B(G106gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(G22gat), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NOR3_X1   g188(.A1(new_n385), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n382), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n374), .B1(new_n370), .B2(new_n372), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n383), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n382), .A3(new_n384), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n388), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n265), .A2(new_n244), .ZN(new_n398));
  OR3_X1    g197(.A1(new_n253), .A2(new_n244), .A3(new_n254), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n399), .A3(KEYINPUT39), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT39), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n265), .A2(new_n401), .A3(new_n244), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n400), .A2(new_n274), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT40), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n403), .B(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n271), .A2(new_n272), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT80), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n271), .A2(new_n270), .A3(new_n272), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n346), .B1(new_n339), .B2(new_n340), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT71), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT71), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n412), .B(new_n346), .C1(new_n339), .C2(new_n340), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT30), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n356), .A2(new_n415), .A3(new_n358), .ZN(new_n416));
  OR2_X1    g215(.A1(new_n355), .A2(new_n415), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n414), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n397), .B1(new_n409), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n367), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n267), .A2(new_n268), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n280), .B1(new_n421), .B2(new_n279), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n414), .A2(new_n416), .A3(new_n417), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n396), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n321), .A2(new_n239), .A3(new_n322), .ZN(new_n425));
  AND2_X1   g224(.A1(new_n311), .A2(new_n318), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n298), .A2(new_n303), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n246), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(G227gat), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n429), .A2(new_n283), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n425), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT32), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT33), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(KEYINPUT67), .B(G71gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n437), .B(G99gat), .ZN(new_n438));
  XOR2_X1   g237(.A(G15gat), .B(G43gat), .Z(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  AND2_X1   g241(.A1(new_n425), .A2(new_n428), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT34), .B1(new_n443), .B2(new_n430), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n430), .B1(new_n425), .B2(new_n428), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT34), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n442), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n440), .B1(new_n431), .B2(new_n435), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n445), .A2(new_n446), .ZN(new_n450));
  AOI211_X1 g249(.A(KEYINPUT34), .B(new_n430), .C1(new_n425), .C2(new_n428), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n434), .B1(new_n448), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n448), .A2(new_n434), .A3(new_n452), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n454), .A2(KEYINPUT36), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT68), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n448), .A2(new_n434), .A3(new_n452), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n459), .A2(new_n453), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n460), .A2(KEYINPUT68), .A3(KEYINPUT36), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT36), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n463), .B1(new_n459), .B2(new_n453), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT69), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT69), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n466), .B(new_n463), .C1(new_n459), .C2(new_n453), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n424), .B1(new_n462), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n389), .B1(new_n385), .B2(new_n386), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n393), .A2(new_n388), .A3(new_n394), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n454), .A2(new_n470), .A3(new_n471), .A4(new_n455), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n472), .A2(KEYINPUT35), .A3(new_n418), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n281), .A2(new_n280), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n407), .A2(new_n408), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT81), .B1(new_n475), .B2(new_n269), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n473), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n423), .A2(new_n422), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT35), .B1(new_n478), .B2(new_n472), .ZN(new_n479));
  AOI22_X1  g278(.A1(new_n420), .A2(new_n469), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(G113gat), .B(G141gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n481), .B(G197gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(KEYINPUT11), .B(G169gat), .ZN(new_n483));
  XOR2_X1   g282(.A(new_n482), .B(new_n483), .Z(new_n484));
  XNOR2_X1  g283(.A(new_n484), .B(KEYINPUT12), .ZN(new_n485));
  XNOR2_X1  g284(.A(G15gat), .B(G22gat), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT16), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(G1gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT88), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n486), .A2(new_n491), .A3(KEYINPUT16), .A4(new_n489), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(KEYINPUT89), .A2(G8gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(KEYINPUT89), .A2(G8gat), .ZN(new_n498));
  INV_X1    g297(.A(new_n496), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n493), .B(new_n494), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT17), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT15), .ZN(new_n503));
  OR2_X1    g302(.A1(G43gat), .A2(G50gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(G43gat), .A2(G50gat), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  AND2_X1   g306(.A1(KEYINPUT85), .A2(G36gat), .ZN(new_n508));
  NOR2_X1   g307(.A1(KEYINPUT85), .A2(G36gat), .ZN(new_n509));
  OAI21_X1  g308(.A(G29gat), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT14), .ZN(new_n511));
  OR3_X1    g310(.A1(new_n511), .A2(G29gat), .A3(G36gat), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n511), .B1(G29gat), .B2(G36gat), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n510), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n505), .A2(new_n503), .ZN(new_n515));
  AND2_X1   g314(.A1(KEYINPUT86), .A2(G43gat), .ZN(new_n516));
  NOR2_X1   g315(.A1(KEYINPUT86), .A2(G43gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(G50gat), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n507), .B1(new_n514), .B2(new_n520), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n506), .A2(new_n510), .A3(new_n513), .A4(new_n512), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT87), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n502), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT87), .A4(KEYINPUT17), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n501), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n523), .B1(new_n497), .B2(new_n500), .ZN(new_n528));
  NAND2_X1  g327(.A1(G229gat), .A2(G233gat), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NOR3_X1   g329(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n485), .B1(new_n531), .B2(KEYINPUT18), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n497), .A2(new_n500), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(new_n523), .ZN(new_n534));
  INV_X1    g333(.A(new_n528), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(new_n529), .B(KEYINPUT13), .Z(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n525), .A2(new_n526), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n533), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n540), .A2(KEYINPUT18), .A3(new_n535), .A4(new_n529), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n532), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT18), .ZN(new_n544));
  NOR4_X1   g343(.A1(new_n527), .A2(new_n544), .A3(new_n528), .A4(new_n530), .ZN(new_n545));
  INV_X1    g344(.A(new_n537), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n546), .B1(new_n534), .B2(new_n535), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT90), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n531), .A2(KEYINPUT18), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT90), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n538), .A2(new_n541), .A3(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n485), .B(KEYINPUT84), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n543), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G183gat), .B(G211gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT93), .ZN(new_n556));
  XNOR2_X1  g355(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(new_n204), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n556), .B(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(G71gat), .B(G78gat), .Z(new_n561));
  AOI21_X1  g360(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n562));
  INV_X1    g361(.A(G57gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(G64gat), .ZN(new_n564));
  INV_X1    g363(.A(G64gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(G57gat), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n562), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT91), .ZN(new_n568));
  OAI211_X1 g367(.A(KEYINPUT92), .B(new_n561), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT92), .ZN(new_n570));
  NAND2_X1  g369(.A1(G71gat), .A2(G78gat), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT9), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n565), .A2(G57gat), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n563), .A2(G64gat), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n570), .B1(new_n576), .B2(KEYINPUT91), .ZN(new_n577));
  XNOR2_X1  g376(.A(G71gat), .B(G78gat), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n578), .B1(new_n567), .B2(KEYINPUT92), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n569), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n580), .A2(KEYINPUT21), .ZN(new_n581));
  NAND2_X1  g380(.A1(G231gat), .A2(G233gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n583), .A2(new_n226), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n226), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n501), .B1(KEYINPUT21), .B2(new_n580), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n584), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n587), .B1(new_n584), .B2(new_n585), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n560), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n590), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n592), .A2(new_n588), .A3(new_n559), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G232gat), .A2(G233gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT94), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n596), .A2(KEYINPUT41), .ZN(new_n597));
  XNOR2_X1  g396(.A(G134gat), .B(G162gat), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n597), .B(new_n598), .Z(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G190gat), .B(G218gat), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT97), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n602), .A2(KEYINPUT98), .ZN(new_n603));
  OR2_X1    g402(.A1(KEYINPUT95), .A2(G92gat), .ZN(new_n604));
  INV_X1    g403(.A(G85gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(KEYINPUT95), .A2(G92gat), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G85gat), .A2(G92gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT7), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT7), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n610), .A2(G85gat), .A3(G92gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(G99gat), .ZN(new_n613));
  INV_X1    g412(.A(G106gat), .ZN(new_n614));
  OAI21_X1  g413(.A(KEYINPUT8), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n607), .A2(new_n612), .A3(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(G99gat), .B(G106gat), .Z(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n617), .A2(new_n607), .A3(new_n612), .A4(new_n615), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n603), .B1(new_n539), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n602), .A2(KEYINPUT98), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n621), .A2(new_n521), .A3(new_n522), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n596), .A2(KEYINPUT41), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT96), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n625), .A2(KEYINPUT96), .A3(new_n626), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AND3_X1   g430(.A1(new_n623), .A2(new_n624), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n624), .B1(new_n623), .B2(new_n631), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n600), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n630), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT96), .B1(new_n625), .B2(new_n626), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n621), .B1(new_n525), .B2(new_n526), .ZN(new_n638));
  OAI211_X1 g437(.A(KEYINPUT98), .B(new_n602), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n624), .A3(new_n631), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n639), .A2(new_n599), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n634), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n594), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(G230gat), .A2(G233gat), .ZN(new_n645));
  XOR2_X1   g444(.A(KEYINPUT100), .B(KEYINPUT10), .Z(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT99), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n616), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n580), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n621), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n622), .A2(new_n580), .A3(new_n649), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n647), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n580), .A2(new_n621), .A3(KEYINPUT10), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(KEYINPUT101), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT101), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n580), .A2(new_n621), .A3(new_n656), .A4(KEYINPUT10), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n645), .B1(new_n653), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n645), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n651), .A2(new_n652), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(G120gat), .B(G148gat), .Z(new_n662));
  XOR2_X1   g461(.A(G176gat), .B(G204gat), .Z(new_n663));
  XOR2_X1   g462(.A(new_n662), .B(new_n663), .Z(new_n664));
  NAND3_X1  g463(.A1(new_n659), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n665), .A2(KEYINPUT102), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT102), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n659), .A2(new_n667), .A3(new_n661), .A4(new_n664), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT104), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n659), .A2(new_n661), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n664), .B(KEYINPUT103), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n670), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  AOI211_X1 g473(.A(KEYINPUT104), .B(new_n672), .C1(new_n659), .C2(new_n661), .ZN(new_n675));
  OAI22_X1  g474(.A1(new_n666), .A2(new_n669), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n644), .A2(new_n677), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n480), .A2(new_n554), .A3(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n422), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g481(.A1(new_n679), .A2(new_n418), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n683), .A2(KEYINPUT105), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(KEYINPUT105), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n684), .A2(G8gat), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT42), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT16), .B(G8gat), .ZN(new_n688));
  OR3_X1    g487(.A1(new_n683), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n688), .B1(new_n684), .B2(new_n685), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n686), .B(new_n689), .C1(new_n690), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g490(.A(new_n679), .ZN(new_n692));
  INV_X1    g491(.A(new_n460), .ZN(new_n693));
  OR3_X1    g492(.A1(new_n692), .A2(G15gat), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n462), .A2(new_n468), .ZN(new_n695));
  OAI21_X1  g494(.A(G15gat), .B1(new_n692), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(G1326gat));
  NAND2_X1  g496(.A1(new_n679), .A2(new_n397), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT43), .B(G22gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  NAND2_X1  g499(.A1(new_n420), .A2(new_n469), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n477), .A2(new_n479), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n642), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n594), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n704), .A2(new_n676), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n554), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(G29gat), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n708), .A2(new_n709), .A3(new_n680), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT45), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n701), .A2(new_n702), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n712), .A2(KEYINPUT44), .A3(new_n643), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n714), .B1(new_n480), .B2(new_n642), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n707), .ZN(new_n717));
  OAI21_X1  g516(.A(G29gat), .B1(new_n717), .B2(new_n422), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n711), .A2(new_n718), .ZN(G1328gat));
  OR2_X1    g518(.A1(new_n508), .A2(new_n509), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n720), .B1(new_n717), .B2(new_n423), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n552), .A2(new_n553), .ZN(new_n722));
  INV_X1    g521(.A(new_n543), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR4_X1   g523(.A1(new_n706), .A2(new_n423), .A3(new_n720), .A4(new_n642), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n712), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n726), .B(KEYINPUT46), .Z(new_n727));
  NAND2_X1  g526(.A1(new_n721), .A2(new_n727), .ZN(G1329gat));
  INV_X1    g527(.A(new_n695), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n716), .A2(new_n729), .A3(new_n707), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n730), .A2(KEYINPUT106), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(KEYINPUT106), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n731), .A2(new_n732), .A3(new_n518), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n708), .A2(new_n460), .A3(new_n518), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT47), .ZN(new_n735));
  INV_X1    g534(.A(new_n518), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n730), .A2(new_n736), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n737), .A2(new_n734), .ZN(new_n738));
  OAI22_X1  g537(.A1(new_n733), .A2(new_n735), .B1(KEYINPUT47), .B2(new_n738), .ZN(G1330gat));
  NAND2_X1  g538(.A1(new_n397), .A2(G50gat), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n708), .A2(new_n397), .ZN(new_n741));
  OAI22_X1  g540(.A1(new_n717), .A2(new_n740), .B1(new_n741), .B2(G50gat), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT48), .ZN(G1331gat));
  AND4_X1   g542(.A1(new_n712), .A2(new_n554), .A3(new_n644), .A4(new_n676), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n680), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n418), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT49), .B(G64gat), .Z(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n747), .B2(new_n749), .ZN(G1333gat));
  NAND2_X1  g549(.A1(new_n744), .A2(new_n729), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n693), .A2(G71gat), .ZN(new_n752));
  AOI22_X1  g551(.A1(new_n751), .A2(G71gat), .B1(new_n744), .B2(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1334gat));
  NAND2_X1  g554(.A1(new_n744), .A2(new_n397), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g556(.A1(new_n594), .A2(new_n554), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n758), .A2(new_n677), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n716), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(G85gat), .B1(new_n760), .B2(new_n422), .ZN(new_n761));
  INV_X1    g560(.A(new_n758), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT51), .B1(new_n703), .B2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT51), .ZN(new_n764));
  NOR4_X1   g563(.A1(new_n480), .A2(new_n764), .A3(new_n642), .A4(new_n758), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n680), .A2(new_n605), .A3(new_n676), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n761), .B1(new_n766), .B2(new_n767), .ZN(G1336gat));
  NAND4_X1  g567(.A1(new_n713), .A2(new_n715), .A3(new_n418), .A4(new_n759), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n604), .A2(new_n606), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n423), .A2(new_n677), .A3(G92gat), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n774), .B1(new_n766), .B2(new_n776), .ZN(new_n777));
  OAI211_X1 g576(.A(KEYINPUT110), .B(new_n775), .C1(new_n763), .C2(new_n765), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n773), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n712), .A2(new_n643), .A3(new_n762), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n764), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT109), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n703), .A2(KEYINPUT51), .A3(new_n762), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n763), .A2(KEYINPUT109), .ZN(new_n785));
  XOR2_X1   g584(.A(new_n775), .B(KEYINPUT108), .Z(new_n786));
  NAND3_X1  g585(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n772), .B1(new_n787), .B2(new_n771), .ZN(new_n788));
  OAI21_X1  g587(.A(KEYINPUT111), .B1(new_n779), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT52), .B1(new_n769), .B2(new_n770), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n781), .A2(new_n783), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT110), .B1(new_n791), .B2(new_n775), .ZN(new_n792));
  INV_X1    g591(.A(new_n778), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n790), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n769), .A2(new_n770), .ZN(new_n796));
  AOI211_X1 g595(.A(new_n782), .B(KEYINPUT51), .C1(new_n703), .C2(new_n762), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n797), .B1(new_n766), .B2(new_n782), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n796), .B1(new_n798), .B2(new_n786), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n794), .B(new_n795), .C1(new_n799), .C2(new_n772), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n789), .A2(new_n800), .ZN(G1337gat));
  OAI21_X1  g600(.A(G99gat), .B1(new_n760), .B2(new_n695), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n460), .A2(new_n613), .A3(new_n676), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(KEYINPUT112), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n766), .B2(new_n804), .ZN(G1338gat));
  NAND3_X1  g604(.A1(new_n716), .A2(new_n397), .A3(new_n759), .ZN(new_n806));
  XNOR2_X1  g605(.A(KEYINPUT113), .B(G106gat), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n396), .A2(new_n677), .A3(G106gat), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT53), .B1(new_n791), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  AOI22_X1  g610(.A1(new_n798), .A2(new_n809), .B1(new_n806), .B2(new_n807), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n811), .B1(new_n812), .B2(new_n813), .ZN(G1339gat));
  NAND3_X1  g613(.A1(new_n644), .A2(new_n554), .A3(new_n677), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT10), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n561), .B1(new_n576), .B2(new_n570), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT92), .B1(new_n567), .B2(new_n568), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n817), .B1(new_n820), .B2(new_n569), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n656), .B1(new_n821), .B2(new_n621), .ZN(new_n822));
  INV_X1    g621(.A(new_n657), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AND4_X1   g623(.A1(new_n580), .A2(new_n619), .A3(new_n620), .A4(new_n649), .ZN(new_n825));
  AOI22_X1  g624(.A1(new_n580), .A2(new_n649), .B1(new_n619), .B2(new_n620), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n646), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n816), .B1(new_n828), .B2(new_n645), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n824), .A2(new_n827), .A3(new_n660), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n824), .A2(new_n827), .A3(KEYINPUT114), .A4(new_n660), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n829), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n816), .B(new_n645), .C1(new_n653), .C2(new_n658), .ZN(new_n835));
  INV_X1    g634(.A(new_n664), .ZN(new_n836));
  AND3_X1   g635(.A1(new_n835), .A2(KEYINPUT55), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n665), .A2(KEYINPUT102), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n668), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n835), .A2(new_n836), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT55), .B1(new_n834), .B2(new_n842), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n534), .A2(new_n535), .A3(new_n546), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n529), .B1(new_n540), .B2(new_n535), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n484), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n846), .B1(new_n532), .B2(new_n542), .ZN(new_n847));
  NOR4_X1   g646(.A1(new_n841), .A2(new_n843), .A3(new_n642), .A4(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n847), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n676), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n842), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT55), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI22_X1  g652(.A1(new_n834), .A2(new_n837), .B1(new_n839), .B2(new_n668), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n850), .B1(new_n855), .B2(new_n554), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n848), .B1(new_n856), .B2(new_n642), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n815), .B1(new_n857), .B2(new_n704), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n858), .A2(new_n680), .ZN(new_n859));
  AND4_X1   g658(.A1(new_n396), .A2(new_n859), .A3(new_n423), .A4(new_n460), .ZN(new_n860));
  AOI21_X1  g659(.A(G113gat), .B1(new_n860), .B2(new_n724), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n858), .A2(new_n396), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n422), .A2(new_n418), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(new_n693), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n724), .A2(G113gat), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n861), .B1(new_n865), .B2(new_n866), .ZN(G1340gat));
  AOI21_X1  g666(.A(G120gat), .B1(new_n860), .B2(new_n676), .ZN(new_n868));
  INV_X1    g667(.A(new_n864), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n693), .A2(new_n677), .A3(new_n236), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(G1341gat));
  NAND3_X1  g670(.A1(new_n860), .A2(new_n226), .A3(new_n704), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n864), .A2(new_n693), .A3(new_n594), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n226), .B2(new_n873), .ZN(G1342gat));
  NAND3_X1  g673(.A1(new_n860), .A2(new_n230), .A3(new_n643), .ZN(new_n875));
  XOR2_X1   g674(.A(new_n875), .B(KEYINPUT56), .Z(new_n876));
  NOR3_X1   g675(.A1(new_n864), .A2(new_n693), .A3(new_n642), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(new_n227), .B2(new_n877), .ZN(G1343gat));
  NOR2_X1   g677(.A1(new_n729), .A2(new_n396), .ZN(new_n879));
  AND3_X1   g678(.A1(new_n859), .A2(new_n423), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n207), .A3(new_n724), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n695), .A2(new_n863), .ZN(new_n882));
  XOR2_X1   g681(.A(KEYINPUT115), .B(KEYINPUT57), .Z(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n884), .B1(new_n858), .B2(new_n397), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n397), .A2(KEYINPUT57), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT116), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n887), .B1(new_n841), .B2(new_n843), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n853), .A2(new_n854), .A3(KEYINPUT116), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(new_n724), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n643), .B1(new_n890), .B2(new_n850), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n594), .B1(new_n891), .B2(new_n848), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n886), .B1(new_n892), .B2(new_n815), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT117), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n885), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n815), .ZN(new_n896));
  INV_X1    g695(.A(new_n848), .ZN(new_n897));
  INV_X1    g696(.A(new_n850), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n554), .B1(new_n855), .B2(new_n887), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n899), .B2(new_n889), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n897), .B1(new_n900), .B2(new_n643), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n896), .B1(new_n901), .B2(new_n594), .ZN(new_n902));
  OAI21_X1  g701(.A(KEYINPUT117), .B1(new_n902), .B2(new_n886), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n882), .B1(new_n895), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n207), .B1(new_n904), .B2(new_n724), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n881), .B1(new_n905), .B2(KEYINPUT118), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT118), .ZN(new_n907));
  AOI211_X1 g706(.A(new_n907), .B(new_n207), .C1(new_n904), .C2(new_n724), .ZN(new_n908));
  OAI21_X1  g707(.A(KEYINPUT58), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT119), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n881), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT58), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n912), .B1(new_n881), .B2(new_n910), .ZN(new_n913));
  OR3_X1    g712(.A1(new_n905), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n909), .A2(new_n914), .ZN(G1344gat));
  NAND3_X1  g714(.A1(new_n880), .A2(new_n208), .A3(new_n676), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT59), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT120), .ZN(new_n918));
  INV_X1    g717(.A(new_n855), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(new_n643), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n855), .A2(KEYINPUT120), .A3(new_n642), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n920), .A2(new_n921), .A3(new_n847), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n594), .B1(new_n922), .B2(new_n891), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(new_n815), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT57), .B1(new_n924), .B2(new_n397), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n858), .A2(new_n397), .A3(new_n884), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n927), .A2(new_n695), .A3(new_n676), .A4(new_n863), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n917), .B1(new_n928), .B2(G148gat), .ZN(new_n929));
  AOI211_X1 g728(.A(KEYINPUT59), .B(new_n208), .C1(new_n904), .C2(new_n676), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n916), .B1(new_n929), .B2(new_n930), .ZN(G1345gat));
  NAND3_X1  g730(.A1(new_n880), .A2(new_n204), .A3(new_n704), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n904), .A2(new_n704), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n933), .B2(new_n204), .ZN(G1346gat));
  NAND3_X1  g733(.A1(new_n880), .A2(new_n205), .A3(new_n643), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n904), .A2(new_n643), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n935), .B1(new_n936), .B2(new_n205), .ZN(G1347gat));
  AND2_X1   g736(.A1(new_n858), .A2(new_n422), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n472), .A2(new_n423), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(G169gat), .B1(new_n941), .B2(new_n724), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n422), .A2(new_n418), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n943), .A2(new_n693), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT121), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n862), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n554), .A2(new_n314), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n942), .B1(new_n946), .B2(new_n947), .ZN(G1348gat));
  INV_X1    g747(.A(new_n946), .ZN(new_n949));
  OAI21_X1  g748(.A(G176gat), .B1(new_n949), .B2(new_n677), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n941), .A2(new_n315), .A3(new_n676), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(G1349gat));
  OAI21_X1  g751(.A(G183gat), .B1(new_n949), .B2(new_n594), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n941), .A2(new_n305), .A3(new_n704), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT60), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n956), .A2(KEYINPUT122), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n955), .B(new_n957), .ZN(G1350gat));
  NAND3_X1  g757(.A1(new_n941), .A2(new_n306), .A3(new_n643), .ZN(new_n959));
  OAI21_X1  g758(.A(G190gat), .B1(new_n949), .B2(new_n642), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n960), .A2(KEYINPUT61), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n960), .A2(KEYINPUT61), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(G1351gat));
  NAND2_X1  g762(.A1(new_n879), .A2(new_n418), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT123), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(new_n938), .ZN(new_n966));
  OR3_X1    g765(.A1(new_n966), .A2(G197gat), .A3(new_n554), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n729), .A2(new_n943), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n927), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g768(.A(KEYINPUT124), .B1(new_n969), .B2(new_n554), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(G197gat), .ZN(new_n971));
  NOR3_X1   g770(.A1(new_n969), .A2(KEYINPUT124), .A3(new_n554), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n967), .B1(new_n971), .B2(new_n972), .ZN(G1352gat));
  NOR3_X1   g772(.A1(new_n966), .A2(G204gat), .A3(new_n677), .ZN(new_n974));
  NAND2_X1  g773(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g775(.A(G204gat), .B1(new_n969), .B2(new_n677), .ZN(new_n977));
  XOR2_X1   g776(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n978));
  OAI211_X1 g777(.A(new_n976), .B(new_n977), .C1(new_n974), .C2(new_n978), .ZN(G1353gat));
  NOR3_X1   g778(.A1(new_n966), .A2(G211gat), .A3(new_n594), .ZN(new_n980));
  OAI211_X1 g779(.A(new_n704), .B(new_n968), .C1(new_n925), .C2(new_n926), .ZN(new_n981));
  AOI21_X1  g780(.A(KEYINPUT63), .B1(new_n981), .B2(G211gat), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT126), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OR2_X1    g783(.A1(new_n982), .A2(new_n983), .ZN(new_n985));
  AND3_X1   g784(.A1(new_n981), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n984), .B1(new_n985), .B2(new_n986), .ZN(G1354gat));
  OAI21_X1  g786(.A(G218gat), .B1(new_n969), .B2(new_n642), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n643), .A2(new_n330), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n988), .B1(new_n966), .B2(new_n989), .ZN(G1355gat));
endmodule


