

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X2 U549 ( .A(n652), .ZN(n633) );
  NAND2_X2 U550 ( .A1(n698), .A2(n591), .ZN(n652) );
  NOR2_X1 U551 ( .A1(G651), .A2(G543), .ZN(n781) );
  NAND2_X1 U552 ( .A1(n652), .A2(G1341), .ZN(n513) );
  XOR2_X1 U553 ( .A(KEYINPUT78), .B(n610), .Z(n514) );
  XOR2_X1 U554 ( .A(KEYINPUT76), .B(n596), .Z(n515) );
  NOR2_X1 U555 ( .A1(n986), .A2(n606), .ZN(n607) );
  INV_X1 U556 ( .A(KEYINPUT102), .ZN(n649) );
  AND2_X2 U557 ( .A1(n520), .A2(G2104), .ZN(n882) );
  XNOR2_X1 U558 ( .A(n614), .B(KEYINPUT15), .ZN(n1000) );
  NOR2_X1 U559 ( .A1(n524), .A2(n523), .ZN(G160) );
  NOR2_X1 U560 ( .A1(G2104), .A2(G2105), .ZN(n516) );
  XOR2_X2 U561 ( .A(KEYINPUT17), .B(n516), .Z(n881) );
  NAND2_X1 U562 ( .A1(n881), .A2(G137), .ZN(n519) );
  INV_X1 U563 ( .A(G2105), .ZN(n520) );
  NAND2_X1 U564 ( .A1(G101), .A2(n882), .ZN(n517) );
  XOR2_X1 U565 ( .A(KEYINPUT23), .B(n517), .Z(n518) );
  NAND2_X1 U566 ( .A1(n519), .A2(n518), .ZN(n524) );
  AND2_X1 U567 ( .A1(G2104), .A2(G2105), .ZN(n877) );
  NAND2_X1 U568 ( .A1(G113), .A2(n877), .ZN(n522) );
  NOR2_X1 U569 ( .A1(G2104), .A2(n520), .ZN(n878) );
  NAND2_X1 U570 ( .A1(G125), .A2(n878), .ZN(n521) );
  NAND2_X1 U571 ( .A1(n522), .A2(n521), .ZN(n523) );
  INV_X1 U572 ( .A(G651), .ZN(n534) );
  NOR2_X1 U573 ( .A1(G543), .A2(n534), .ZN(n525) );
  XOR2_X1 U574 ( .A(KEYINPUT1), .B(n525), .Z(n775) );
  XOR2_X1 U575 ( .A(G543), .B(KEYINPUT0), .Z(n535) );
  NOR2_X1 U576 ( .A1(G651), .A2(n535), .ZN(n526) );
  XOR2_X2 U577 ( .A(KEYINPUT65), .B(n526), .Z(n776) );
  NAND2_X1 U578 ( .A1(G49), .A2(n776), .ZN(n528) );
  NAND2_X1 U579 ( .A1(G74), .A2(G651), .ZN(n527) );
  NAND2_X1 U580 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U581 ( .A1(n775), .A2(n529), .ZN(n532) );
  NAND2_X1 U582 ( .A1(G87), .A2(n535), .ZN(n530) );
  XOR2_X1 U583 ( .A(KEYINPUT85), .B(n530), .Z(n531) );
  NAND2_X1 U584 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U585 ( .A(KEYINPUT86), .B(n533), .ZN(G288) );
  NOR2_X1 U586 ( .A1(n535), .A2(n534), .ZN(n780) );
  NAND2_X1 U587 ( .A1(G78), .A2(n780), .ZN(n537) );
  NAND2_X1 U588 ( .A1(G91), .A2(n781), .ZN(n536) );
  NAND2_X1 U589 ( .A1(n537), .A2(n536), .ZN(n540) );
  NAND2_X1 U590 ( .A1(n775), .A2(G65), .ZN(n538) );
  XOR2_X1 U591 ( .A(KEYINPUT70), .B(n538), .Z(n539) );
  NOR2_X1 U592 ( .A1(n540), .A2(n539), .ZN(n542) );
  NAND2_X1 U593 ( .A1(n776), .A2(G53), .ZN(n541) );
  NAND2_X1 U594 ( .A1(n542), .A2(n541), .ZN(G299) );
  NAND2_X1 U595 ( .A1(n775), .A2(G64), .ZN(n543) );
  XNOR2_X1 U596 ( .A(KEYINPUT67), .B(n543), .ZN(n552) );
  NAND2_X1 U597 ( .A1(n781), .A2(G90), .ZN(n544) );
  XNOR2_X1 U598 ( .A(n544), .B(KEYINPUT68), .ZN(n546) );
  NAND2_X1 U599 ( .A1(G77), .A2(n780), .ZN(n545) );
  NAND2_X1 U600 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U601 ( .A(KEYINPUT69), .B(n547), .Z(n548) );
  XNOR2_X1 U602 ( .A(n548), .B(KEYINPUT9), .ZN(n550) );
  NAND2_X1 U603 ( .A1(G52), .A2(n776), .ZN(n549) );
  NAND2_X1 U604 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U605 ( .A1(n552), .A2(n551), .ZN(G171) );
  NAND2_X1 U606 ( .A1(G63), .A2(n775), .ZN(n554) );
  NAND2_X1 U607 ( .A1(G51), .A2(n776), .ZN(n553) );
  NAND2_X1 U608 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U609 ( .A(KEYINPUT6), .B(n555), .ZN(n562) );
  NAND2_X1 U610 ( .A1(n781), .A2(G89), .ZN(n556) );
  XNOR2_X1 U611 ( .A(n556), .B(KEYINPUT4), .ZN(n558) );
  NAND2_X1 U612 ( .A1(G76), .A2(n780), .ZN(n557) );
  NAND2_X1 U613 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U614 ( .A(KEYINPUT79), .B(n559), .ZN(n560) );
  XNOR2_X1 U615 ( .A(KEYINPUT5), .B(n560), .ZN(n561) );
  NOR2_X1 U616 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U617 ( .A(KEYINPUT7), .B(n563), .Z(G168) );
  XOR2_X1 U618 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U619 ( .A1(G75), .A2(n780), .ZN(n565) );
  NAND2_X1 U620 ( .A1(G88), .A2(n781), .ZN(n564) );
  NAND2_X1 U621 ( .A1(n565), .A2(n564), .ZN(n568) );
  NAND2_X1 U622 ( .A1(G50), .A2(n776), .ZN(n566) );
  XNOR2_X1 U623 ( .A(KEYINPUT87), .B(n566), .ZN(n567) );
  NOR2_X1 U624 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U625 ( .A1(n775), .A2(G62), .ZN(n569) );
  NAND2_X1 U626 ( .A1(n570), .A2(n569), .ZN(G303) );
  INV_X1 U627 ( .A(G303), .ZN(G166) );
  NAND2_X1 U628 ( .A1(G61), .A2(n775), .ZN(n572) );
  NAND2_X1 U629 ( .A1(G48), .A2(n776), .ZN(n571) );
  NAND2_X1 U630 ( .A1(n572), .A2(n571), .ZN(n575) );
  NAND2_X1 U631 ( .A1(n780), .A2(G73), .ZN(n573) );
  XOR2_X1 U632 ( .A(KEYINPUT2), .B(n573), .Z(n574) );
  NOR2_X1 U633 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U634 ( .A1(n781), .A2(G86), .ZN(n576) );
  NAND2_X1 U635 ( .A1(n577), .A2(n576), .ZN(G305) );
  NAND2_X1 U636 ( .A1(G47), .A2(n776), .ZN(n579) );
  NAND2_X1 U637 ( .A1(G85), .A2(n781), .ZN(n578) );
  NAND2_X1 U638 ( .A1(n579), .A2(n578), .ZN(n582) );
  NAND2_X1 U639 ( .A1(G72), .A2(n780), .ZN(n580) );
  XOR2_X1 U640 ( .A(KEYINPUT66), .B(n580), .Z(n581) );
  NOR2_X1 U641 ( .A1(n582), .A2(n581), .ZN(n584) );
  NAND2_X1 U642 ( .A1(n775), .A2(G60), .ZN(n583) );
  NAND2_X1 U643 ( .A1(n584), .A2(n583), .ZN(G290) );
  NAND2_X1 U644 ( .A1(G138), .A2(n881), .ZN(n590) );
  AND2_X1 U645 ( .A1(G102), .A2(n882), .ZN(n588) );
  NAND2_X1 U646 ( .A1(G114), .A2(n877), .ZN(n586) );
  NAND2_X1 U647 ( .A1(G126), .A2(n878), .ZN(n585) );
  NAND2_X1 U648 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U649 ( .A1(n588), .A2(n587), .ZN(n589) );
  AND2_X1 U650 ( .A1(n590), .A2(n589), .ZN(G164) );
  NOR2_X2 U651 ( .A1(G164), .A2(G1384), .ZN(n698) );
  AND2_X1 U652 ( .A1(G160), .A2(G40), .ZN(n591) );
  NAND2_X1 U653 ( .A1(G8), .A2(n652), .ZN(n692) );
  NOR2_X1 U654 ( .A1(G1976), .A2(G288), .ZN(n673) );
  NAND2_X1 U655 ( .A1(n673), .A2(KEYINPUT33), .ZN(n592) );
  NOR2_X1 U656 ( .A1(n692), .A2(n592), .ZN(n681) );
  XOR2_X1 U657 ( .A(KEYINPUT14), .B(KEYINPUT75), .Z(n594) );
  NAND2_X1 U658 ( .A1(G56), .A2(n775), .ZN(n593) );
  XNOR2_X1 U659 ( .A(n594), .B(n593), .ZN(n595) );
  XNOR2_X1 U660 ( .A(KEYINPUT74), .B(n595), .ZN(n603) );
  NAND2_X1 U661 ( .A1(n776), .A2(G43), .ZN(n596) );
  NAND2_X1 U662 ( .A1(n781), .A2(G81), .ZN(n597) );
  XNOR2_X1 U663 ( .A(n597), .B(KEYINPUT12), .ZN(n599) );
  NAND2_X1 U664 ( .A1(G68), .A2(n780), .ZN(n598) );
  NAND2_X1 U665 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U666 ( .A(KEYINPUT13), .B(n600), .Z(n601) );
  NOR2_X1 U667 ( .A1(n515), .A2(n601), .ZN(n602) );
  NAND2_X1 U668 ( .A1(n603), .A2(n602), .ZN(n986) );
  XOR2_X1 U669 ( .A(G1996), .B(KEYINPUT99), .Z(n942) );
  NAND2_X1 U670 ( .A1(n633), .A2(n942), .ZN(n604) );
  XNOR2_X1 U671 ( .A(n604), .B(KEYINPUT26), .ZN(n605) );
  NAND2_X1 U672 ( .A1(n605), .A2(n513), .ZN(n606) );
  XOR2_X1 U673 ( .A(KEYINPUT64), .B(n607), .Z(n620) );
  NAND2_X1 U674 ( .A1(G92), .A2(n781), .ZN(n613) );
  NAND2_X1 U675 ( .A1(G66), .A2(n775), .ZN(n609) );
  NAND2_X1 U676 ( .A1(G54), .A2(n776), .ZN(n608) );
  NAND2_X1 U677 ( .A1(n609), .A2(n608), .ZN(n611) );
  NAND2_X1 U678 ( .A1(n780), .A2(G79), .ZN(n610) );
  NOR2_X1 U679 ( .A1(n611), .A2(n514), .ZN(n612) );
  NAND2_X1 U680 ( .A1(n613), .A2(n612), .ZN(n614) );
  INV_X1 U681 ( .A(n1000), .ZN(n752) );
  OR2_X1 U682 ( .A1(n620), .A2(n752), .ZN(n619) );
  NAND2_X1 U683 ( .A1(G1348), .A2(n652), .ZN(n616) );
  NAND2_X1 U684 ( .A1(G2067), .A2(n633), .ZN(n615) );
  NAND2_X1 U685 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U686 ( .A(n617), .B(KEYINPUT100), .ZN(n618) );
  NAND2_X1 U687 ( .A1(n619), .A2(n618), .ZN(n622) );
  NAND2_X1 U688 ( .A1(n620), .A2(n752), .ZN(n621) );
  NAND2_X1 U689 ( .A1(n622), .A2(n621), .ZN(n627) );
  INV_X1 U690 ( .A(G299), .ZN(n999) );
  NAND2_X1 U691 ( .A1(n633), .A2(G2072), .ZN(n623) );
  XNOR2_X1 U692 ( .A(n623), .B(KEYINPUT27), .ZN(n625) );
  AND2_X1 U693 ( .A1(G1956), .A2(n652), .ZN(n624) );
  NOR2_X1 U694 ( .A1(n625), .A2(n624), .ZN(n628) );
  NAND2_X1 U695 ( .A1(n999), .A2(n628), .ZN(n626) );
  NAND2_X1 U696 ( .A1(n627), .A2(n626), .ZN(n631) );
  NOR2_X1 U697 ( .A1(n999), .A2(n628), .ZN(n629) );
  XOR2_X1 U698 ( .A(n629), .B(KEYINPUT28), .Z(n630) );
  NAND2_X1 U699 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U700 ( .A(n632), .B(KEYINPUT29), .ZN(n638) );
  NAND2_X1 U701 ( .A1(n652), .A2(G1961), .ZN(n635) );
  XOR2_X1 U702 ( .A(KEYINPUT25), .B(G2078), .Z(n936) );
  NAND2_X1 U703 ( .A1(n633), .A2(n936), .ZN(n634) );
  NAND2_X1 U704 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U705 ( .A(n636), .B(KEYINPUT98), .Z(n642) );
  AND2_X1 U706 ( .A1(G171), .A2(n642), .ZN(n637) );
  NOR2_X1 U707 ( .A1(n638), .A2(n637), .ZN(n648) );
  NOR2_X1 U708 ( .A1(G1966), .A2(n692), .ZN(n664) );
  NOR2_X1 U709 ( .A1(G2084), .A2(n652), .ZN(n666) );
  NOR2_X1 U710 ( .A1(n664), .A2(n666), .ZN(n639) );
  NAND2_X1 U711 ( .A1(G8), .A2(n639), .ZN(n640) );
  XNOR2_X1 U712 ( .A(KEYINPUT30), .B(n640), .ZN(n641) );
  NOR2_X1 U713 ( .A1(G168), .A2(n641), .ZN(n644) );
  NOR2_X1 U714 ( .A1(G171), .A2(n642), .ZN(n643) );
  NOR2_X1 U715 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U716 ( .A(n645), .B(KEYINPUT101), .Z(n646) );
  XNOR2_X1 U717 ( .A(KEYINPUT31), .B(n646), .ZN(n647) );
  NOR2_X1 U718 ( .A1(n648), .A2(n647), .ZN(n650) );
  XNOR2_X1 U719 ( .A(n650), .B(n649), .ZN(n663) );
  NAND2_X1 U720 ( .A1(n663), .A2(G286), .ZN(n660) );
  INV_X1 U721 ( .A(G8), .ZN(n658) );
  NOR2_X1 U722 ( .A1(G1971), .A2(n692), .ZN(n651) );
  XNOR2_X1 U723 ( .A(KEYINPUT103), .B(n651), .ZN(n656) );
  NOR2_X1 U724 ( .A1(G2090), .A2(n652), .ZN(n653) );
  XNOR2_X1 U725 ( .A(KEYINPUT104), .B(n653), .ZN(n654) );
  NOR2_X1 U726 ( .A1(G166), .A2(n654), .ZN(n655) );
  NAND2_X1 U727 ( .A1(n656), .A2(n655), .ZN(n657) );
  OR2_X1 U728 ( .A1(n658), .A2(n657), .ZN(n659) );
  AND2_X1 U729 ( .A1(n660), .A2(n659), .ZN(n662) );
  XOR2_X1 U730 ( .A(KEYINPUT32), .B(KEYINPUT105), .Z(n661) );
  XNOR2_X1 U731 ( .A(n662), .B(n661), .ZN(n683) );
  INV_X1 U732 ( .A(n663), .ZN(n665) );
  NOR2_X1 U733 ( .A1(n665), .A2(n664), .ZN(n668) );
  NAND2_X1 U734 ( .A1(G8), .A2(n666), .ZN(n667) );
  NAND2_X1 U735 ( .A1(n668), .A2(n667), .ZN(n684) );
  NAND2_X1 U736 ( .A1(G1976), .A2(G288), .ZN(n991) );
  AND2_X1 U737 ( .A1(n684), .A2(n991), .ZN(n670) );
  INV_X1 U738 ( .A(n692), .ZN(n669) );
  AND2_X1 U739 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U740 ( .A1(n683), .A2(n671), .ZN(n678) );
  INV_X1 U741 ( .A(n991), .ZN(n675) );
  NOR2_X1 U742 ( .A1(G1971), .A2(G303), .ZN(n672) );
  NOR2_X1 U743 ( .A1(n673), .A2(n672), .ZN(n992) );
  XNOR2_X1 U744 ( .A(KEYINPUT106), .B(n992), .ZN(n674) );
  OR2_X1 U745 ( .A1(n675), .A2(n674), .ZN(n676) );
  OR2_X1 U746 ( .A1(n692), .A2(n676), .ZN(n677) );
  NAND2_X1 U747 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U748 ( .A1(n679), .A2(KEYINPUT33), .ZN(n680) );
  NOR2_X1 U749 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U750 ( .A(G1981), .B(G305), .Z(n983) );
  AND2_X1 U751 ( .A1(n682), .A2(n983), .ZN(n696) );
  NAND2_X1 U752 ( .A1(n684), .A2(n683), .ZN(n687) );
  NOR2_X1 U753 ( .A1(G2090), .A2(G303), .ZN(n685) );
  NAND2_X1 U754 ( .A1(G8), .A2(n685), .ZN(n686) );
  AND2_X1 U755 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U756 ( .A(KEYINPUT107), .B(n688), .ZN(n689) );
  NAND2_X1 U757 ( .A1(n689), .A2(n692), .ZN(n694) );
  NOR2_X1 U758 ( .A1(G1981), .A2(G305), .ZN(n690) );
  XOR2_X1 U759 ( .A(n690), .B(KEYINPUT24), .Z(n691) );
  OR2_X1 U760 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U761 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U762 ( .A1(n696), .A2(n695), .ZN(n730) );
  NAND2_X1 U763 ( .A1(G160), .A2(G40), .ZN(n697) );
  NOR2_X1 U764 ( .A1(n698), .A2(n697), .ZN(n742) );
  XOR2_X1 U765 ( .A(KEYINPUT36), .B(KEYINPUT94), .Z(n710) );
  NAND2_X1 U766 ( .A1(G140), .A2(n881), .ZN(n700) );
  NAND2_X1 U767 ( .A1(G104), .A2(n882), .ZN(n699) );
  NAND2_X1 U768 ( .A1(n700), .A2(n699), .ZN(n702) );
  XOR2_X1 U769 ( .A(KEYINPUT34), .B(KEYINPUT93), .Z(n701) );
  XNOR2_X1 U770 ( .A(n702), .B(n701), .ZN(n707) );
  NAND2_X1 U771 ( .A1(G116), .A2(n877), .ZN(n704) );
  NAND2_X1 U772 ( .A1(G128), .A2(n878), .ZN(n703) );
  NAND2_X1 U773 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U774 ( .A(KEYINPUT35), .B(n705), .Z(n706) );
  NOR2_X1 U775 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U776 ( .A(n708), .B(KEYINPUT95), .ZN(n709) );
  XNOR2_X1 U777 ( .A(n710), .B(n709), .ZN(n872) );
  XNOR2_X1 U778 ( .A(G2067), .B(KEYINPUT37), .ZN(n740) );
  NOR2_X1 U779 ( .A1(n872), .A2(n740), .ZN(n975) );
  NAND2_X1 U780 ( .A1(n742), .A2(n975), .ZN(n738) );
  NAND2_X1 U781 ( .A1(G131), .A2(n881), .ZN(n712) );
  NAND2_X1 U782 ( .A1(G95), .A2(n882), .ZN(n711) );
  NAND2_X1 U783 ( .A1(n712), .A2(n711), .ZN(n716) );
  NAND2_X1 U784 ( .A1(G107), .A2(n877), .ZN(n714) );
  NAND2_X1 U785 ( .A1(G119), .A2(n878), .ZN(n713) );
  NAND2_X1 U786 ( .A1(n714), .A2(n713), .ZN(n715) );
  OR2_X1 U787 ( .A1(n716), .A2(n715), .ZN(n888) );
  NAND2_X1 U788 ( .A1(G1991), .A2(n888), .ZN(n726) );
  NAND2_X1 U789 ( .A1(G129), .A2(n878), .ZN(n723) );
  NAND2_X1 U790 ( .A1(G141), .A2(n881), .ZN(n718) );
  NAND2_X1 U791 ( .A1(G117), .A2(n877), .ZN(n717) );
  NAND2_X1 U792 ( .A1(n718), .A2(n717), .ZN(n721) );
  NAND2_X1 U793 ( .A1(n882), .A2(G105), .ZN(n719) );
  XOR2_X1 U794 ( .A(KEYINPUT38), .B(n719), .Z(n720) );
  NOR2_X1 U795 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U796 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U797 ( .A(n724), .B(KEYINPUT96), .ZN(n861) );
  NAND2_X1 U798 ( .A1(G1996), .A2(n861), .ZN(n725) );
  NAND2_X1 U799 ( .A1(n726), .A2(n725), .ZN(n962) );
  NAND2_X1 U800 ( .A1(n962), .A2(n742), .ZN(n727) );
  XNOR2_X1 U801 ( .A(n727), .B(KEYINPUT97), .ZN(n735) );
  INV_X1 U802 ( .A(n735), .ZN(n728) );
  NAND2_X1 U803 ( .A1(n738), .A2(n728), .ZN(n729) );
  NOR2_X1 U804 ( .A1(n730), .A2(n729), .ZN(n732) );
  XNOR2_X1 U805 ( .A(G1986), .B(G290), .ZN(n1004) );
  NAND2_X1 U806 ( .A1(n1004), .A2(n742), .ZN(n731) );
  NAND2_X1 U807 ( .A1(n732), .A2(n731), .ZN(n745) );
  NOR2_X1 U808 ( .A1(G1996), .A2(n861), .ZN(n955) );
  NOR2_X1 U809 ( .A1(G1986), .A2(G290), .ZN(n733) );
  NOR2_X1 U810 ( .A1(G1991), .A2(n888), .ZN(n958) );
  NOR2_X1 U811 ( .A1(n733), .A2(n958), .ZN(n734) );
  NOR2_X1 U812 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U813 ( .A1(n955), .A2(n736), .ZN(n737) );
  XNOR2_X1 U814 ( .A(n737), .B(KEYINPUT39), .ZN(n739) );
  NAND2_X1 U815 ( .A1(n739), .A2(n738), .ZN(n741) );
  NAND2_X1 U816 ( .A1(n872), .A2(n740), .ZN(n972) );
  NAND2_X1 U817 ( .A1(n741), .A2(n972), .ZN(n743) );
  NAND2_X1 U818 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U819 ( .A1(n745), .A2(n744), .ZN(n747) );
  XNOR2_X1 U820 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n746) );
  XNOR2_X1 U821 ( .A(n747), .B(n746), .ZN(G329) );
  AND2_X1 U822 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U823 ( .A(G120), .ZN(G236) );
  INV_X1 U824 ( .A(G69), .ZN(G235) );
  INV_X1 U825 ( .A(G108), .ZN(G238) );
  NAND2_X1 U826 ( .A1(G7), .A2(G661), .ZN(n749) );
  XNOR2_X1 U827 ( .A(n749), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U828 ( .A(G223), .ZN(n816) );
  NAND2_X1 U829 ( .A1(n816), .A2(G567), .ZN(n750) );
  XNOR2_X1 U830 ( .A(n750), .B(KEYINPUT11), .ZN(n751) );
  XNOR2_X1 U831 ( .A(KEYINPUT73), .B(n751), .ZN(G234) );
  XNOR2_X1 U832 ( .A(G860), .B(KEYINPUT77), .ZN(n758) );
  OR2_X1 U833 ( .A1(n986), .A2(n758), .ZN(G153) );
  INV_X1 U834 ( .A(G171), .ZN(G301) );
  NAND2_X1 U835 ( .A1(G868), .A2(G301), .ZN(n754) );
  INV_X1 U836 ( .A(G868), .ZN(n755) );
  NAND2_X1 U837 ( .A1(n752), .A2(n755), .ZN(n753) );
  NAND2_X1 U838 ( .A1(n754), .A2(n753), .ZN(G284) );
  NOR2_X1 U839 ( .A1(G286), .A2(n755), .ZN(n757) );
  NOR2_X1 U840 ( .A1(G868), .A2(G299), .ZN(n756) );
  NOR2_X1 U841 ( .A1(n757), .A2(n756), .ZN(G297) );
  NAND2_X1 U842 ( .A1(n758), .A2(G559), .ZN(n759) );
  NAND2_X1 U843 ( .A1(n759), .A2(n1000), .ZN(n760) );
  XNOR2_X1 U844 ( .A(n760), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U845 ( .A1(G868), .A2(n986), .ZN(n763) );
  NAND2_X1 U846 ( .A1(n1000), .A2(G868), .ZN(n761) );
  NOR2_X1 U847 ( .A1(G559), .A2(n761), .ZN(n762) );
  NOR2_X1 U848 ( .A1(n763), .A2(n762), .ZN(G282) );
  NAND2_X1 U849 ( .A1(G111), .A2(n877), .ZN(n770) );
  NAND2_X1 U850 ( .A1(G135), .A2(n881), .ZN(n765) );
  NAND2_X1 U851 ( .A1(G99), .A2(n882), .ZN(n764) );
  NAND2_X1 U852 ( .A1(n765), .A2(n764), .ZN(n768) );
  NAND2_X1 U853 ( .A1(n878), .A2(G123), .ZN(n766) );
  XOR2_X1 U854 ( .A(KEYINPUT18), .B(n766), .Z(n767) );
  NOR2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U856 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U857 ( .A(n771), .B(KEYINPUT80), .ZN(n960) );
  XOR2_X1 U858 ( .A(n960), .B(G2096), .Z(n773) );
  XNOR2_X1 U859 ( .A(G2100), .B(KEYINPUT81), .ZN(n772) );
  NAND2_X1 U860 ( .A1(n773), .A2(n772), .ZN(G156) );
  NAND2_X1 U861 ( .A1(G559), .A2(n1000), .ZN(n774) );
  XNOR2_X1 U862 ( .A(n986), .B(n774), .ZN(n797) );
  NOR2_X1 U863 ( .A1(G860), .A2(n797), .ZN(n788) );
  NAND2_X1 U864 ( .A1(G67), .A2(n775), .ZN(n778) );
  NAND2_X1 U865 ( .A1(G55), .A2(n776), .ZN(n777) );
  NAND2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U867 ( .A(KEYINPUT84), .B(n779), .ZN(n786) );
  NAND2_X1 U868 ( .A1(G80), .A2(n780), .ZN(n783) );
  NAND2_X1 U869 ( .A1(G93), .A2(n781), .ZN(n782) );
  NAND2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n784) );
  XOR2_X1 U871 ( .A(KEYINPUT83), .B(n784), .Z(n785) );
  NOR2_X1 U872 ( .A1(n786), .A2(n785), .ZN(n791) );
  XNOR2_X1 U873 ( .A(n791), .B(KEYINPUT82), .ZN(n787) );
  XNOR2_X1 U874 ( .A(n788), .B(n787), .ZN(G145) );
  NOR2_X1 U875 ( .A1(G868), .A2(n791), .ZN(n789) );
  XNOR2_X1 U876 ( .A(n789), .B(KEYINPUT89), .ZN(n800) );
  XNOR2_X1 U877 ( .A(n999), .B(KEYINPUT19), .ZN(n790) );
  XNOR2_X1 U878 ( .A(n790), .B(KEYINPUT88), .ZN(n792) );
  XOR2_X1 U879 ( .A(n792), .B(n791), .Z(n794) );
  XNOR2_X1 U880 ( .A(G166), .B(G288), .ZN(n793) );
  XNOR2_X1 U881 ( .A(n794), .B(n793), .ZN(n795) );
  XNOR2_X1 U882 ( .A(n795), .B(G290), .ZN(n796) );
  XNOR2_X1 U883 ( .A(n796), .B(G305), .ZN(n894) );
  XOR2_X1 U884 ( .A(n894), .B(n797), .Z(n798) );
  NAND2_X1 U885 ( .A1(G868), .A2(n798), .ZN(n799) );
  NAND2_X1 U886 ( .A1(n800), .A2(n799), .ZN(G295) );
  NAND2_X1 U887 ( .A1(G2078), .A2(G2084), .ZN(n801) );
  XOR2_X1 U888 ( .A(KEYINPUT20), .B(n801), .Z(n802) );
  NAND2_X1 U889 ( .A1(G2090), .A2(n802), .ZN(n803) );
  XNOR2_X1 U890 ( .A(KEYINPUT21), .B(n803), .ZN(n804) );
  NAND2_X1 U891 ( .A1(n804), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U892 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U893 ( .A(KEYINPUT72), .B(G82), .Z(G220) );
  XNOR2_X1 U894 ( .A(KEYINPUT71), .B(G132), .ZN(G219) );
  NOR2_X1 U895 ( .A1(G235), .A2(G236), .ZN(n805) );
  XOR2_X1 U896 ( .A(KEYINPUT90), .B(n805), .Z(n806) );
  NOR2_X1 U897 ( .A1(G238), .A2(n806), .ZN(n807) );
  NAND2_X1 U898 ( .A1(G57), .A2(n807), .ZN(n820) );
  NAND2_X1 U899 ( .A1(G567), .A2(n820), .ZN(n808) );
  XOR2_X1 U900 ( .A(KEYINPUT91), .B(n808), .Z(n813) );
  NOR2_X1 U901 ( .A1(G220), .A2(G219), .ZN(n809) );
  XOR2_X1 U902 ( .A(KEYINPUT22), .B(n809), .Z(n810) );
  NOR2_X1 U903 ( .A1(G218), .A2(n810), .ZN(n811) );
  NAND2_X1 U904 ( .A1(G96), .A2(n811), .ZN(n821) );
  NAND2_X1 U905 ( .A1(G2106), .A2(n821), .ZN(n812) );
  NAND2_X1 U906 ( .A1(n813), .A2(n812), .ZN(n832) );
  NAND2_X1 U907 ( .A1(G661), .A2(G483), .ZN(n814) );
  NOR2_X1 U908 ( .A1(n832), .A2(n814), .ZN(n819) );
  NAND2_X1 U909 ( .A1(G36), .A2(n819), .ZN(n815) );
  XNOR2_X1 U910 ( .A(n815), .B(KEYINPUT92), .ZN(G176) );
  NAND2_X1 U911 ( .A1(G2106), .A2(n816), .ZN(G217) );
  AND2_X1 U912 ( .A1(G15), .A2(G2), .ZN(n817) );
  NAND2_X1 U913 ( .A1(G661), .A2(n817), .ZN(G259) );
  NAND2_X1 U914 ( .A1(G3), .A2(G1), .ZN(n818) );
  NAND2_X1 U915 ( .A1(n819), .A2(n818), .ZN(G188) );
  INV_X1 U917 ( .A(G96), .ZN(G221) );
  NOR2_X1 U918 ( .A1(n821), .A2(n820), .ZN(G325) );
  INV_X1 U919 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U920 ( .A(G1348), .B(G2454), .ZN(n822) );
  XNOR2_X1 U921 ( .A(n822), .B(G2430), .ZN(n823) );
  XNOR2_X1 U922 ( .A(n823), .B(G1341), .ZN(n829) );
  XOR2_X1 U923 ( .A(G2443), .B(G2427), .Z(n825) );
  XNOR2_X1 U924 ( .A(G2438), .B(G2446), .ZN(n824) );
  XNOR2_X1 U925 ( .A(n825), .B(n824), .ZN(n827) );
  XOR2_X1 U926 ( .A(G2451), .B(G2435), .Z(n826) );
  XNOR2_X1 U927 ( .A(n827), .B(n826), .ZN(n828) );
  XNOR2_X1 U928 ( .A(n829), .B(n828), .ZN(n830) );
  NAND2_X1 U929 ( .A1(n830), .A2(G14), .ZN(n831) );
  XNOR2_X1 U930 ( .A(KEYINPUT109), .B(n831), .ZN(n903) );
  XNOR2_X1 U931 ( .A(n903), .B(KEYINPUT110), .ZN(G401) );
  XNOR2_X1 U932 ( .A(KEYINPUT111), .B(n832), .ZN(G319) );
  XOR2_X1 U933 ( .A(G2096), .B(KEYINPUT43), .Z(n834) );
  XNOR2_X1 U934 ( .A(G2090), .B(KEYINPUT112), .ZN(n833) );
  XNOR2_X1 U935 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U936 ( .A(n835), .B(G2678), .Z(n837) );
  XNOR2_X1 U937 ( .A(G2067), .B(G2072), .ZN(n836) );
  XNOR2_X1 U938 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U939 ( .A(KEYINPUT42), .B(G2100), .Z(n839) );
  XNOR2_X1 U940 ( .A(G2078), .B(G2084), .ZN(n838) );
  XNOR2_X1 U941 ( .A(n839), .B(n838), .ZN(n840) );
  XNOR2_X1 U942 ( .A(n841), .B(n840), .ZN(G227) );
  XOR2_X1 U943 ( .A(G1981), .B(G1961), .Z(n843) );
  XNOR2_X1 U944 ( .A(G1996), .B(G1986), .ZN(n842) );
  XNOR2_X1 U945 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U946 ( .A(G1976), .B(G1971), .Z(n845) );
  XNOR2_X1 U947 ( .A(G1966), .B(G1956), .ZN(n844) );
  XNOR2_X1 U948 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U949 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U950 ( .A(G2474), .B(KEYINPUT41), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n849), .B(n848), .ZN(n851) );
  XOR2_X1 U952 ( .A(G1991), .B(KEYINPUT113), .Z(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(G229) );
  NAND2_X1 U954 ( .A1(n878), .A2(G124), .ZN(n852) );
  XNOR2_X1 U955 ( .A(n852), .B(KEYINPUT44), .ZN(n854) );
  NAND2_X1 U956 ( .A1(G136), .A2(n881), .ZN(n853) );
  NAND2_X1 U957 ( .A1(n854), .A2(n853), .ZN(n855) );
  XOR2_X1 U958 ( .A(KEYINPUT114), .B(n855), .Z(n857) );
  NAND2_X1 U959 ( .A1(n882), .A2(G100), .ZN(n856) );
  NAND2_X1 U960 ( .A1(n857), .A2(n856), .ZN(n860) );
  NAND2_X1 U961 ( .A1(G112), .A2(n877), .ZN(n858) );
  XNOR2_X1 U962 ( .A(KEYINPUT115), .B(n858), .ZN(n859) );
  NOR2_X1 U963 ( .A1(n860), .A2(n859), .ZN(G162) );
  XNOR2_X1 U964 ( .A(n861), .B(n960), .ZN(n876) );
  XOR2_X1 U965 ( .A(KEYINPUT48), .B(KEYINPUT116), .Z(n863) );
  XNOR2_X1 U966 ( .A(G162), .B(KEYINPUT46), .ZN(n862) );
  XNOR2_X1 U967 ( .A(n863), .B(n862), .ZN(n871) );
  NAND2_X1 U968 ( .A1(G139), .A2(n881), .ZN(n865) );
  NAND2_X1 U969 ( .A1(G103), .A2(n882), .ZN(n864) );
  NAND2_X1 U970 ( .A1(n865), .A2(n864), .ZN(n870) );
  NAND2_X1 U971 ( .A1(G115), .A2(n877), .ZN(n867) );
  NAND2_X1 U972 ( .A1(G127), .A2(n878), .ZN(n866) );
  NAND2_X1 U973 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U974 ( .A(KEYINPUT47), .B(n868), .Z(n869) );
  NOR2_X1 U975 ( .A1(n870), .A2(n869), .ZN(n965) );
  XOR2_X1 U976 ( .A(n871), .B(n965), .Z(n874) );
  XNOR2_X1 U977 ( .A(G164), .B(n872), .ZN(n873) );
  XNOR2_X1 U978 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U979 ( .A(n876), .B(n875), .ZN(n892) );
  NAND2_X1 U980 ( .A1(G118), .A2(n877), .ZN(n880) );
  NAND2_X1 U981 ( .A1(G130), .A2(n878), .ZN(n879) );
  NAND2_X1 U982 ( .A1(n880), .A2(n879), .ZN(n887) );
  NAND2_X1 U983 ( .A1(G142), .A2(n881), .ZN(n884) );
  NAND2_X1 U984 ( .A1(G106), .A2(n882), .ZN(n883) );
  NAND2_X1 U985 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U986 ( .A(n885), .B(KEYINPUT45), .Z(n886) );
  NOR2_X1 U987 ( .A1(n887), .A2(n886), .ZN(n889) );
  XNOR2_X1 U988 ( .A(n889), .B(n888), .ZN(n890) );
  XOR2_X1 U989 ( .A(G160), .B(n890), .Z(n891) );
  XNOR2_X1 U990 ( .A(n892), .B(n891), .ZN(n893) );
  NOR2_X1 U991 ( .A1(G37), .A2(n893), .ZN(G395) );
  XOR2_X1 U992 ( .A(KEYINPUT117), .B(n894), .Z(n896) );
  XNOR2_X1 U993 ( .A(G171), .B(G286), .ZN(n895) );
  XNOR2_X1 U994 ( .A(n896), .B(n895), .ZN(n898) );
  XNOR2_X1 U995 ( .A(n986), .B(n1000), .ZN(n897) );
  XNOR2_X1 U996 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U997 ( .A1(G37), .A2(n899), .ZN(G397) );
  NOR2_X1 U998 ( .A1(G227), .A2(G229), .ZN(n900) );
  XOR2_X1 U999 ( .A(KEYINPUT49), .B(n900), .Z(n901) );
  NAND2_X1 U1000 ( .A1(G319), .A2(n901), .ZN(n902) );
  NOR2_X1 U1001 ( .A1(n903), .A2(n902), .ZN(n905) );
  NOR2_X1 U1002 ( .A1(G395), .A2(G397), .ZN(n904) );
  NAND2_X1 U1003 ( .A1(n905), .A2(n904), .ZN(G225) );
  INV_X1 U1004 ( .A(G225), .ZN(G308) );
  INV_X1 U1005 ( .A(G57), .ZN(G237) );
  XOR2_X1 U1006 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n916) );
  XNOR2_X1 U1007 ( .A(G1341), .B(G19), .ZN(n907) );
  XNOR2_X1 U1008 ( .A(G6), .B(G1981), .ZN(n906) );
  NOR2_X1 U1009 ( .A1(n907), .A2(n906), .ZN(n914) );
  XOR2_X1 U1010 ( .A(KEYINPUT124), .B(G4), .Z(n909) );
  XNOR2_X1 U1011 ( .A(G1348), .B(KEYINPUT59), .ZN(n908) );
  XNOR2_X1 U1012 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1013 ( .A(KEYINPUT123), .B(n910), .Z(n912) );
  XNOR2_X1 U1014 ( .A(G1956), .B(G20), .ZN(n911) );
  NOR2_X1 U1015 ( .A1(n912), .A2(n911), .ZN(n913) );
  NAND2_X1 U1016 ( .A1(n914), .A2(n913), .ZN(n915) );
  XNOR2_X1 U1017 ( .A(n916), .B(n915), .ZN(n919) );
  XNOR2_X1 U1018 ( .A(G1966), .B(KEYINPUT126), .ZN(n917) );
  XNOR2_X1 U1019 ( .A(G21), .B(n917), .ZN(n918) );
  NOR2_X1 U1020 ( .A1(n919), .A2(n918), .ZN(n927) );
  XNOR2_X1 U1021 ( .A(G1986), .B(G24), .ZN(n921) );
  XNOR2_X1 U1022 ( .A(G22), .B(G1971), .ZN(n920) );
  NOR2_X1 U1023 ( .A1(n921), .A2(n920), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(G1976), .B(KEYINPUT127), .ZN(n922) );
  XNOR2_X1 U1025 ( .A(n922), .B(G23), .ZN(n923) );
  NAND2_X1 U1026 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1027 ( .A(KEYINPUT58), .B(n925), .Z(n926) );
  NAND2_X1 U1028 ( .A1(n927), .A2(n926), .ZN(n929) );
  XNOR2_X1 U1029 ( .A(G5), .B(G1961), .ZN(n928) );
  NOR2_X1 U1030 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1031 ( .A(KEYINPUT61), .B(n930), .Z(n931) );
  NOR2_X1 U1032 ( .A1(G16), .A2(n931), .ZN(n1012) );
  XNOR2_X1 U1033 ( .A(G2084), .B(G34), .ZN(n932) );
  XNOR2_X1 U1034 ( .A(n932), .B(KEYINPUT54), .ZN(n947) );
  XNOR2_X1 U1035 ( .A(G2067), .B(G26), .ZN(n934) );
  XNOR2_X1 U1036 ( .A(G1991), .B(G25), .ZN(n933) );
  NOR2_X1 U1037 ( .A1(n934), .A2(n933), .ZN(n941) );
  XOR2_X1 U1038 ( .A(G2072), .B(G33), .Z(n935) );
  NAND2_X1 U1039 ( .A1(n935), .A2(G28), .ZN(n939) );
  XOR2_X1 U1040 ( .A(G27), .B(n936), .Z(n937) );
  XNOR2_X1 U1041 ( .A(KEYINPUT121), .B(n937), .ZN(n938) );
  NOR2_X1 U1042 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1043 ( .A1(n941), .A2(n940), .ZN(n944) );
  XNOR2_X1 U1044 ( .A(G32), .B(n942), .ZN(n943) );
  NOR2_X1 U1045 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1046 ( .A(n945), .B(KEYINPUT53), .ZN(n946) );
  NOR2_X1 U1047 ( .A1(n947), .A2(n946), .ZN(n950) );
  XOR2_X1 U1048 ( .A(G2090), .B(KEYINPUT120), .Z(n948) );
  XNOR2_X1 U1049 ( .A(G35), .B(n948), .ZN(n949) );
  NAND2_X1 U1050 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1051 ( .A(KEYINPUT55), .B(n951), .Z(n952) );
  INV_X1 U1052 ( .A(G29), .ZN(n980) );
  NAND2_X1 U1053 ( .A1(n952), .A2(n980), .ZN(n953) );
  NAND2_X1 U1054 ( .A1(G11), .A2(n953), .ZN(n982) );
  XNOR2_X1 U1055 ( .A(KEYINPUT119), .B(KEYINPUT52), .ZN(n977) );
  XOR2_X1 U1056 ( .A(G2090), .B(G162), .Z(n954) );
  NOR2_X1 U1057 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1058 ( .A(KEYINPUT51), .B(n956), .Z(n964) );
  XOR2_X1 U1059 ( .A(G160), .B(G2084), .Z(n957) );
  NOR2_X1 U1060 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1061 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1062 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1063 ( .A1(n964), .A2(n963), .ZN(n971) );
  XOR2_X1 U1064 ( .A(G2072), .B(n965), .Z(n967) );
  XOR2_X1 U1065 ( .A(G164), .B(G2078), .Z(n966) );
  NOR2_X1 U1066 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1067 ( .A(KEYINPUT118), .B(n968), .Z(n969) );
  XNOR2_X1 U1068 ( .A(KEYINPUT50), .B(n969), .ZN(n970) );
  NOR2_X1 U1069 ( .A1(n971), .A2(n970), .ZN(n973) );
  NAND2_X1 U1070 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1072 ( .A(n977), .B(n976), .ZN(n978) );
  NOR2_X1 U1073 ( .A1(n978), .A2(KEYINPUT55), .ZN(n979) );
  NOR2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n1010) );
  XNOR2_X1 U1076 ( .A(G16), .B(KEYINPUT56), .ZN(n1008) );
  XNOR2_X1 U1077 ( .A(G1966), .B(G168), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1079 ( .A(n985), .B(KEYINPUT57), .ZN(n990) );
  XNOR2_X1 U1080 ( .A(G301), .B(G1961), .ZN(n988) );
  XNOR2_X1 U1081 ( .A(n986), .B(G1341), .ZN(n987) );
  NOR2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n998) );
  NAND2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n995) );
  INV_X1 U1085 ( .A(G1971), .ZN(n993) );
  NOR2_X1 U1086 ( .A1(G166), .A2(n993), .ZN(n994) );
  NOR2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1088 ( .A(KEYINPUT122), .B(n996), .Z(n997) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n1006) );
  XNOR2_X1 U1090 ( .A(n999), .B(G1956), .ZN(n1002) );
  XNOR2_X1 U1091 ( .A(n1000), .B(G1348), .ZN(n1001) );
  NAND2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NOR2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1098 ( .A(n1013), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1099 ( .A(G311), .ZN(G150) );
endmodule

