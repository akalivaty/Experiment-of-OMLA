//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 0 0 0 1 0 0 0 1 0 1 0 0 0 1 0 1 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n785, new_n786,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n865, new_n866, new_n867, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n986, new_n987, new_n988;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT32), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT67), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT66), .ZN(new_n205));
  INV_X1    g004(.A(G169gat), .ZN(new_n206));
  INV_X1    g005(.A(G176gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n209));
  AND3_X1   g008(.A1(new_n208), .A2(KEYINPUT23), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n211), .B(KEYINPUT65), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n204), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n211), .B(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n208), .A2(KEYINPUT23), .A3(new_n209), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT67), .ZN(new_n217));
  NOR2_X1   g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT25), .B1(new_n218), .B2(KEYINPUT23), .ZN(new_n219));
  NAND3_X1  g018(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n219), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n213), .A2(new_n217), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT25), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n218), .A2(KEYINPUT23), .ZN(new_n227));
  XOR2_X1   g026(.A(KEYINPUT64), .B(G169gat), .Z(new_n228));
  NAND2_X1  g027(.A1(new_n207), .A2(KEYINPUT23), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n227), .B(new_n211), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  AND2_X1   g029(.A1(new_n223), .A2(new_n220), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n226), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n225), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G183gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT27), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT27), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G183gat), .ZN(new_n237));
  INV_X1    g036(.A(G190gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT28), .ZN(new_n240));
  OR2_X1    g039(.A1(new_n240), .A2(KEYINPUT68), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(KEYINPUT68), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n239), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT27), .B(G183gat), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n244), .A2(KEYINPUT68), .A3(new_n240), .A4(new_n238), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n243), .A2(new_n245), .A3(new_n222), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT26), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n208), .A2(new_n247), .A3(new_n209), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n208), .A2(KEYINPUT69), .A3(new_n247), .A4(new_n209), .ZN(new_n251));
  OAI21_X1  g050(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n250), .A2(new_n211), .A3(new_n251), .A4(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n246), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n233), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT75), .ZN(new_n256));
  INV_X1    g055(.A(G134gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(G127gat), .ZN(new_n258));
  INV_X1    g057(.A(G127gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(G134gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G113gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n263), .A2(G120gat), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT74), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(G120gat), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G120gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n268), .A2(G113gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT74), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n262), .B1(new_n267), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT72), .B1(new_n264), .B2(new_n269), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n268), .A2(G113gat), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT72), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n274), .A2(new_n266), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n273), .A2(new_n261), .A3(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(KEYINPUT70), .B1(new_n259), .B2(G134gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n279), .A2(new_n257), .A3(G127gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n259), .A2(KEYINPUT71), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT71), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(G127gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n282), .A2(new_n284), .A3(G134gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  AND3_X1   g085(.A1(new_n277), .A2(KEYINPUT73), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT73), .B1(new_n277), .B2(new_n286), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n272), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n255), .A2(new_n256), .A3(new_n289), .ZN(new_n290));
  AOI22_X1  g089(.A1(new_n225), .A2(new_n232), .B1(new_n246), .B2(new_n253), .ZN(new_n291));
  XNOR2_X1  g090(.A(G113gat), .B(G120gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n261), .B1(new_n292), .B2(new_n275), .ZN(new_n293));
  INV_X1    g092(.A(new_n276), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n286), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT73), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n277), .A2(KEYINPUT73), .A3(new_n286), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n271), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT75), .B1(new_n291), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n291), .A2(new_n299), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n290), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G227gat), .A2(G233gat), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n203), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT33), .B1(new_n302), .B2(new_n304), .ZN(new_n306));
  XOR2_X1   g105(.A(G15gat), .B(G43gat), .Z(new_n307));
  XNOR2_X1  g106(.A(G71gat), .B(G99gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NOR3_X1   g109(.A1(new_n305), .A2(new_n306), .A3(new_n310), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n290), .B(new_n303), .C1(new_n300), .C2(new_n301), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n312), .B(KEYINPUT34), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n302), .A2(new_n304), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n309), .B(KEYINPUT76), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT33), .ZN(new_n316));
  OR2_X1    g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AND3_X1   g116(.A1(new_n314), .A2(KEYINPUT32), .A3(new_n317), .ZN(new_n318));
  NOR3_X1   g117(.A1(new_n311), .A2(new_n313), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT34), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n312), .B(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n314), .A2(KEYINPUT32), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n314), .A2(new_n316), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n322), .A2(new_n323), .A3(new_n309), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n305), .A2(new_n317), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n321), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n319), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT77), .B(KEYINPUT36), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT77), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n330), .B(KEYINPUT36), .C1(new_n319), .C2(new_n326), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G197gat), .B(G204gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(G211gat), .A2(G218gat), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT78), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT22), .ZN(new_n336));
  AND3_X1   g135(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n335), .B1(new_n334), .B2(new_n336), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n333), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G211gat), .B(G218gat), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT79), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n333), .B(new_n340), .C1(new_n337), .C2(new_n338), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n339), .A2(KEYINPUT79), .A3(new_n341), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G141gat), .B(G148gat), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G155gat), .A2(G162gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT2), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT82), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT82), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n350), .A2(new_n353), .A3(KEYINPUT2), .ZN(new_n354));
  XNOR2_X1  g153(.A(G155gat), .B(G162gat), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n349), .A2(new_n352), .A3(new_n354), .A4(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(G155gat), .A2(G162gat), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n350), .B1(new_n357), .B2(KEYINPUT81), .ZN(new_n358));
  OR2_X1    g157(.A1(new_n350), .A2(KEYINPUT81), .ZN(new_n359));
  INV_X1    g158(.A(new_n351), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n358), .B(new_n359), .C1(new_n360), .C2(new_n348), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT3), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n356), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT29), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n347), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n356), .A2(new_n361), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT29), .B1(new_n342), .B2(new_n344), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n367), .B1(new_n368), .B2(KEYINPUT3), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(G228gat), .A2(G233gat), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n371), .B1(new_n347), .B2(new_n365), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n367), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n345), .A2(new_n364), .A3(new_n346), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n375), .B1(new_n376), .B2(new_n362), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(G22gat), .B1(new_n372), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n370), .A2(new_n371), .ZN(new_n380));
  INV_X1    g179(.A(G22gat), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n380), .B(new_n381), .C1(new_n377), .C2(new_n374), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G78gat), .B(G106gat), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n379), .A2(new_n382), .A3(new_n384), .ZN(new_n387));
  XOR2_X1   g186(.A(KEYINPUT31), .B(G50gat), .Z(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n386), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n389), .B1(new_n386), .B2(new_n387), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(G225gat), .A2(G233gat), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n297), .A2(new_n298), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n375), .B1(new_n395), .B2(new_n272), .ZN(new_n396));
  AOI211_X1 g195(.A(new_n367), .B(new_n271), .C1(new_n297), .C2(new_n298), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n394), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT85), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI211_X1 g199(.A(KEYINPUT85), .B(new_n394), .C1(new_n396), .C2(new_n397), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n400), .A2(KEYINPUT5), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT83), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n367), .A2(KEYINPUT3), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n363), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n403), .B1(new_n299), .B2(new_n405), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n356), .A2(new_n361), .A3(new_n362), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n362), .B1(new_n356), .B2(new_n361), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n289), .A2(new_n409), .A3(KEYINPUT83), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n375), .B(new_n272), .C1(new_n287), .C2(new_n288), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT4), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT4), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n395), .A2(new_n414), .A3(new_n375), .A4(new_n272), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n411), .A2(new_n393), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(KEYINPUT84), .A2(KEYINPUT5), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n406), .A2(new_n410), .B1(new_n413), .B2(new_n415), .ZN(new_n420));
  INV_X1    g219(.A(new_n418), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(new_n393), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n402), .A2(new_n419), .A3(new_n422), .ZN(new_n423));
  XOR2_X1   g222(.A(G1gat), .B(G29gat), .Z(new_n424));
  XNOR2_X1  g223(.A(G57gat), .B(G85gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT86), .B(KEYINPUT0), .ZN(new_n427));
  XOR2_X1   g226(.A(new_n426), .B(new_n427), .Z(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n423), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT6), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n402), .A2(new_n419), .A3(new_n428), .A4(new_n422), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n402), .A2(new_n419), .A3(new_n422), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT87), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n434), .A2(new_n435), .A3(KEYINPUT6), .A4(new_n428), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT87), .B1(new_n432), .B2(new_n431), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n433), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(G226gat), .ZN(new_n439));
  INV_X1    g238(.A(G233gat), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n255), .A2(KEYINPUT80), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n441), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n443), .B1(new_n291), .B2(KEYINPUT29), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT80), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n445), .B1(new_n291), .B2(new_n443), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n442), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n347), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n255), .A2(new_n441), .ZN(new_n449));
  INV_X1    g248(.A(new_n347), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n444), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(KEYINPUT90), .B(KEYINPUT37), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n448), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(G8gat), .B(G36gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(G64gat), .B(G92gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n455), .B(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT37), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n459), .B1(new_n448), .B2(new_n451), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT38), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n457), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n448), .A2(new_n451), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n450), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n444), .A2(new_n449), .A3(new_n347), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(KEYINPUT37), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT38), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n466), .A2(new_n454), .A3(new_n467), .A4(new_n457), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n461), .A2(new_n463), .A3(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n438), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n411), .A2(new_n416), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT39), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n471), .A2(new_n472), .A3(new_n394), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n289), .A2(new_n367), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n474), .A2(new_n393), .A3(new_n412), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT89), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n474), .A2(KEYINPUT89), .A3(new_n393), .A4(new_n412), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n420), .A2(new_n393), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n429), .B(new_n473), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT40), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n477), .B(new_n478), .C1(new_n393), .C2(new_n420), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n484), .A2(KEYINPUT40), .A3(new_n429), .A4(new_n473), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n432), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT30), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n448), .A2(new_n487), .A3(new_n451), .A4(new_n462), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n463), .A2(KEYINPUT30), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n462), .B1(new_n448), .B2(new_n451), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT88), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT88), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n493), .B(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n486), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n392), .B1(new_n470), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n392), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(new_n491), .A3(new_n438), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n332), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT35), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n438), .A2(new_n500), .A3(new_n492), .A4(new_n494), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT91), .B1(new_n319), .B2(new_n326), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n313), .B1(new_n311), .B2(new_n318), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT91), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n324), .A2(new_n321), .A3(new_n325), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n502), .A2(new_n392), .A3(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n392), .A2(new_n438), .A3(new_n327), .A4(new_n491), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n508), .A2(KEYINPUT92), .B1(KEYINPUT35), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT92), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n511), .B1(new_n501), .B2(new_n507), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n499), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT16), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n514), .A2(G1gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(G15gat), .B(G22gat), .ZN(new_n516));
  MUX2_X1   g315(.A(G1gat), .B(new_n515), .S(new_n516), .Z(new_n517));
  XNOR2_X1  g316(.A(new_n517), .B(G8gat), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT15), .ZN(new_n519));
  XNOR2_X1  g318(.A(G43gat), .B(G50gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT94), .ZN(new_n521));
  OR2_X1    g320(.A1(G43gat), .A2(G50gat), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT94), .ZN(new_n523));
  NAND2_X1  g322(.A1(G43gat), .A2(G50gat), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n519), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n520), .A2(KEYINPUT15), .ZN(new_n528));
  NAND2_X1  g327(.A1(G29gat), .A2(G36gat), .ZN(new_n529));
  OAI21_X1  g328(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NOR3_X1   g330(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n527), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT95), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n526), .A2(new_n536), .A3(new_n533), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n536), .B1(new_n526), .B2(new_n533), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n535), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n540), .A2(KEYINPUT96), .A3(KEYINPUT17), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT17), .B1(new_n540), .B2(KEYINPUT96), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n518), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G229gat), .A2(G233gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n526), .A2(new_n533), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT95), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n547), .A2(new_n537), .B1(new_n527), .B2(new_n534), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n548), .A2(new_n518), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n544), .A2(new_n545), .A3(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT18), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G113gat), .B(G141gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT11), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(new_n206), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(G197gat), .ZN(new_n557));
  XOR2_X1   g356(.A(KEYINPUT93), .B(KEYINPUT12), .Z(new_n558));
  XOR2_X1   g357(.A(new_n557), .B(new_n558), .Z(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n544), .A2(KEYINPUT18), .A3(new_n545), .A4(new_n550), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n540), .B(new_n518), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n545), .B(KEYINPUT13), .Z(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n553), .A2(new_n560), .A3(new_n561), .A4(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n561), .A2(new_n565), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT17), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT96), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n569), .B1(new_n548), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(new_n541), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n549), .B1(new_n572), .B2(new_n518), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT18), .B1(new_n573), .B2(new_n545), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n559), .B1(new_n568), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT97), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g376(.A(KEYINPUT97), .B(new_n559), .C1(new_n568), .C2(new_n574), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n567), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n202), .B1(new_n513), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n501), .ZN(new_n581));
  INV_X1    g380(.A(new_n507), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(new_n582), .A3(KEYINPUT92), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n509), .A2(KEYINPUT35), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n583), .A2(new_n512), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n496), .A2(new_n498), .ZN(new_n586));
  INV_X1    g385(.A(new_n332), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n553), .A2(new_n561), .A3(new_n565), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT97), .B1(new_n590), .B2(new_n559), .ZN(new_n591));
  INV_X1    g390(.A(new_n578), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n566), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n589), .A2(KEYINPUT98), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n580), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G127gat), .B(G155gat), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT100), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(G64gat), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n600), .A2(G57gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT99), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT99), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n603), .B1(G57gat), .B2(new_n600), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n602), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G71gat), .B(G78gat), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n599), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n600), .A2(G57gat), .ZN(new_n608));
  OAI21_X1  g407(.A(KEYINPUT9), .B1(new_n608), .B2(new_n601), .ZN(new_n609));
  INV_X1    g408(.A(new_n606), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n613), .A2(KEYINPUT21), .ZN(new_n614));
  NAND2_X1  g413(.A1(G231gat), .A2(G233gat), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n596), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n616), .A2(new_n617), .A3(new_n596), .ZN(new_n620));
  XOR2_X1   g419(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  AND3_X1   g421(.A1(new_n619), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n622), .B1(new_n619), .B2(new_n620), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n518), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n626), .B1(KEYINPUT21), .B2(new_n613), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  NOR3_X1   g428(.A1(new_n623), .A2(new_n624), .A3(new_n627), .ZN(new_n630));
  XOR2_X1   g429(.A(G183gat), .B(G211gat), .Z(new_n631));
  OR3_X1    g430(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n631), .B1(new_n629), .B2(new_n630), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G99gat), .A2(G106gat), .ZN(new_n635));
  INV_X1    g434(.A(G85gat), .ZN(new_n636));
  INV_X1    g435(.A(G92gat), .ZN(new_n637));
  AOI22_X1  g436(.A1(KEYINPUT8), .A2(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G85gat), .A2(G92gat), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n639), .A2(KEYINPUT103), .A3(KEYINPUT7), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n640), .B1(KEYINPUT7), .B2(new_n639), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT103), .B1(new_n639), .B2(KEYINPUT7), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n638), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(G99gat), .B(G106gat), .ZN(new_n644));
  OR2_X1    g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n571), .B2(new_n541), .ZN(new_n648));
  NAND3_X1  g447(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n649));
  INV_X1    g448(.A(new_n647), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n649), .B1(new_n548), .B2(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G190gat), .B(G218gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT104), .ZN(new_n654));
  OAI21_X1  g453(.A(KEYINPUT105), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT105), .ZN(new_n656));
  INV_X1    g455(.A(new_n654), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n656), .B(new_n657), .C1(new_n648), .C2(new_n651), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n652), .A2(new_n654), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n655), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT101), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(G134gat), .B(G162gat), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n664), .B(KEYINPUT102), .Z(new_n665));
  INV_X1    g464(.A(new_n662), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n655), .A2(new_n658), .A3(new_n659), .A4(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n663), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n665), .B1(new_n663), .B2(new_n667), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(G120gat), .B(G148gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(G176gat), .B(G204gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n643), .A2(KEYINPUT106), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n675), .A2(new_n644), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n675), .A2(new_n644), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n613), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n647), .A2(new_n612), .ZN(new_n679));
  AOI21_X1  g478(.A(KEYINPUT10), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n647), .A2(KEYINPUT10), .A3(new_n613), .ZN(new_n681));
  INV_X1    g480(.A(G230gat), .ZN(new_n682));
  OAI22_X1  g481(.A1(new_n680), .A2(new_n681), .B1(new_n682), .B2(new_n440), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n682), .A2(new_n440), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n678), .A2(new_n679), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n674), .B1(new_n684), .B2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n686), .B(KEYINPUT107), .ZN(new_n689));
  INV_X1    g488(.A(new_n674), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n689), .A2(new_n683), .A3(new_n690), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n634), .A2(new_n671), .A3(new_n693), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n595), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n438), .A2(KEYINPUT108), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n438), .A2(KEYINPUT108), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g500(.A1(new_n492), .A2(new_n494), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n595), .A2(new_n702), .A3(new_n694), .ZN(new_n703));
  XNOR2_X1  g502(.A(KEYINPUT16), .B(G8gat), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n704), .B(KEYINPUT109), .Z(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n703), .A2(KEYINPUT42), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n695), .A2(new_n702), .A3(new_n705), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT42), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n709), .B1(new_n703), .B2(G8gat), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n707), .B1(new_n708), .B2(new_n710), .ZN(G1325gat));
  INV_X1    g510(.A(G15gat), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n502), .A2(new_n506), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n695), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n695), .A2(new_n332), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n715), .B1(new_n716), .B2(new_n712), .ZN(G1326gat));
  NAND2_X1  g516(.A1(new_n695), .A2(new_n497), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT43), .B(G22gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1327gat));
  NAND2_X1  g519(.A1(new_n634), .A2(new_n692), .ZN(new_n721));
  INV_X1    g520(.A(new_n670), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n668), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n698), .A2(G29gat), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n595), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT45), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n595), .A2(KEYINPUT45), .A3(new_n724), .A4(new_n725), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n513), .B2(new_n723), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n589), .A2(KEYINPUT44), .A3(new_n671), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n721), .A2(new_n579), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n731), .A2(new_n699), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(G29gat), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n728), .A2(new_n729), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT110), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n728), .A2(new_n729), .A3(new_n738), .A4(new_n735), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(G1328gat));
  AND2_X1   g539(.A1(new_n731), .A2(new_n732), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n741), .A2(new_n702), .A3(new_n733), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G36gat), .ZN(new_n743));
  INV_X1    g542(.A(G36gat), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n595), .A2(new_n744), .A3(new_n702), .A4(new_n724), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n745), .A2(new_n746), .A3(KEYINPUT46), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n746), .B1(new_n745), .B2(KEYINPUT46), .ZN(new_n748));
  OAI221_X1 g547(.A(new_n743), .B1(KEYINPUT46), .B2(new_n745), .C1(new_n747), .C2(new_n748), .ZN(G1329gat));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n731), .A2(new_n332), .A3(new_n732), .A4(new_n733), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G43gat), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n713), .A2(G43gat), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n595), .A2(new_n724), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n750), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT47), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n755), .B(new_n756), .ZN(G1330gat));
  NAND3_X1  g556(.A1(new_n595), .A2(new_n497), .A3(new_n724), .ZN(new_n758));
  INV_X1    g557(.A(G50gat), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n741), .A2(G50gat), .A3(new_n497), .A4(new_n733), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(KEYINPUT48), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT48), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n760), .A2(new_n761), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(G1331gat));
  NOR2_X1   g565(.A1(new_n634), .A2(new_n671), .ZN(new_n767));
  AND4_X1   g566(.A1(new_n579), .A2(new_n589), .A3(new_n767), .A4(new_n693), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n699), .ZN(new_n769));
  XNOR2_X1  g568(.A(KEYINPUT113), .B(G57gat), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n769), .B(new_n770), .ZN(G1332gat));
  XNOR2_X1  g570(.A(new_n702), .B(KEYINPUT114), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT49), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n774), .B2(new_n600), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT115), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n768), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n774), .A2(new_n600), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n777), .B(new_n778), .ZN(G1333gat));
  AOI21_X1  g578(.A(G71gat), .B1(new_n768), .B2(new_n714), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n332), .A2(G71gat), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n780), .B1(new_n768), .B2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n782), .B(new_n783), .ZN(G1334gat));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n497), .ZN(new_n785));
  XNOR2_X1  g584(.A(KEYINPUT116), .B(G78gat), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(G1335gat));
  NAND2_X1  g586(.A1(new_n632), .A2(new_n633), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n788), .A2(new_n593), .A3(new_n692), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n741), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(G85gat), .B1(new_n790), .B2(new_n698), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n723), .B1(new_n585), .B2(new_n588), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n788), .A2(new_n593), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n792), .A2(KEYINPUT51), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT51), .B1(new_n792), .B2(new_n793), .ZN(new_n795));
  OR2_X1    g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n796), .A2(new_n636), .A3(new_n693), .A4(new_n699), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n791), .A2(new_n797), .ZN(G1336gat));
  OAI21_X1  g597(.A(G92gat), .B1(new_n790), .B2(new_n772), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n772), .A2(G92gat), .A3(new_n692), .ZN(new_n800));
  AOI21_X1  g599(.A(KEYINPUT52), .B1(new_n796), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n741), .A2(new_n702), .A3(new_n789), .ZN(new_n803));
  AOI22_X1  g602(.A1(new_n803), .A2(G92gat), .B1(new_n796), .B2(new_n800), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(G1337gat));
  OAI21_X1  g605(.A(G99gat), .B1(new_n790), .B2(new_n587), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n713), .A2(G99gat), .A3(new_n692), .ZN(new_n808));
  XOR2_X1   g607(.A(new_n808), .B(KEYINPUT117), .Z(new_n809));
  NAND2_X1  g608(.A1(new_n796), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n807), .A2(new_n810), .ZN(G1338gat));
  INV_X1    g610(.A(KEYINPUT119), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n731), .A2(new_n497), .A3(new_n732), .A4(new_n789), .ZN(new_n813));
  XOR2_X1   g612(.A(KEYINPUT118), .B(G106gat), .Z(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n392), .A2(G106gat), .A3(new_n692), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n817), .B1(new_n794), .B2(new_n795), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n812), .B1(new_n819), .B2(KEYINPUT53), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n821));
  AOI211_X1 g620(.A(KEYINPUT119), .B(new_n821), .C1(new_n816), .C2(new_n818), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n813), .A2(KEYINPUT120), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n813), .A2(KEYINPUT120), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n814), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n818), .A2(new_n821), .ZN(new_n826));
  OAI22_X1  g625(.A1(new_n820), .A2(new_n822), .B1(new_n825), .B2(new_n826), .ZN(G1339gat));
  NAND2_X1  g626(.A1(new_n562), .A2(new_n564), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT121), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n573), .A2(new_n545), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n557), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n693), .A2(new_n566), .A3(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n680), .A2(new_n681), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n685), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n836), .A2(KEYINPUT54), .A3(new_n683), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n674), .B1(new_n683), .B2(KEYINPUT54), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n834), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n839), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n841), .A2(KEYINPUT55), .A3(new_n837), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n840), .A2(new_n691), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n833), .B1(new_n579), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n723), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n832), .A2(new_n566), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n722), .A2(new_n847), .A3(new_n668), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n634), .ZN(new_n850));
  AND4_X1   g649(.A1(new_n579), .A2(new_n788), .A3(new_n723), .A4(new_n692), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n773), .A2(new_n698), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n853), .A2(new_n582), .A3(new_n854), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n855), .A2(new_n263), .A3(new_n579), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n853), .A2(new_n854), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n392), .A2(new_n327), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n593), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n856), .B1(new_n860), .B2(new_n263), .ZN(G1340gat));
  NOR3_X1   g660(.A1(new_n855), .A2(new_n268), .A3(new_n692), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n859), .A2(new_n693), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n863), .B2(new_n268), .ZN(G1341gat));
  NAND4_X1  g663(.A1(new_n859), .A2(new_n282), .A3(new_n284), .A4(new_n788), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n282), .A2(new_n284), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n866), .B1(new_n855), .B2(new_n634), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(G1342gat));
  OAI21_X1  g667(.A(G134gat), .B1(new_n855), .B2(new_n723), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n788), .B1(new_n845), .B2(new_n848), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n870), .A2(new_n851), .ZN(new_n871));
  NOR4_X1   g670(.A1(new_n871), .A2(new_n702), .A3(new_n723), .A4(new_n698), .ZN(new_n872));
  INV_X1    g671(.A(new_n858), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n872), .A2(new_n257), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(KEYINPUT122), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT122), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n872), .A2(new_n876), .A3(new_n257), .A4(new_n873), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n875), .A2(KEYINPUT56), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT56), .B1(new_n875), .B2(new_n877), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n869), .B1(new_n878), .B2(new_n879), .ZN(G1343gat));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n854), .A2(new_n587), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(G141gat), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n579), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT57), .B1(new_n853), .B2(new_n497), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT57), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n871), .A2(new_n887), .A3(new_n392), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n883), .B(new_n885), .C1(new_n886), .C2(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n332), .A2(new_n392), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n853), .A2(new_n854), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n884), .B1(new_n891), .B2(new_n579), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n889), .A2(KEYINPUT58), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(KEYINPUT58), .B1(new_n889), .B2(new_n892), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n881), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n889), .A2(new_n892), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT58), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n889), .A2(KEYINPUT58), .A3(new_n892), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n898), .A2(KEYINPUT123), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n895), .A2(new_n900), .ZN(G1344gat));
  INV_X1    g700(.A(new_n891), .ZN(new_n902));
  INV_X1    g701(.A(G148gat), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(new_n903), .A3(new_n693), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n853), .A2(KEYINPUT57), .A3(new_n497), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n887), .B1(new_n871), .B2(new_n392), .ZN(new_n907));
  AOI211_X1 g706(.A(new_n692), .B(new_n882), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n903), .A2(KEYINPUT59), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n905), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n883), .B1(new_n886), .B2(new_n888), .ZN(new_n912));
  OAI211_X1 g711(.A(KEYINPUT124), .B(new_n909), .C1(new_n912), .C2(new_n692), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT59), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n846), .A2(new_n692), .ZN(new_n916));
  INV_X1    g715(.A(new_n843), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n593), .B2(new_n917), .ZN(new_n918));
  OAI211_X1 g717(.A(KEYINPUT125), .B(new_n848), .C1(new_n918), .C2(new_n671), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(KEYINPUT125), .B1(new_n845), .B2(new_n848), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n634), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(new_n852), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT57), .B1(new_n923), .B2(new_n497), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n693), .B(new_n883), .C1(new_n924), .C2(new_n888), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n915), .B1(new_n925), .B2(G148gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n904), .B1(new_n914), .B2(new_n926), .ZN(G1345gat));
  OAI21_X1  g726(.A(G155gat), .B1(new_n912), .B2(new_n634), .ZN(new_n928));
  OR3_X1    g727(.A1(new_n891), .A2(G155gat), .A3(new_n634), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(G1346gat));
  OAI21_X1  g729(.A(G162gat), .B1(new_n912), .B2(new_n723), .ZN(new_n931));
  INV_X1    g730(.A(G162gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n872), .A2(new_n932), .A3(new_n890), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1347gat));
  NOR3_X1   g733(.A1(new_n871), .A2(new_n699), .A3(new_n772), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n935), .A2(new_n873), .ZN(new_n936));
  INV_X1    g735(.A(new_n228), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n936), .A2(new_n593), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n698), .A2(new_n702), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n939), .A2(new_n507), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n853), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(KEYINPUT126), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n853), .A2(new_n940), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n945), .A2(new_n579), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n938), .B1(new_n946), .B2(new_n206), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT127), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI211_X1 g748(.A(KEYINPUT127), .B(new_n938), .C1(new_n946), .C2(new_n206), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1348gat));
  OAI21_X1  g750(.A(G176gat), .B1(new_n945), .B2(new_n692), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n936), .A2(new_n207), .A3(new_n693), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1349gat));
  NAND3_X1  g753(.A1(new_n936), .A2(new_n244), .A3(new_n788), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n945), .A2(new_n634), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n955), .B1(new_n956), .B2(new_n234), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(KEYINPUT60), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT60), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n959), .B(new_n955), .C1(new_n956), .C2(new_n234), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(G1350gat));
  NAND3_X1  g760(.A1(new_n936), .A2(new_n238), .A3(new_n671), .ZN(new_n962));
  OAI21_X1  g761(.A(G190gat), .B1(new_n945), .B2(new_n723), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n963), .A2(KEYINPUT61), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n963), .A2(KEYINPUT61), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(G1351gat));
  AND2_X1   g765(.A1(new_n935), .A2(new_n890), .ZN(new_n967));
  AOI21_X1  g766(.A(G197gat), .B1(new_n967), .B2(new_n593), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n924), .A2(new_n888), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n939), .A2(new_n332), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n593), .A2(G197gat), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n968), .B1(new_n972), .B2(new_n973), .ZN(G1352gat));
  INV_X1    g773(.A(G204gat), .ZN(new_n975));
  AND4_X1   g774(.A1(new_n975), .A2(new_n935), .A3(new_n693), .A4(new_n890), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n976), .B(KEYINPUT62), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n969), .A2(new_n692), .A3(new_n971), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n977), .B1(new_n975), .B2(new_n978), .ZN(G1353gat));
  INV_X1    g778(.A(G211gat), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n967), .A2(new_n980), .A3(new_n788), .ZN(new_n981));
  OAI211_X1 g780(.A(new_n788), .B(new_n970), .C1(new_n924), .C2(new_n888), .ZN(new_n982));
  AND3_X1   g781(.A1(new_n982), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n983));
  AOI21_X1  g782(.A(KEYINPUT63), .B1(new_n982), .B2(G211gat), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n981), .B1(new_n983), .B2(new_n984), .ZN(G1354gat));
  INV_X1    g784(.A(G218gat), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n967), .A2(new_n986), .A3(new_n671), .ZN(new_n987));
  NOR3_X1   g786(.A1(new_n969), .A2(new_n723), .A3(new_n971), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n987), .B1(new_n988), .B2(new_n986), .ZN(G1355gat));
endmodule


