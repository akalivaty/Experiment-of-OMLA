//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 0 1 1 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 1 1 1 0 1 1 0 1 1 0 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n551, new_n552, new_n553, new_n554, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n564, new_n566,
    new_n567, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n618,
    new_n620, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1145, new_n1146, new_n1147;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT65), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT67), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT68), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT70), .Z(G217));
  NOR4_X1   g027(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT71), .Z(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  AND2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT72), .B(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND4_X1  g041(.A1(new_n464), .A2(new_n466), .A3(KEYINPUT73), .A4(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(KEYINPUT73), .B1(new_n470), .B2(G125), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n462), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT75), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(KEYINPUT3), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n465), .A2(KEYINPUT75), .ZN(new_n476));
  OAI21_X1  g051(.A(G2104), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  XOR2_X1   g052(.A(KEYINPUT72), .B(G2105), .Z(new_n478));
  NAND2_X1  g053(.A1(new_n463), .A2(KEYINPUT74), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT74), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2104), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n479), .A2(new_n481), .A3(KEYINPUT3), .ZN(new_n482));
  NAND4_X1  g057(.A1(new_n477), .A2(G137), .A3(new_n478), .A4(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(G2105), .B1(new_n479), .B2(new_n481), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G101), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n473), .A2(new_n486), .ZN(G160));
  AND2_X1   g062(.A1(new_n477), .A2(new_n482), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(new_n462), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  OAI221_X1 g066(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n478), .C2(G112), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n488), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n493), .B1(G136), .B2(new_n496), .ZN(G162));
  AND2_X1   g072(.A1(G126), .A2(G2105), .ZN(new_n498));
  XNOR2_X1  g073(.A(KEYINPUT75), .B(KEYINPUT3), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n482), .B(new_n498), .C1(new_n463), .C2(new_n499), .ZN(new_n500));
  MUX2_X1   g075(.A(G102), .B(G114), .S(G2105), .Z(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G2104), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n477), .A2(G138), .A3(new_n478), .A4(new_n482), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n464), .A2(new_n466), .A3(G138), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT76), .B(KEYINPUT4), .ZN(new_n507));
  NOR3_X1   g082(.A1(new_n506), .A2(new_n462), .A3(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n503), .B1(new_n505), .B2(new_n509), .ZN(G164));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT77), .B1(new_n511), .B2(G651), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT77), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n513), .A2(new_n514), .A3(KEYINPUT6), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g091(.A(KEYINPUT78), .B1(new_n514), .B2(KEYINPUT6), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT78), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(new_n511), .A3(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AND3_X1   g095(.A1(new_n516), .A2(new_n520), .A3(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G50), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT79), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT79), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n521), .A2(new_n524), .A3(G50), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n516), .A2(new_n520), .ZN(new_n527));
  OR2_X1    g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(KEYINPUT5), .A2(G543), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(G75), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(new_n530), .ZN(new_n533));
  INV_X1    g108(.A(G62), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n531), .A2(G88), .B1(G651), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n526), .A2(new_n536), .ZN(G303));
  INV_X1    g112(.A(G303), .ZN(G166));
  NAND2_X1  g113(.A1(new_n521), .A2(G51), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(KEYINPUT7), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(KEYINPUT7), .ZN(new_n542));
  AND2_X1   g117(.A1(G63), .A2(G651), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n541), .A2(new_n542), .B1(new_n530), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n527), .A2(new_n530), .ZN(new_n545));
  INV_X1    g120(.A(G89), .ZN(new_n546));
  OAI211_X1 g121(.A(new_n539), .B(new_n544), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(KEYINPUT80), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(KEYINPUT80), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(G168));
  NAND2_X1  g125(.A1(new_n531), .A2(G90), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n521), .A2(G52), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n530), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(new_n514), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(G301));
  INV_X1    g130(.A(G301), .ZN(G171));
  NAND2_X1  g131(.A1(new_n521), .A2(G43), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n530), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G81), .ZN(new_n559));
  OAI221_X1 g134(.A(new_n557), .B1(new_n514), .B2(new_n558), .C1(new_n545), .C2(new_n559), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT81), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(new_n562));
  XOR2_X1   g137(.A(new_n562), .B(KEYINPUT82), .Z(G153));
  AND3_X1   g138(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G36), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n564), .A2(new_n567), .ZN(G188));
  NAND2_X1  g143(.A1(new_n521), .A2(G53), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT9), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n530), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT83), .B1(new_n571), .B2(new_n514), .ZN(new_n572));
  INV_X1    g147(.A(G91), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n545), .B2(new_n573), .ZN(new_n574));
  NOR3_X1   g149(.A1(new_n571), .A2(KEYINPUT83), .A3(new_n514), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n570), .A2(new_n576), .ZN(G299));
  INV_X1    g152(.A(G168), .ZN(G286));
  INV_X1    g153(.A(G74), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n528), .A2(new_n579), .A3(new_n529), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G651), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT84), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n580), .A2(KEYINPUT84), .A3(G651), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n516), .A2(new_n520), .A3(G87), .A4(new_n530), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n516), .A2(new_n520), .A3(G49), .A4(G543), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(G288));
  NAND4_X1  g163(.A1(new_n516), .A2(new_n520), .A3(G86), .A4(new_n530), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n516), .A2(new_n520), .A3(G48), .A4(G543), .ZN(new_n590));
  INV_X1    g165(.A(G61), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n591), .B1(new_n528), .B2(new_n529), .ZN(new_n592));
  AND2_X1   g167(.A1(G73), .A2(G543), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n589), .A2(new_n590), .A3(new_n594), .ZN(G305));
  NAND2_X1  g170(.A1(new_n531), .A2(G85), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n521), .A2(G47), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n530), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n598), .A2(new_n514), .ZN(new_n599));
  AND3_X1   g174(.A1(new_n596), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G290));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NOR2_X1   g177(.A1(G301), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n531), .A2(G92), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n604), .B(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n533), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(G54), .A2(new_n521), .B1(new_n609), .B2(G651), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n603), .B1(new_n612), .B2(new_n602), .ZN(G284));
  AOI21_X1  g188(.A(new_n603), .B1(new_n612), .B2(new_n602), .ZN(G321));
  NAND2_X1  g189(.A1(G299), .A2(new_n602), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G168), .B2(new_n602), .ZN(G297));
  OAI21_X1  g191(.A(new_n615), .B1(G168), .B2(new_n602), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n612), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n561), .A2(new_n602), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n612), .A2(new_n618), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n602), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT85), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n484), .A2(new_n470), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT13), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2100), .ZN(new_n629));
  OAI221_X1 g204(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n478), .C2(G111), .ZN(new_n630));
  INV_X1    g205(.A(G135), .ZN(new_n631));
  INV_X1    g206(.A(G123), .ZN(new_n632));
  OAI221_X1 g207(.A(new_n630), .B1(new_n495), .B2(new_n631), .C1(new_n632), .C2(new_n489), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(G2096), .Z(new_n634));
  NAND2_X1  g209(.A1(new_n629), .A2(new_n634), .ZN(G156));
  XOR2_X1   g210(.A(KEYINPUT15), .B(G2435), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2427), .ZN(new_n638));
  INV_X1    g213(.A(G2430), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(KEYINPUT14), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT87), .ZN(new_n643));
  XOR2_X1   g218(.A(G1341), .B(G1348), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2451), .B(G2454), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n645), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(G14), .A3(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(G401));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  NOR3_X1   g233(.A1(new_n655), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT18), .ZN(new_n660));
  INV_X1    g235(.A(new_n656), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(KEYINPUT17), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n657), .B1(new_n663), .B2(new_n654), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n664), .B1(new_n655), .B2(new_n662), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n655), .A2(new_n658), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n661), .B1(new_n666), .B2(KEYINPUT17), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n660), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2096), .ZN(new_n669));
  XOR2_X1   g244(.A(KEYINPUT88), .B(G2100), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G227));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1956), .B(G2474), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1961), .B(G1966), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n674), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n674), .A2(new_n677), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT20), .Z(new_n681));
  AOI211_X1 g256(.A(new_n679), .B(new_n681), .C1(new_n674), .C2(new_n678), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1991), .B(G1996), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n684), .B(new_n687), .ZN(G229));
  NOR2_X1   g263(.A1(G16), .A2(G24), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n600), .B2(G16), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT91), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT90), .B(G1986), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(G25), .A2(G29), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n496), .A2(G131), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n490), .A2(G119), .ZN(new_n696));
  OAI221_X1 g271(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n478), .C2(G107), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n694), .B1(new_n699), .B2(G29), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT35), .B(G1991), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(G16), .A2(G23), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT92), .Z(new_n704));
  NAND2_X1  g279(.A1(G288), .A2(KEYINPUT93), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT93), .ZN(new_n706));
  NAND4_X1  g281(.A1(new_n585), .A2(new_n706), .A3(new_n586), .A4(new_n587), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n704), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT33), .B(G1976), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  MUX2_X1   g287(.A(G6), .B(G305), .S(G16), .Z(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT32), .B(G1981), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(G16), .A2(G22), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G166), .B2(G16), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n715), .B1(new_n717), .B2(G1971), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n712), .B(new_n718), .C1(G1971), .C2(new_n717), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n693), .B(new_n702), .C1(KEYINPUT34), .C2(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT94), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(KEYINPUT34), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT95), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT36), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n723), .B(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n709), .A2(G19), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n561), .B2(new_n709), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(G1341), .Z(new_n730));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n633), .A2(new_n731), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT97), .Z(new_n733));
  INV_X1    g308(.A(G2084), .ZN(new_n734));
  NAND2_X1  g309(.A1(G160), .A2(G29), .ZN(new_n735));
  INV_X1    g310(.A(G34), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n736), .A2(KEYINPUT24), .ZN(new_n737));
  AOI21_X1  g312(.A(G29), .B1(new_n736), .B2(KEYINPUT24), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(KEYINPUT96), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(KEYINPUT96), .B2(new_n738), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n735), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n733), .B1(new_n734), .B2(new_n741), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT31), .B(G11), .Z(new_n743));
  INV_X1    g318(.A(KEYINPUT30), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n731), .B1(new_n744), .B2(G28), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n746), .A2(KEYINPUT98), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n746), .A2(KEYINPUT98), .B1(new_n744), .B2(G28), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n743), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n731), .A2(G32), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT26), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n751), .A2(new_n752), .ZN(new_n754));
  AOI22_X1  g329(.A1(G105), .A2(new_n484), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G141), .ZN(new_n756));
  INV_X1    g331(.A(G129), .ZN(new_n757));
  OAI221_X1 g332(.A(new_n755), .B1(new_n495), .B2(new_n756), .C1(new_n757), .C2(new_n489), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n750), .B1(new_n758), .B2(G29), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT27), .B(G1996), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n742), .B(new_n749), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n496), .A2(G139), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n478), .A2(G103), .A3(G2104), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT25), .Z(new_n764));
  AOI22_X1  g339(.A1(new_n470), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n762), .B(new_n764), .C1(new_n478), .C2(new_n765), .ZN(new_n766));
  MUX2_X1   g341(.A(G33), .B(new_n766), .S(G29), .Z(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(G2072), .Z(new_n768));
  NOR2_X1   g343(.A1(G171), .A2(new_n709), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G5), .B2(new_n709), .ZN(new_n770));
  INV_X1    g345(.A(G1961), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n770), .A2(new_n771), .B1(new_n759), .B2(new_n760), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n768), .B(new_n772), .C1(new_n734), .C2(new_n741), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n731), .A2(G26), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT28), .Z(new_n775));
  OAI221_X1 g350(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n478), .C2(G116), .ZN(new_n776));
  INV_X1    g351(.A(G140), .ZN(new_n777));
  INV_X1    g352(.A(G128), .ZN(new_n778));
  OAI221_X1 g353(.A(new_n776), .B1(new_n495), .B2(new_n777), .C1(new_n778), .C2(new_n489), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n775), .B1(new_n779), .B2(G29), .ZN(new_n780));
  INV_X1    g355(.A(G2067), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n731), .A2(G27), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT100), .Z(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G164), .B2(new_n731), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G2078), .ZN(new_n786));
  NOR4_X1   g361(.A1(new_n761), .A2(new_n773), .A3(new_n782), .A4(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(G4), .A2(G16), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n612), .B2(G16), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1348), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n709), .A2(G20), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT23), .Z(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G299), .B2(G16), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1956), .ZN(new_n794));
  NOR2_X1   g369(.A1(G29), .A2(G35), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G162), .B2(G29), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT29), .Z(new_n797));
  INV_X1    g372(.A(G2090), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n794), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AOI211_X1 g374(.A(new_n790), .B(new_n799), .C1(new_n798), .C2(new_n797), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n770), .A2(new_n771), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT99), .Z(new_n802));
  NOR2_X1   g377(.A1(G16), .A2(G21), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G168), .B2(G16), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n804), .A2(G1966), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n804), .A2(G1966), .ZN(new_n806));
  NOR3_X1   g381(.A1(new_n802), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  AND4_X1   g382(.A1(new_n730), .A2(new_n787), .A3(new_n800), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n727), .A2(new_n808), .ZN(G150));
  INV_X1    g384(.A(G150), .ZN(G311));
  NOR2_X1   g385(.A1(new_n611), .A2(new_n618), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT38), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n531), .A2(G93), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n521), .A2(G55), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n530), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(new_n514), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n813), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n561), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n560), .A2(new_n814), .A3(new_n813), .A4(new_n816), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n812), .B(new_n821), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n822), .A2(KEYINPUT39), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n822), .A2(KEYINPUT39), .ZN(new_n824));
  NOR3_X1   g399(.A1(new_n823), .A2(new_n824), .A3(G860), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n817), .A2(G860), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT101), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT37), .Z(new_n828));
  OR2_X1    g403(.A1(new_n825), .A2(new_n828), .ZN(G145));
  INV_X1    g404(.A(G37), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n698), .B(KEYINPUT102), .Z(new_n831));
  OAI221_X1 g406(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n478), .C2(G118), .ZN(new_n832));
  INV_X1    g407(.A(G130), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n489), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(G142), .B2(new_n496), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(new_n627), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n831), .B(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n766), .B(new_n758), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n779), .B(G164), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n837), .A2(new_n840), .ZN(new_n842));
  AND2_X1   g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(G162), .B(G160), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n633), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n841), .A2(KEYINPUT103), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n847), .A2(new_n842), .A3(new_n846), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n841), .A2(KEYINPUT103), .ZN(new_n849));
  OAI221_X1 g424(.A(new_n830), .B1(new_n843), .B2(new_n846), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g426(.A1(new_n817), .A2(G868), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n708), .B(new_n600), .Z(new_n853));
  XOR2_X1   g428(.A(G303), .B(G305), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(G299), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n611), .A2(new_n857), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n858), .A2(KEYINPUT104), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(KEYINPUT104), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n612), .A2(G299), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT41), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n820), .B(new_n621), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n862), .A2(KEYINPUT41), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(KEYINPUT105), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT105), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n865), .A2(new_n866), .A3(new_n867), .A4(new_n870), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n863), .A2(new_n866), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n869), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT42), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n873), .A2(KEYINPUT42), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n856), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n873), .A2(KEYINPUT42), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n878), .A2(new_n855), .A3(new_n874), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n852), .B1(new_n880), .B2(G868), .ZN(G295));
  AOI21_X1  g456(.A(new_n852), .B1(new_n880), .B2(G868), .ZN(G331));
  NOR2_X1   g457(.A1(G286), .A2(G301), .ZN(new_n883));
  NOR2_X1   g458(.A1(G168), .A2(G171), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n821), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n883), .A2(new_n884), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n820), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n886), .A2(new_n862), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n865), .A2(new_n867), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n885), .A2(KEYINPUT106), .A3(new_n821), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT106), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n892), .B1(new_n887), .B2(new_n820), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n891), .A2(new_n888), .A3(new_n893), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n889), .B(new_n856), .C1(new_n890), .C2(new_n894), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n895), .A2(new_n830), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n886), .A2(new_n888), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n865), .A2(new_n867), .A3(new_n897), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n891), .A2(new_n893), .A3(new_n862), .A4(new_n888), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n855), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT107), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT107), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n900), .A2(new_n903), .A3(new_n855), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n896), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n889), .B1(new_n890), .B2(new_n894), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n855), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n896), .A2(KEYINPUT43), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n907), .A2(new_n908), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n904), .A2(new_n830), .A3(new_n895), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n903), .B1(new_n900), .B2(new_n855), .ZN(new_n914));
  OAI211_X1 g489(.A(KEYINPUT108), .B(KEYINPUT43), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n896), .A2(new_n906), .A3(new_n910), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(KEYINPUT44), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT108), .B1(new_n905), .B2(KEYINPUT43), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n912), .B1(new_n917), .B2(new_n918), .ZN(G397));
  INV_X1    g494(.A(KEYINPUT45), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(G164), .B2(G1384), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n472), .A2(G40), .A3(new_n485), .A4(new_n483), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n779), .B(new_n781), .ZN(new_n924));
  INV_X1    g499(.A(G1996), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n758), .B(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  XOR2_X1   g502(.A(new_n698), .B(new_n701), .Z(new_n928));
  OAI21_X1  g503(.A(new_n923), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AND2_X1   g504(.A1(G290), .A2(G1986), .ZN(new_n930));
  NOR2_X1   g505(.A1(G290), .A2(G1986), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n923), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(KEYINPUT109), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT63), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT55), .ZN(new_n937));
  INV_X1    g512(.A(G8), .ZN(new_n938));
  AOI211_X1 g513(.A(new_n937), .B(new_n938), .C1(new_n526), .C2(new_n536), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT50), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(G164), .B2(G1384), .ZN(new_n942));
  INV_X1    g517(.A(G1384), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n508), .B1(new_n504), .B2(KEYINPUT4), .ZN(new_n944));
  OAI211_X1 g519(.A(KEYINPUT50), .B(new_n943), .C1(new_n944), .C2(new_n503), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n922), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n922), .ZN(new_n947));
  OAI211_X1 g522(.A(KEYINPUT45), .B(new_n943), .C1(new_n944), .C2(new_n503), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n921), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G1971), .ZN(new_n950));
  AOI22_X1  g525(.A1(new_n798), .A2(new_n946), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n940), .B1(new_n951), .B2(new_n938), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT118), .ZN(new_n953));
  XOR2_X1   g528(.A(KEYINPUT110), .B(G8), .Z(new_n954));
  NAND2_X1  g529(.A1(new_n505), .A2(new_n509), .ZN(new_n955));
  INV_X1    g530(.A(new_n503), .ZN(new_n956));
  AOI21_X1  g531(.A(G1384), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n954), .B1(new_n957), .B2(new_n947), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n705), .A2(G1976), .A3(new_n707), .ZN(new_n959));
  XOR2_X1   g534(.A(KEYINPUT111), .B(G1976), .Z(new_n960));
  AOI21_X1  g535(.A(KEYINPUT52), .B1(G288), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT112), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT112), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n958), .A2(new_n964), .A3(new_n959), .A4(new_n961), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g541(.A(KEYINPUT113), .B(G86), .Z(new_n967));
  NAND4_X1  g542(.A1(new_n516), .A2(new_n967), .A3(new_n520), .A4(new_n530), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n968), .A2(new_n590), .A3(new_n594), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(G1981), .ZN(new_n970));
  INV_X1    g545(.A(G1981), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n589), .A2(new_n590), .A3(new_n594), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT49), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n970), .A2(KEYINPUT49), .A3(new_n972), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n954), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n943), .B1(new_n944), .B2(new_n503), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n978), .B1(new_n979), .B2(new_n922), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT114), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n958), .A2(new_n982), .A3(new_n976), .A4(new_n975), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n958), .A2(new_n959), .ZN(new_n984));
  AOI22_X1  g559(.A1(new_n981), .A2(new_n983), .B1(new_n984), .B2(KEYINPUT52), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n952), .A2(new_n953), .A3(new_n966), .A4(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1966), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT117), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n921), .A2(new_n988), .A3(new_n947), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n948), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n922), .B1(new_n979), .B2(new_n920), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n991), .A2(new_n988), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n987), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n946), .A2(new_n734), .ZN(new_n994));
  AOI211_X1 g569(.A(G286), .B(new_n954), .C1(new_n993), .C2(new_n994), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n986), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n985), .A2(new_n966), .ZN(new_n997));
  OR2_X1    g572(.A1(new_n936), .A2(new_n939), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n949), .A2(new_n950), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n942), .A2(new_n945), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n947), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n999), .B1(new_n1001), .B2(G2090), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n998), .B1(new_n1002), .B2(G8), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT118), .B1(new_n997), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n935), .B1(new_n996), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n997), .A2(new_n935), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1002), .A2(new_n998), .A3(G8), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT116), .ZN(new_n1010));
  XOR2_X1   g585(.A(new_n972), .B(KEYINPUT115), .Z(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n981), .A2(new_n983), .ZN(new_n1013));
  NOR2_X1   g588(.A1(G288), .A2(G1976), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1010), .B(new_n1012), .C1(new_n1013), .C2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1015), .B1(new_n981), .B2(new_n983), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT116), .B1(new_n1017), .B2(new_n1011), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1016), .A2(new_n958), .A3(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n940), .B1(new_n951), .B2(new_n954), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1007), .A2(new_n1020), .A3(new_n966), .A4(new_n985), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n993), .A2(new_n994), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1022), .A2(new_n935), .A3(G168), .A4(new_n978), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1009), .B(new_n1019), .C1(new_n1021), .C2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT119), .B1(new_n1005), .B2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1004), .A2(new_n986), .A3(new_n995), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT63), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n1009), .A2(new_n1019), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT119), .ZN(new_n1029));
  OR2_X1    g604(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1025), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT127), .ZN(new_n1033));
  INV_X1    g608(.A(G1956), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1001), .A2(KEYINPUT120), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT120), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1036), .B1(new_n946), .B2(G1956), .ZN(new_n1037));
  XOR2_X1   g612(.A(KEYINPUT56), .B(G2072), .Z(new_n1038));
  OR2_X1    g613(.A1(new_n949), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1035), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  AND2_X1   g615(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1041));
  NOR2_X1   g616(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G1348), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n957), .A2(new_n947), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1001), .A2(new_n1046), .B1(new_n781), .B2(new_n1048), .ZN(new_n1049));
  OR2_X1    g624(.A1(new_n1049), .A2(new_n611), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1045), .A2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1043), .A2(new_n1035), .A3(new_n1037), .A4(new_n1039), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT121), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1051), .A2(KEYINPUT121), .A3(new_n1052), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT123), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1045), .A2(KEYINPUT61), .A3(new_n1052), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT58), .B(G1341), .ZN(new_n1060));
  OAI22_X1  g635(.A1(new_n949), .A2(G1996), .B1(new_n1048), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1061), .A2(KEYINPUT122), .A3(new_n561), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT59), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1061), .A2(KEYINPUT122), .A3(new_n561), .A4(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1059), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT61), .B1(new_n1045), .B2(new_n1052), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1058), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1045), .A2(new_n1052), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT61), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1072), .A2(KEYINPUT123), .A3(new_n1059), .A4(new_n1066), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1069), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1049), .A2(KEYINPUT60), .ZN(new_n1075));
  OR3_X1    g650(.A1(new_n1075), .A2(KEYINPUT124), .A3(new_n612), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT124), .B1(new_n1075), .B2(new_n612), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1075), .A2(new_n612), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n1049), .A2(KEYINPUT60), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1057), .B1(new_n1074), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(new_n949), .B2(G2078), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1001), .A2(new_n771), .ZN(new_n1086));
  OR2_X1    g661(.A1(new_n991), .A2(new_n988), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n991), .A2(new_n988), .B1(KEYINPUT45), .B2(new_n957), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G2078), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT53), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1085), .B(new_n1086), .C1(new_n1089), .C2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(G171), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n991), .A2(KEYINPUT53), .A3(new_n1090), .A4(new_n948), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1086), .A2(new_n1085), .A3(G301), .A4(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT126), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1095), .A2(KEYINPUT126), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1083), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n1092), .A2(G171), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1086), .A2(new_n1085), .A3(new_n1094), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1083), .B1(new_n1101), .B2(G171), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1021), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  AND2_X1   g678(.A1(new_n1099), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1022), .A2(G286), .A3(new_n978), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT51), .ZN(new_n1106));
  AOI21_X1  g681(.A(G1966), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1107));
  INV_X1    g682(.A(new_n994), .ZN(new_n1108));
  OAI21_X1  g683(.A(G8), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(G286), .A2(new_n978), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1106), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT125), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1022), .A2(new_n978), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1114), .A2(new_n1106), .A3(new_n1110), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1105), .B1(new_n1113), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1104), .A2(new_n1117), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1032), .B(new_n1033), .C1(new_n1082), .C2(new_n1118), .ZN(new_n1119));
  OR2_X1    g694(.A1(new_n1117), .A2(KEYINPUT62), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1117), .A2(KEYINPUT62), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1021), .A2(new_n1093), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1119), .A2(new_n1123), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1069), .A2(new_n1073), .B1(new_n1080), .B2(new_n1079), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1104), .B(new_n1117), .C1(new_n1125), .C2(new_n1057), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1033), .B1(new_n1126), .B2(new_n1032), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n934), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n931), .A2(KEYINPUT48), .A3(new_n923), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n929), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT48), .B1(new_n931), .B2(new_n923), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n924), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n923), .B1(new_n1133), .B2(new_n758), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n923), .A2(new_n925), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1135), .A2(KEYINPUT46), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1135), .A2(KEYINPUT46), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1134), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  XOR2_X1   g713(.A(new_n1138), .B(KEYINPUT47), .Z(new_n1139));
  NAND2_X1  g714(.A1(new_n699), .A2(new_n701), .ZN(new_n1140));
  OAI22_X1  g715(.A1(new_n927), .A2(new_n1140), .B1(G2067), .B2(new_n779), .ZN(new_n1141));
  AOI211_X1 g716(.A(new_n1132), .B(new_n1139), .C1(new_n923), .C2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1128), .A2(new_n1142), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g718(.A(G319), .ZN(new_n1145));
  NOR3_X1   g719(.A1(G229), .A2(G227), .A3(new_n1145), .ZN(new_n1146));
  AND3_X1   g720(.A1(new_n850), .A2(new_n652), .A3(new_n1146), .ZN(new_n1147));
  NAND3_X1  g721(.A1(new_n907), .A2(new_n1147), .A3(new_n911), .ZN(G225));
  INV_X1    g722(.A(G225), .ZN(G308));
endmodule


