//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 1 1 1 0 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013;
  XNOR2_X1  g000(.A(G110), .B(G140), .ZN(new_n187));
  INV_X1    g001(.A(G227), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G953), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(G104), .B(G107), .ZN(new_n191));
  INV_X1    g005(.A(G101), .ZN(new_n192));
  OR2_X1    g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G104), .ZN(new_n195));
  AND2_X1   g009(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n196));
  NOR2_X1   g010(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n195), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n198), .B(new_n192), .C1(new_n191), .C2(new_n196), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(G146), .ZN(new_n204));
  NOR3_X1   g018(.A1(new_n200), .A2(KEYINPUT65), .A3(G143), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n201), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(KEYINPUT1), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n203), .A2(G146), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT65), .B1(new_n200), .B2(G143), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n202), .A2(new_n203), .A3(G146), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n207), .B1(new_n201), .B2(KEYINPUT1), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n193), .B(new_n199), .C1(new_n210), .C2(new_n216), .ZN(new_n217));
  AND3_X1   g031(.A1(new_n200), .A2(KEYINPUT64), .A3(G143), .ZN(new_n218));
  AOI21_X1  g032(.A(KEYINPUT64), .B1(new_n200), .B2(G143), .ZN(new_n219));
  OAI22_X1  g033(.A1(new_n218), .A2(new_n219), .B1(G143), .B2(new_n200), .ZN(new_n220));
  INV_X1    g034(.A(new_n215), .ZN(new_n221));
  AOI22_X1  g035(.A1(new_n220), .A2(new_n221), .B1(new_n214), .B2(new_n208), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n199), .A2(new_n193), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n217), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT11), .ZN(new_n226));
  INV_X1    g040(.A(G134), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n226), .B1(new_n227), .B2(G137), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(G137), .ZN(new_n229));
  INV_X1    g043(.A(G137), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n230), .A2(KEYINPUT11), .A3(G134), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n228), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G131), .ZN(new_n233));
  INV_X1    g047(.A(G131), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n228), .A2(new_n231), .A3(new_n234), .A4(new_n229), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n225), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT12), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n225), .A2(KEYINPUT12), .A3(new_n236), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OR2_X1    g055(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n242));
  NAND2_X1  g056(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n242), .A2(new_n243), .B1(G104), .B2(new_n194), .ZN(new_n244));
  INV_X1    g058(.A(G104), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G107), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n196), .B1(new_n246), .B2(new_n195), .ZN(new_n247));
  OAI21_X1  g061(.A(G101), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(new_n199), .A3(KEYINPUT4), .ZN(new_n249));
  NAND2_X1  g063(.A1(KEYINPUT0), .A2(G128), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n220), .A2(new_n253), .B1(new_n214), .B2(new_n251), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n255), .B(G101), .C1(new_n244), .C2(new_n247), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n249), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT79), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT79), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n249), .A2(new_n259), .A3(new_n254), .A4(new_n256), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n233), .A2(new_n235), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT10), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n222), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n223), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n263), .A2(new_n217), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n261), .A2(new_n262), .A3(new_n266), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n241), .A2(KEYINPUT80), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT80), .B1(new_n241), .B2(new_n267), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n190), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n261), .A2(new_n262), .A3(new_n266), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n262), .B1(new_n261), .B2(new_n266), .ZN(new_n272));
  NOR3_X1   g086(.A1(new_n271), .A2(new_n272), .A3(new_n190), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n270), .A2(G469), .A3(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n190), .B1(new_n271), .B2(new_n272), .ZN(new_n276));
  INV_X1    g090(.A(new_n190), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n241), .A2(new_n277), .A3(new_n267), .ZN(new_n278));
  AOI21_X1  g092(.A(G902), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G469), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G902), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n275), .A2(new_n281), .A3(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(KEYINPUT9), .B(G234), .ZN(new_n286));
  OAI21_X1  g100(.A(G221), .B1(new_n286), .B2(G902), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(G214), .B1(G237), .B2(G902), .ZN(new_n289));
  NOR3_X1   g103(.A1(KEYINPUT67), .A2(KEYINPUT2), .A3(G113), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT67), .B1(KEYINPUT2), .B2(G113), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n291), .A2(new_n292), .B1(KEYINPUT2), .B2(G113), .ZN(new_n293));
  INV_X1    g107(.A(G119), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n294), .A2(G116), .ZN(new_n295));
  XNOR2_X1  g109(.A(KEYINPUT69), .B(G119), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n295), .B1(new_n296), .B2(G116), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT68), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n293), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n295), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n294), .A2(KEYINPUT69), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT69), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G119), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G116), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n300), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(KEYINPUT2), .A2(G113), .ZN(new_n307));
  INV_X1    g121(.A(new_n292), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n307), .B1(new_n308), .B2(new_n290), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n306), .A2(new_n309), .A3(KEYINPUT68), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n299), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(new_n249), .A3(new_n256), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n293), .A2(new_n297), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT5), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n296), .A2(new_n314), .A3(G116), .ZN(new_n315));
  OAI211_X1 g129(.A(G113), .B(new_n315), .C1(new_n306), .C2(new_n314), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n265), .A2(new_n313), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(G110), .B(G122), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n312), .A2(new_n319), .A3(new_n317), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(KEYINPUT6), .A3(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G125), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n222), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT64), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n326), .B1(new_n203), .B2(G146), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n200), .A2(KEYINPUT64), .A3(G143), .ZN(new_n328));
  AOI22_X1  g142(.A1(new_n327), .A2(new_n328), .B1(new_n203), .B2(G146), .ZN(new_n329));
  OR2_X1    g143(.A1(new_n251), .A2(new_n252), .ZN(new_n330));
  OAI22_X1  g144(.A1(new_n206), .A2(new_n250), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G125), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n325), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G953), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G224), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n333), .B(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT6), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n318), .A2(new_n338), .A3(new_n320), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n323), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(G210), .B1(G237), .B2(G902), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT83), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT7), .B1(new_n335), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n345), .B1(new_n344), .B2(new_n335), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n325), .A2(new_n332), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT84), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT84), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n325), .A2(new_n332), .A3(new_n349), .A4(new_n346), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n319), .B(KEYINPUT81), .ZN(new_n352));
  XOR2_X1   g166(.A(new_n352), .B(KEYINPUT8), .Z(new_n353));
  INV_X1    g167(.A(new_n317), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n265), .B1(new_n313), .B2(new_n316), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT7), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n336), .B1(KEYINPUT82), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n358), .B1(KEYINPUT82), .B2(new_n357), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n333), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n351), .A2(new_n356), .A3(new_n322), .A4(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n282), .ZN(new_n362));
  NOR3_X1   g176(.A1(new_n341), .A2(new_n343), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n362), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n342), .B1(new_n364), .B2(new_n340), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n289), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n305), .A2(G122), .ZN(new_n367));
  XNOR2_X1  g181(.A(KEYINPUT91), .B(G122), .ZN(new_n368));
  OAI221_X1 g182(.A(new_n367), .B1(KEYINPUT14), .B2(new_n194), .C1(new_n368), .C2(new_n305), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n367), .B1(new_n368), .B2(new_n305), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT14), .B1(new_n368), .B2(new_n305), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n371), .A3(G107), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n203), .A2(G128), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n207), .A2(G143), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n375), .A2(KEYINPUT92), .ZN(new_n376));
  XNOR2_X1  g190(.A(G128), .B(G143), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT92), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NOR3_X1   g193(.A1(new_n376), .A2(new_n379), .A3(new_n227), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n375), .A2(KEYINPUT92), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n377), .A2(new_n378), .ZN(new_n382));
  AOI21_X1  g196(.A(G134), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n369), .B(new_n372), .C1(new_n380), .C2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n377), .A2(KEYINPUT13), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n385), .B(G134), .C1(KEYINPUT13), .C2(new_n373), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n227), .B1(new_n376), .B2(new_n379), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n370), .A2(G107), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n370), .A2(G107), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n386), .B(new_n387), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G217), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n286), .A2(new_n391), .A3(G953), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n384), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n392), .B1(new_n384), .B2(new_n390), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G478), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n396), .B(new_n282), .C1(KEYINPUT15), .C2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT93), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n400), .B1(new_n395), .B2(G902), .ZN(new_n401));
  OAI211_X1 g215(.A(KEYINPUT93), .B(new_n282), .C1(new_n393), .C2(new_n394), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n397), .A2(KEYINPUT15), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n399), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(G475), .A2(G902), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT16), .ZN(new_n407));
  INV_X1    g221(.A(G140), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(new_n408), .A3(G125), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(G125), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n324), .A2(G140), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n409), .B1(new_n412), .B2(new_n407), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n200), .ZN(new_n414));
  OAI211_X1 g228(.A(G146), .B(new_n409), .C1(new_n412), .C2(new_n407), .ZN(new_n415));
  NOR2_X1   g229(.A1(G237), .A2(G953), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(G143), .A3(G214), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(G143), .B1(new_n416), .B2(G214), .ZN(new_n419));
  OAI211_X1 g233(.A(KEYINPUT17), .B(G131), .C1(new_n418), .C2(new_n419), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n414), .A2(new_n415), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT87), .ZN(new_n422));
  INV_X1    g236(.A(G237), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n423), .A2(new_n334), .A3(G214), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n203), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n417), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n422), .B1(new_n426), .B2(G131), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT17), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n425), .A2(KEYINPUT87), .A3(new_n234), .A4(new_n417), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n426), .A2(G131), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n427), .A2(new_n428), .A3(new_n429), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n421), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(G113), .B(G122), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n433), .B(new_n245), .ZN(new_n434));
  NAND2_X1  g248(.A1(KEYINPUT18), .A2(G131), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n425), .A2(new_n435), .A3(new_n417), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT86), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT86), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n425), .A2(new_n438), .A3(new_n435), .A4(new_n417), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n412), .A2(G146), .ZN(new_n441));
  XNOR2_X1  g255(.A(G125), .B(G140), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n200), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NOR3_X1   g258(.A1(new_n418), .A2(new_n419), .A3(KEYINPUT85), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT85), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n446), .B1(new_n425), .B2(new_n417), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n440), .B(new_n444), .C1(new_n448), .C2(new_n435), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n432), .A2(new_n434), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n427), .A2(new_n429), .A3(new_n430), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT19), .ZN(new_n452));
  AOI21_X1  g266(.A(KEYINPUT19), .B1(new_n410), .B2(new_n411), .ZN(new_n453));
  OR2_X1    g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT88), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(new_n455), .A3(new_n200), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n200), .B1(new_n452), .B2(new_n453), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT88), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n451), .A2(new_n456), .A3(new_n458), .A4(new_n415), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n434), .B1(new_n459), .B2(new_n449), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n406), .B1(new_n450), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT20), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT20), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n463), .B(new_n406), .C1(new_n450), .C2(new_n460), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n434), .B1(new_n432), .B2(new_n449), .ZN(new_n466));
  NOR3_X1   g280(.A1(new_n450), .A2(new_n466), .A3(KEYINPUT89), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(KEYINPUT89), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n282), .ZN(new_n469));
  OAI21_X1  g283(.A(G475), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT90), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT90), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n465), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(G234), .A2(G237), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n475), .A2(G952), .A3(new_n334), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n475), .A2(G902), .A3(G953), .ZN(new_n477));
  XNOR2_X1  g291(.A(KEYINPUT21), .B(G898), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n405), .A2(new_n472), .A3(new_n474), .A4(new_n480), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n288), .A2(new_n366), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n334), .A2(G221), .A3(G234), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n483), .B(KEYINPUT74), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT22), .B(G137), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n484), .B(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n414), .A2(new_n415), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n296), .A2(G128), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n294), .A2(G128), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT23), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT73), .ZN(new_n493));
  OR2_X1    g307(.A1(new_n493), .A2(KEYINPUT23), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(KEYINPUT23), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n304), .A2(new_n207), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(G110), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n490), .B1(new_n296), .B2(G128), .ZN(new_n498));
  XOR2_X1   g312(.A(KEYINPUT24), .B(G110), .Z(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n488), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n415), .A2(new_n443), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n494), .A2(new_n495), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n504), .B1(G128), .B2(new_n296), .ZN(new_n505));
  INV_X1    g319(.A(G110), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n505), .A2(new_n506), .A3(new_n489), .A4(new_n491), .ZN(new_n507));
  OR2_X1    g321(.A1(new_n498), .A2(new_n499), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n503), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n487), .B1(new_n502), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n509), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(new_n501), .A3(new_n486), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n391), .B1(G234), .B2(new_n282), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n514), .A2(G902), .ZN(new_n515));
  XOR2_X1   g329(.A(new_n515), .B(KEYINPUT77), .Z(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n510), .A2(new_n512), .A3(new_n282), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT76), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT25), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT75), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT25), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n522), .B1(new_n523), .B2(KEYINPUT76), .ZN(new_n524));
  AOI21_X1  g338(.A(KEYINPUT25), .B1(new_n520), .B2(KEYINPUT75), .ZN(new_n525));
  OAI22_X1  g339(.A1(new_n521), .A2(new_n524), .B1(new_n519), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n518), .B1(new_n526), .B2(new_n514), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT66), .B1(new_n230), .B2(G134), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT66), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n529), .A2(new_n227), .A3(G137), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n230), .A2(G134), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n528), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(G131), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n533), .A2(new_n235), .ZN(new_n534));
  OAI22_X1  g348(.A1(new_n206), .A2(new_n209), .B1(new_n329), .B2(new_n215), .ZN(new_n535));
  AOI22_X1  g349(.A1(new_n534), .A2(new_n535), .B1(new_n254), .B2(new_n236), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n299), .A2(KEYINPUT70), .A3(new_n310), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT70), .B1(new_n299), .B2(new_n310), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT28), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n533), .A2(new_n235), .ZN(new_n542));
  OAI22_X1  g356(.A1(new_n262), .A2(new_n331), .B1(new_n222), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n311), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n536), .B(KEYINPUT28), .C1(new_n537), .C2(new_n538), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n541), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n423), .A2(new_n334), .A3(G210), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT27), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(KEYINPUT26), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(new_n192), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n546), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT30), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n543), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n254), .A2(new_n236), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n556), .B(KEYINPUT30), .C1(new_n222), .C2(new_n542), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n555), .A2(new_n311), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n558), .A2(new_n551), .A3(new_n539), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(KEYINPUT31), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT31), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n558), .A2(new_n551), .A3(new_n561), .A4(new_n539), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n553), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT71), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT71), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n553), .A2(new_n560), .A3(new_n565), .A4(new_n562), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(G472), .A2(G902), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT32), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n541), .A2(new_n545), .ZN(new_n572));
  OR3_X1    g386(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n572), .A2(KEYINPUT29), .A3(new_n551), .A4(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n572), .A2(new_n551), .A3(new_n544), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT72), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n558), .A2(new_n539), .ZN(new_n578));
  AOI21_X1  g392(.A(KEYINPUT29), .B1(new_n578), .B2(new_n552), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n579), .B1(new_n575), .B2(new_n576), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n282), .B(new_n574), .C1(new_n577), .C2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(G472), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n567), .A2(KEYINPUT32), .A3(new_n568), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n571), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n482), .A2(new_n527), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(G101), .ZN(G3));
  AOI21_X1  g400(.A(G902), .B1(new_n564), .B2(new_n566), .ZN(new_n587));
  INV_X1    g401(.A(G472), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(KEYINPUT94), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n587), .B(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n288), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n590), .A2(new_n591), .A3(new_n527), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n472), .A2(new_n474), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT33), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n594), .B1(new_n393), .B2(new_n394), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n384), .A2(new_n390), .ZN(new_n596));
  INV_X1    g410(.A(new_n392), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n384), .A2(new_n390), .A3(new_n392), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(KEYINPUT33), .A3(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n397), .A2(G902), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n595), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT95), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT95), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n595), .A2(new_n600), .A3(new_n604), .A4(new_n601), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT96), .B(G478), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n403), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n593), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n343), .B1(new_n341), .B2(new_n362), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n364), .A2(new_n342), .A3(new_n340), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n613), .A2(new_n289), .A3(new_n480), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n592), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT34), .B(G104), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(KEYINPUT97), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n616), .B(new_n618), .ZN(G6));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n464), .A2(KEYINPUT98), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n620), .B1(new_n464), .B2(KEYINPUT98), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n462), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n464), .A2(KEYINPUT98), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(KEYINPUT99), .ZN(new_n625));
  INV_X1    g439(.A(new_n462), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n464), .A2(KEYINPUT98), .A3(new_n620), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT15), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n403), .A2(new_n630), .A3(G478), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n398), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n629), .A2(new_n470), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(KEYINPUT100), .B1(new_n633), .B2(new_n614), .ZN(new_n634));
  INV_X1    g448(.A(new_n289), .ZN(new_n635));
  AOI211_X1 g449(.A(new_n635), .B(new_n479), .C1(new_n611), .C2(new_n612), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n637));
  INV_X1    g451(.A(new_n470), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n623), .B2(new_n628), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n636), .A2(new_n637), .A3(new_n632), .A4(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n634), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n592), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT35), .B(G107), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  NOR3_X1   g458(.A1(new_n587), .A2(KEYINPUT94), .A3(new_n588), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n502), .A2(new_n509), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n487), .A2(KEYINPUT36), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n648), .A2(new_n649), .A3(new_n517), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n526), .B2(new_n514), .ZN(new_n651));
  AOI211_X1 g465(.A(G902), .B(new_n589), .C1(new_n564), .C2(new_n566), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n645), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT101), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n482), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NOR4_X1   g469(.A1(new_n645), .A2(new_n652), .A3(KEYINPUT101), .A4(new_n651), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT37), .B(G110), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G12));
  AOI21_X1  g473(.A(KEYINPUT32), .B1(new_n567), .B2(new_n568), .ZN(new_n660));
  INV_X1    g474(.A(new_n568), .ZN(new_n661));
  AOI211_X1 g475(.A(new_n570), .B(new_n661), .C1(new_n564), .C2(new_n566), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n651), .B1(new_n663), .B2(new_n582), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT102), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n635), .B1(new_n611), .B2(new_n612), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n285), .A2(new_n666), .A3(new_n287), .ZN(new_n667));
  INV_X1    g481(.A(G900), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n476), .B1(new_n477), .B2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n639), .A2(new_n632), .A3(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n664), .A2(new_n665), .A3(new_n667), .A4(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n651), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n584), .A2(new_n667), .A3(new_n673), .A4(new_n671), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(KEYINPUT102), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT103), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G128), .ZN(G30));
  XOR2_X1   g492(.A(new_n669), .B(KEYINPUT39), .Z(new_n679));
  NAND2_X1  g493(.A1(new_n591), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n680), .B(KEYINPUT40), .Z(new_n681));
  NAND2_X1  g495(.A1(new_n578), .A2(new_n551), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n552), .A2(new_n539), .A3(new_n573), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n682), .A2(new_n683), .A3(new_n282), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(G472), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n571), .A2(new_n583), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT104), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n663), .A2(KEYINPUT104), .A3(new_n685), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n613), .B(KEYINPUT38), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n465), .A2(new_n470), .A3(new_n473), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n473), .B1(new_n465), .B2(new_n470), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n632), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n694), .A2(new_n673), .A3(new_n635), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n681), .A2(new_n690), .A3(new_n691), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G143), .ZN(G45));
  OAI211_X1 g511(.A(new_n609), .B(new_n670), .C1(new_n692), .C2(new_n693), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(KEYINPUT105), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT105), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n593), .A2(new_n700), .A3(new_n609), .A4(new_n670), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n664), .A2(new_n667), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  INV_X1    g518(.A(new_n278), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n254), .A2(new_n256), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n259), .B1(new_n706), .B2(new_n249), .ZN(new_n707));
  INV_X1    g521(.A(new_n260), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n266), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n236), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n277), .B1(new_n710), .B2(new_n267), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n282), .B1(new_n705), .B2(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n280), .A2(KEYINPUT106), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n713), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n279), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n287), .A3(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n584), .A2(new_n615), .A3(new_n527), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT41), .B(G113), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G15));
  AND4_X1   g535(.A1(new_n527), .A2(new_n641), .A3(new_n584), .A4(new_n718), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(new_n305), .ZN(G18));
  NAND4_X1  g537(.A1(new_n666), .A2(new_n287), .A3(new_n716), .A4(new_n714), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(new_n481), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(new_n584), .A3(new_n673), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G119), .ZN(G21));
  NAND2_X1  g541(.A1(new_n560), .A2(new_n562), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n551), .B1(new_n572), .B2(new_n573), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n568), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n527), .B(new_n730), .C1(new_n587), .C2(new_n588), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n731), .A2(new_n479), .A3(new_n717), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n733), .B1(new_n694), .B2(new_n366), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n593), .A2(new_n666), .A3(KEYINPUT107), .A4(new_n632), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  NOR2_X1   g552(.A1(new_n717), .A2(new_n366), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n567), .A2(new_n282), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(G472), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n739), .A2(new_n673), .A3(new_n741), .A4(new_n730), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n699), .A2(new_n701), .ZN(new_n743));
  OAI21_X1  g557(.A(KEYINPUT108), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n673), .B(new_n730), .C1(new_n587), .C2(new_n588), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n724), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n702), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G125), .ZN(G27));
  NAND3_X1  g564(.A1(new_n611), .A2(new_n289), .A3(new_n612), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n288), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n584), .A3(new_n527), .ZN(new_n753));
  AND2_X1   g567(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n754));
  NOR2_X1   g568(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n755));
  OAI22_X1  g569(.A1(new_n753), .A2(new_n743), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n584), .A2(new_n527), .ZN(new_n757));
  INV_X1    g571(.A(new_n755), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n757), .A2(new_n702), .A3(new_n752), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G131), .ZN(G33));
  INV_X1    g575(.A(KEYINPUT110), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n757), .A2(new_n762), .A3(new_n671), .A4(new_n752), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n639), .A2(new_n632), .A3(new_n670), .ZN(new_n764));
  OAI21_X1  g578(.A(KEYINPUT110), .B1(new_n753), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G134), .ZN(G36));
  INV_X1    g581(.A(KEYINPUT45), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n241), .A2(new_n267), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT80), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n241), .A2(KEYINPUT80), .A3(new_n267), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n277), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n768), .B1(new_n773), .B2(new_n273), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n270), .A2(KEYINPUT45), .A3(new_n274), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(G469), .A3(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT111), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n270), .A2(new_n274), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n280), .B1(new_n779), .B2(new_n768), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(KEYINPUT111), .A3(new_n775), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n283), .B1(new_n778), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n281), .B1(new_n782), .B2(KEYINPUT46), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT46), .ZN(new_n784));
  AOI211_X1 g598(.A(new_n784), .B(new_n283), .C1(new_n778), .C2(new_n781), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n287), .B(new_n679), .C1(new_n783), .C2(new_n785), .ZN(new_n786));
  XOR2_X1   g600(.A(new_n786), .B(KEYINPUT112), .Z(new_n787));
  NAND3_X1  g601(.A1(new_n472), .A2(new_n609), .A3(new_n474), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n788), .A2(KEYINPUT43), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(KEYINPUT43), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n673), .B1(new_n645), .B2(new_n652), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT44), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(KEYINPUT44), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(new_n751), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n787), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT113), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(new_n230), .ZN(G39));
  OAI21_X1  g613(.A(new_n287), .B1(new_n783), .B2(new_n785), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(KEYINPUT47), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT47), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n802), .B(new_n287), .C1(new_n783), .C2(new_n785), .ZN(new_n803));
  NOR4_X1   g617(.A1(new_n743), .A2(new_n584), .A3(new_n527), .A4(new_n751), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n801), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G140), .ZN(G42));
  INV_X1    g620(.A(KEYINPUT121), .ZN(new_n807));
  INV_X1    g621(.A(G952), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n334), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT120), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n674), .A2(KEYINPUT102), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n674), .A2(KEYINPUT102), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n749), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n688), .A2(new_n689), .ZN(new_n815));
  AOI211_X1 g629(.A(new_n650), .B(new_n669), .C1(new_n526), .C2(new_n514), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n285), .A2(new_n287), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT116), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n285), .A2(new_n816), .A3(new_n819), .A4(new_n287), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n736), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n703), .B1(new_n815), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n811), .B1(new_n814), .B2(new_n822), .ZN(new_n823));
  OAI211_X1 g637(.A(KEYINPUT52), .B(new_n703), .C1(new_n815), .C2(new_n821), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n823), .B1(new_n814), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n719), .B1(new_n655), .B2(new_n656), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n472), .A2(new_n632), .A3(new_n474), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n614), .B1(new_n610), .B2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n828), .A2(new_n590), .A3(new_n527), .A4(new_n591), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n585), .A2(new_n737), .A3(new_n829), .A4(new_n726), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n826), .A2(new_n830), .A3(new_n722), .ZN(new_n831));
  INV_X1    g645(.A(new_n664), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n639), .A2(new_n405), .A3(new_n670), .ZN(new_n833));
  OAI22_X1  g647(.A1(new_n832), .A2(new_n833), .B1(new_n743), .B2(new_n746), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n752), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n756), .A2(new_n759), .B1(new_n763), .B2(new_n765), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n831), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT53), .B1(new_n825), .B2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n831), .A2(new_n836), .A3(KEYINPUT53), .A4(new_n835), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT117), .B1(new_n814), .B2(new_n824), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n672), .A2(new_n675), .B1(new_n744), .B2(new_n748), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT117), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n736), .A2(new_n818), .A3(new_n820), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n584), .A2(new_n667), .A3(new_n673), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n843), .A2(new_n690), .B1(new_n844), .B2(new_n702), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n841), .A2(new_n842), .A3(new_n845), .A4(KEYINPUT52), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n840), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n839), .B1(new_n847), .B2(new_n823), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n838), .A2(new_n848), .A3(KEYINPUT54), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT52), .B1(new_n841), .B2(new_n845), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n852), .B1(new_n840), .B2(new_n846), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n831), .A2(new_n835), .A3(new_n836), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n851), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n825), .A2(new_n837), .A3(KEYINPUT53), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n850), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n849), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n717), .A2(new_n751), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n859), .A2(new_n527), .A3(new_n476), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n593), .A2(new_n609), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n815), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n789), .A2(new_n859), .A3(new_n476), .A4(new_n790), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n863), .A2(new_n746), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(KEYINPUT118), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n863), .A2(new_n866), .A3(new_n746), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n862), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n789), .A2(new_n476), .A3(new_n790), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n731), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n718), .A2(new_n635), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n871), .A2(new_n691), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n870), .A2(KEYINPUT50), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT50), .B1(new_n870), .B2(new_n872), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n868), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n287), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n714), .A2(new_n716), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  AOI22_X1  g693(.A1(new_n801), .A2(new_n803), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n869), .A2(new_n731), .A3(new_n751), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n876), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT51), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n757), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n886), .A2(new_n863), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT48), .ZN(new_n888));
  AOI211_X1 g702(.A(new_n808), .B(G953), .C1(new_n870), .C2(new_n739), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n815), .A2(new_n860), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n889), .B1(new_n610), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n885), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n876), .B(KEYINPUT51), .C1(new_n880), .C2(new_n882), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT119), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n894), .A2(new_n895), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n893), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n810), .B1(new_n858), .B2(new_n899), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n527), .A2(new_n289), .A3(new_n287), .ZN(new_n901));
  INV_X1    g715(.A(new_n788), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT49), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n901), .B(new_n902), .C1(new_n879), .C2(new_n903), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT114), .Z(new_n905));
  NAND2_X1  g719(.A1(new_n879), .A2(new_n903), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT115), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n907), .A2(new_n691), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n905), .A2(new_n815), .A3(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n807), .B1(new_n900), .B2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n892), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n912), .B1(new_n883), .B2(new_n884), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n894), .A2(new_n895), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n913), .B1(new_n914), .B2(new_n896), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n915), .A2(new_n857), .A3(new_n849), .ZN(new_n916));
  OAI211_X1 g730(.A(KEYINPUT121), .B(new_n909), .C1(new_n916), .C2(new_n810), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n911), .A2(new_n917), .ZN(G75));
  XNOR2_X1  g732(.A(KEYINPUT122), .B(KEYINPUT55), .ZN(new_n919));
  OAI211_X1 g733(.A(G210), .B(G902), .C1(new_n838), .C2(new_n848), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n323), .A2(new_n339), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(new_n337), .ZN(new_n922));
  NOR2_X1   g736(.A1(KEYINPUT123), .A2(KEYINPUT56), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n920), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n922), .B1(new_n920), .B2(new_n923), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n919), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n920), .A2(new_n923), .ZN(new_n927));
  INV_X1    g741(.A(new_n922), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n919), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n920), .A2(new_n922), .A3(new_n923), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n334), .A2(G952), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n926), .A2(new_n932), .A3(new_n934), .ZN(G51));
  XNOR2_X1  g749(.A(new_n283), .B(KEYINPUT57), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n825), .A2(new_n837), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n851), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n853), .A2(new_n839), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n850), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n936), .B1(new_n940), .B2(new_n849), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n941), .B1(new_n711), .B2(new_n705), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n282), .B1(new_n938), .B2(new_n939), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n943), .A2(new_n778), .A3(new_n781), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n933), .B1(new_n942), .B2(new_n944), .ZN(G54));
  NAND3_X1  g759(.A1(new_n943), .A2(KEYINPUT58), .A3(G475), .ZN(new_n946));
  OR2_X1    g760(.A1(new_n450), .A2(new_n460), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n946), .A2(new_n948), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n949), .A2(new_n950), .A3(new_n933), .ZN(G60));
  AND2_X1   g765(.A1(new_n595), .A2(new_n600), .ZN(new_n952));
  INV_X1    g766(.A(new_n858), .ZN(new_n953));
  NAND2_X1  g767(.A1(G478), .A2(G902), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT59), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n952), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n952), .B(new_n955), .C1(new_n940), .C2(new_n849), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n934), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n956), .A2(new_n958), .ZN(G63));
  NAND2_X1  g773(.A1(G217), .A2(G902), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT60), .Z(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(new_n838), .B2(new_n848), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n933), .B1(new_n962), .B2(new_n513), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n938), .A2(new_n939), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n648), .A2(new_n649), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n964), .A2(KEYINPUT124), .A3(new_n965), .A4(new_n961), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n965), .B(new_n961), .C1(new_n838), .C2(new_n848), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT124), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n963), .A2(new_n966), .A3(new_n969), .ZN(new_n970));
  XNOR2_X1  g784(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(G66));
  NOR2_X1   g786(.A1(new_n826), .A2(new_n830), .ZN(new_n973));
  INV_X1    g787(.A(new_n722), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(G224), .A2(G953), .ZN(new_n976));
  OAI22_X1  g790(.A1(new_n975), .A2(G953), .B1(new_n478), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n921), .B1(G898), .B2(new_n334), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n977), .B(new_n978), .Z(G69));
  XOR2_X1   g793(.A(new_n836), .B(KEYINPUT127), .Z(new_n980));
  OR2_X1    g794(.A1(new_n980), .A2(G953), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n841), .A2(new_n703), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n757), .A2(new_n736), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n982), .B1(new_n787), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n984), .A2(new_n797), .A3(new_n805), .ZN(new_n985));
  OAI22_X1  g799(.A1(new_n981), .A2(new_n985), .B1(new_n188), .B2(new_n334), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n555), .A2(new_n557), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n454), .B(KEYINPUT126), .Z(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  OR2_X1    g804(.A1(new_n989), .A2(G227), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n334), .B1(new_n991), .B2(G900), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n696), .A2(new_n703), .A3(new_n841), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT62), .Z(new_n994));
  NOR2_X1   g808(.A1(new_n680), .A2(new_n751), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n610), .A2(new_n827), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n995), .A2(new_n757), .A3(new_n996), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n994), .A2(new_n797), .A3(new_n805), .A4(new_n997), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n989), .A2(G953), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n992), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n990), .A2(new_n1000), .ZN(G72));
  NAND2_X1  g815(.A1(G472), .A2(G902), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(KEYINPUT63), .Z(new_n1003));
  OAI21_X1  g817(.A(new_n1003), .B1(new_n998), .B2(new_n975), .ZN(new_n1004));
  INV_X1    g818(.A(new_n682), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n855), .A2(new_n856), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n578), .A2(new_n551), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n1007), .A2(new_n682), .A3(new_n1003), .A4(new_n1009), .ZN(new_n1010));
  OR2_X1    g824(.A1(new_n980), .A2(new_n975), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1003), .B1(new_n1011), .B2(new_n985), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n933), .B1(new_n1012), .B2(new_n1008), .ZN(new_n1013));
  AND3_X1   g827(.A1(new_n1006), .A2(new_n1010), .A3(new_n1013), .ZN(G57));
endmodule


