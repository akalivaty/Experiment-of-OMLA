//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 1 0 1 0 0 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n865, new_n866, new_n867, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n995,
    new_n996, new_n997;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT11), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G169gat), .ZN(new_n204));
  OR2_X1    g003(.A1(new_n202), .A2(KEYINPUT11), .ZN(new_n205));
  INV_X1    g004(.A(G169gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n202), .A2(KEYINPUT11), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  AOI21_X1  g007(.A(G197gat), .B1(new_n204), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n204), .A2(G197gat), .A3(new_n208), .ZN(new_n211));
  AND3_X1   g010(.A1(new_n210), .A2(KEYINPUT12), .A3(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT12), .B1(new_n210), .B2(new_n211), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT15), .ZN(new_n215));
  INV_X1    g014(.A(G50gat), .ZN(new_n216));
  AND2_X1   g015(.A1(KEYINPUT86), .A2(G43gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(KEYINPUT86), .A2(G43gat), .ZN(new_n218));
  OAI211_X1 g017(.A(KEYINPUT87), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G43gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G50gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT86), .B(G43gat), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT87), .B1(new_n223), .B2(new_n216), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n215), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n215), .B1(new_n220), .B2(G50gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n216), .A2(G43gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT14), .ZN(new_n228));
  AOI21_X1  g027(.A(G36gat), .B1(new_n228), .B2(G29gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n226), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G36gat), .ZN(new_n231));
  INV_X1    g030(.A(G29gat), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n231), .B1(new_n232), .B2(KEYINPUT14), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT15), .B1(new_n216), .B2(G43gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n220), .A2(G50gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n230), .A2(new_n236), .A3(KEYINPUT14), .A4(new_n232), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n232), .A2(KEYINPUT14), .ZN(new_n238));
  NOR3_X1   g037(.A1(new_n234), .A2(new_n233), .A3(new_n235), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n229), .B1(new_n226), .B2(new_n227), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n237), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT17), .ZN(new_n243));
  XNOR2_X1  g042(.A(G15gat), .B(G22gat), .ZN(new_n244));
  INV_X1    g043(.A(G1gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT16), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n247), .B1(G1gat), .B2(new_n244), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(G8gat), .ZN(new_n249));
  INV_X1    g048(.A(G8gat), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n247), .B(new_n250), .C1(G1gat), .C2(new_n244), .ZN(new_n251));
  AND2_X1   g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT17), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n225), .A2(new_n241), .A3(new_n253), .A4(new_n237), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n243), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G229gat), .A2(G233gat), .ZN(new_n256));
  INV_X1    g055(.A(new_n242), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n249), .A2(new_n251), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n255), .A2(new_n256), .A3(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT18), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n255), .A2(KEYINPUT18), .A3(new_n256), .A4(new_n259), .ZN(new_n263));
  XOR2_X1   g062(.A(new_n256), .B(KEYINPUT13), .Z(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n252), .A2(new_n242), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n265), .B1(new_n259), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  AND4_X1   g067(.A1(new_n214), .A2(new_n262), .A3(new_n263), .A4(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n267), .B1(new_n260), .B2(new_n261), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n214), .B1(new_n270), .B2(new_n263), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT36), .ZN(new_n273));
  NAND2_X1  g072(.A1(G227gat), .A2(G233gat), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G113gat), .ZN(new_n276));
  INV_X1    g075(.A(G120gat), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT1), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n278), .B1(new_n276), .B2(new_n277), .ZN(new_n279));
  OR2_X1    g078(.A1(G127gat), .A2(G134gat), .ZN(new_n280));
  INV_X1    g079(.A(G134gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT67), .B(G127gat), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n279), .B(new_n280), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(KEYINPUT68), .ZN(new_n284));
  NAND2_X1  g083(.A1(G127gat), .A2(G134gat), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n279), .B1(new_n280), .B2(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT25), .ZN(new_n288));
  NAND3_X1  g087(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n289), .B1(G183gat), .B2(G190gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT24), .ZN(new_n291));
  NAND2_X1  g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT23), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT23), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n296), .B1(G169gat), .B2(G176gat), .ZN(new_n297));
  INV_X1    g096(.A(G176gat), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n295), .B(new_n297), .C1(new_n206), .C2(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n288), .B1(new_n293), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT64), .ZN(new_n301));
  OR2_X1    g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OR2_X1    g101(.A1(new_n292), .A2(KEYINPUT65), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT24), .B1(new_n292), .B2(KEYINPUT65), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n290), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OR3_X1    g104(.A1(new_n305), .A2(new_n288), .A3(new_n299), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n300), .A2(new_n301), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n302), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n206), .A2(new_n298), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT26), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n309), .B1(new_n310), .B2(new_n294), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n311), .B1(new_n310), .B2(new_n294), .ZN(new_n312));
  XOR2_X1   g111(.A(KEYINPUT27), .B(G183gat), .Z(new_n313));
  INV_X1    g112(.A(KEYINPUT66), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT27), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(G183gat), .ZN(new_n317));
  AOI21_X1  g116(.A(G190gat), .B1(new_n317), .B2(KEYINPUT66), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT28), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT28), .ZN(new_n320));
  NOR3_X1   g119(.A1(new_n313), .A2(new_n320), .A3(G190gat), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n292), .B(new_n312), .C1(new_n319), .C2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n287), .A2(new_n308), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n287), .B1(new_n322), .B2(new_n308), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n323), .B1(new_n324), .B2(KEYINPUT69), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n322), .ZN(new_n326));
  INV_X1    g125(.A(new_n287), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT69), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n275), .B1(new_n325), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT32), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT33), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(G15gat), .B(G43gat), .Z(new_n334));
  XNOR2_X1  g133(.A(G71gat), .B(G99gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n331), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n326), .A2(new_n327), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT69), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n340), .A2(new_n274), .A3(new_n328), .A4(new_n323), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT70), .B1(new_n341), .B2(KEYINPUT34), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(KEYINPUT34), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n336), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n330), .B(KEYINPUT32), .C1(new_n332), .C2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n341), .A2(KEYINPUT70), .A3(KEYINPUT34), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n337), .A2(new_n344), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n346), .A2(new_n337), .B1(new_n344), .B2(new_n347), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n273), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT72), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n346), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n344), .A2(new_n347), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(new_n348), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT72), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n356), .A2(new_n357), .A3(new_n273), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT71), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n353), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(new_n347), .A3(new_n344), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n353), .A2(new_n354), .A3(new_n359), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n361), .A2(KEYINPUT36), .A3(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n352), .A2(new_n358), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(G225gat), .A2(G233gat), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT2), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n367), .B1(G155gat), .B2(G162gat), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G148gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n370), .A2(G141gat), .ZN(new_n371));
  INV_X1    g170(.A(G141gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n372), .A2(G148gat), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n369), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G155gat), .B(G162gat), .ZN(new_n375));
  OR2_X1    g174(.A1(new_n375), .A2(KEYINPUT78), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(KEYINPUT78), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n374), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n375), .B(KEYINPUT81), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT79), .B(G148gat), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT80), .B1(new_n380), .B2(new_n372), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n381), .B1(G141gat), .B2(new_n370), .ZN(new_n382));
  NOR3_X1   g181(.A1(new_n380), .A2(KEYINPUT80), .A3(new_n372), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n369), .B(new_n379), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT82), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n384), .A2(new_n385), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n378), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n287), .B1(new_n388), .B2(KEYINPUT3), .ZN(new_n389));
  INV_X1    g188(.A(new_n378), .ZN(new_n390));
  OR2_X1    g189(.A1(new_n384), .A2(new_n385), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n384), .A2(new_n385), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n366), .B1(new_n389), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n393), .A2(new_n287), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT4), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n388), .A2(KEYINPUT83), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT83), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n401), .B(new_n378), .C1(new_n386), .C2(new_n387), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n400), .A2(KEYINPUT4), .A3(new_n287), .A4(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n396), .A2(new_n399), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT5), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n388), .A2(new_n327), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n397), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n405), .B1(new_n407), .B2(new_n366), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n397), .A2(KEYINPUT4), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n400), .A2(new_n287), .A3(new_n402), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n410), .B1(new_n411), .B2(KEYINPUT4), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n412), .A2(new_n405), .A3(new_n396), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G1gat), .B(G29gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(KEYINPUT0), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n416), .B(G57gat), .ZN(new_n417));
  INV_X1    g216(.A(G85gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n414), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT6), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n409), .A2(new_n413), .A3(new_n419), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n414), .A2(KEYINPUT6), .A3(new_n420), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(G226gat), .A2(G233gat), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n326), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n326), .B(KEYINPUT76), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AOI22_X1  g230(.A1(KEYINPUT73), .A2(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n432), .B1(KEYINPUT73), .B2(KEYINPUT22), .ZN(new_n433));
  XNOR2_X1  g232(.A(G211gat), .B(G218gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(G197gat), .B(G204gat), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT75), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n436), .B(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n433), .A2(new_n435), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT74), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n434), .B1(new_n439), .B2(new_n440), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n438), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OR2_X1    g243(.A1(new_n431), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(G8gat), .B(G36gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n446), .B(G64gat), .ZN(new_n447));
  INV_X1    g246(.A(G92gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n447), .B(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n326), .A2(new_n430), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n444), .B(new_n450), .C1(new_n429), .C2(new_n427), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n445), .A2(KEYINPUT30), .A3(new_n449), .A4(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n451), .B1(new_n431), .B2(new_n444), .ZN(new_n453));
  XOR2_X1   g252(.A(new_n449), .B(KEYINPUT77), .Z(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n451), .B(new_n449), .C1(new_n431), .C2(new_n444), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT30), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n452), .A2(new_n455), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n426), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(G22gat), .B(G50gat), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT29), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n464), .B1(new_n388), .B2(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(new_n444), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT84), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(G228gat), .A2(G233gat), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n465), .A2(KEYINPUT84), .A3(new_n444), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n400), .A2(new_n402), .ZN(new_n471));
  INV_X1    g270(.A(new_n434), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n438), .B1(new_n472), .B2(new_n439), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n394), .B1(new_n473), .B2(KEYINPUT29), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n468), .A2(new_n469), .A3(new_n470), .A4(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n444), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n477), .B1(new_n395), .B2(new_n464), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n464), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n393), .B1(new_n479), .B2(new_n394), .ZN(new_n480));
  OAI211_X1 g279(.A(G228gat), .B(G233gat), .C1(new_n478), .C2(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(G78gat), .B(G106gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n482), .B(KEYINPUT31), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n476), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n484), .B1(new_n476), .B2(new_n481), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n463), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n487), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n489), .A2(new_n462), .A3(new_n485), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n461), .A2(new_n491), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n364), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n477), .B(new_n450), .C1(new_n429), .C2(new_n427), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n494), .B(KEYINPUT37), .C1(new_n431), .C2(new_n477), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT37), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n451), .B(new_n496), .C1(new_n431), .C2(new_n444), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT38), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n454), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n495), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n500), .A2(new_n456), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n501), .A2(new_n424), .A3(new_n425), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT85), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT85), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n501), .A2(new_n424), .A3(new_n504), .A4(new_n425), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n449), .B1(new_n453), .B2(KEYINPUT37), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(new_n497), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT38), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n503), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n491), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT40), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n389), .A2(new_n395), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n365), .B1(new_n412), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT39), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT39), .B1(new_n407), .B2(new_n366), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n419), .B1(new_n513), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n511), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n513), .A2(new_n517), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n520), .A2(new_n515), .A3(KEYINPUT40), .A4(new_n419), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n519), .A2(new_n521), .A3(new_n421), .A4(new_n459), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n509), .A2(new_n510), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n493), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n459), .B1(new_n424), .B2(new_n425), .ZN(new_n525));
  INV_X1    g324(.A(new_n356), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT35), .ZN(new_n528));
  AND4_X1   g327(.A1(new_n490), .A2(new_n361), .A3(new_n488), .A4(new_n362), .ZN(new_n529));
  AOI211_X1 g328(.A(new_n528), .B(new_n459), .C1(new_n424), .C2(new_n425), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n527), .A2(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n272), .B1(new_n524), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT101), .ZN(new_n534));
  NAND2_X1  g333(.A1(G71gat), .A2(G78gat), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(G71gat), .A2(G78gat), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT88), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT9), .ZN(new_n539));
  AND3_X1   g338(.A1(new_n535), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n538), .B1(new_n535), .B2(new_n539), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OR2_X1    g341(.A1(G57gat), .A2(G64gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(G57gat), .A2(G64gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  AOI211_X1 g345(.A(new_n536), .B(new_n537), .C1(new_n542), .C2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT89), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n548), .B1(new_n540), .B2(new_n541), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n543), .B(new_n544), .C1(new_n536), .C2(new_n537), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n539), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT88), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n535), .A2(new_n538), .A3(new_n539), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(KEYINPUT89), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n549), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT90), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT90), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n549), .A2(new_n551), .A3(new_n555), .A4(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n547), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n258), .B1(new_n560), .B2(KEYINPUT21), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(G183gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(KEYINPUT92), .B(G211gat), .ZN(new_n565));
  INV_X1    g364(.A(G231gat), .ZN(new_n566));
  INV_X1    g365(.A(G233gat), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OR3_X1    g367(.A1(new_n560), .A2(KEYINPUT21), .A3(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G127gat), .B(G155gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT20), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n568), .B1(new_n560), .B2(KEYINPUT21), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n569), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n572), .B1(new_n569), .B2(new_n573), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n565), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n576), .ZN(new_n578));
  INV_X1    g377(.A(new_n565), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n578), .A2(new_n574), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n564), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n577), .A2(new_n580), .ZN(new_n582));
  INV_X1    g381(.A(new_n563), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n562), .B(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT93), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n587), .A2(G85gat), .A3(G92gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT7), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT7), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n587), .A2(new_n590), .A3(G85gat), .A4(G92gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT8), .ZN(new_n593));
  NOR2_X1   g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT95), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G99gat), .A2(G106gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AND2_X1   g397(.A1(KEYINPUT94), .A2(G92gat), .ZN(new_n599));
  NOR2_X1   g398(.A1(KEYINPUT94), .A2(G92gat), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(new_n418), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n592), .A2(new_n598), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n594), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n597), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n595), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  AOI22_X1  g407(.A1(new_n589), .A2(new_n591), .B1(new_n601), .B2(new_n418), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n609), .A2(new_n606), .A3(new_n598), .ZN(new_n610));
  AND3_X1   g409(.A1(new_n608), .A2(KEYINPUT96), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT96), .B1(new_n608), .B2(new_n610), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n613), .A2(new_n243), .A3(new_n254), .ZN(new_n614));
  XNOR2_X1  g413(.A(G190gat), .B(G218gat), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n257), .B1(new_n611), .B2(new_n612), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n614), .A2(new_n616), .A3(new_n617), .A4(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n619), .A2(KEYINPUT97), .ZN(new_n620));
  XNOR2_X1  g419(.A(G134gat), .B(G162gat), .ZN(new_n621));
  AOI21_X1  g420(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n614), .A2(new_n617), .A3(new_n618), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(new_n615), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n626), .A2(KEYINPUT97), .A3(new_n619), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n626), .A2(new_n619), .A3(new_n623), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT98), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n626), .A2(KEYINPUT98), .A3(new_n619), .A4(new_n623), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n628), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n586), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G176gat), .B(G204gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT100), .ZN(new_n636));
  XNOR2_X1  g435(.A(G120gat), .B(G148gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n636), .B(new_n637), .Z(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(G230gat), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n640), .A2(new_n567), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT10), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n608), .A2(new_n610), .A3(KEYINPUT99), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n606), .B1(new_n609), .B2(new_n598), .ZN(new_n645));
  AND4_X1   g444(.A1(new_n606), .A2(new_n592), .A3(new_n598), .A4(new_n602), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AND3_X1   g446(.A1(new_n560), .A2(new_n643), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n647), .B1(new_n560), .B2(new_n643), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n642), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n560), .A2(KEYINPUT10), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n613), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n641), .B1(new_n650), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n641), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n648), .A2(new_n649), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n639), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n547), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n550), .B1(new_n542), .B2(KEYINPUT89), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n558), .B1(new_n659), .B2(new_n549), .ZN(new_n660));
  INV_X1    g459(.A(new_n559), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n608), .A2(new_n610), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n662), .A2(new_n644), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n560), .A2(new_n643), .A3(new_n647), .ZN(new_n665));
  AOI21_X1  g464(.A(KEYINPUT10), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n655), .B1(new_n666), .B2(new_n652), .ZN(new_n667));
  INV_X1    g466(.A(new_n656), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(new_n668), .A3(new_n638), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n657), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n534), .B1(new_n634), .B2(new_n671), .ZN(new_n672));
  NOR4_X1   g471(.A1(new_n586), .A2(new_n633), .A3(KEYINPUT101), .A4(new_n670), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n533), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n426), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(G1gat), .ZN(G1324gat));
  INV_X1    g477(.A(KEYINPUT102), .ZN(new_n679));
  INV_X1    g478(.A(new_n674), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n532), .A2(new_n679), .A3(new_n459), .A4(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n510), .A2(new_n522), .ZN(new_n682));
  AOI22_X1  g481(.A1(new_n502), .A2(KEYINPUT85), .B1(KEYINPUT38), .B2(new_n507), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n682), .B1(new_n683), .B2(new_n505), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n364), .A2(new_n492), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n531), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n272), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n686), .A2(new_n459), .A3(new_n687), .A4(new_n680), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT102), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT16), .B(G8gat), .Z(new_n690));
  NAND3_X1  g489(.A1(new_n681), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT42), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(KEYINPUT103), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT103), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n691), .A2(new_n695), .A3(new_n692), .ZN(new_n696));
  INV_X1    g495(.A(new_n690), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n688), .A2(new_n692), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n681), .A2(new_n689), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n698), .B1(new_n699), .B2(G8gat), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n694), .A2(new_n696), .A3(new_n700), .ZN(G1325gat));
  AOI21_X1  g500(.A(G15gat), .B1(new_n675), .B2(new_n526), .ZN(new_n702));
  INV_X1    g501(.A(new_n364), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(G15gat), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT104), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n702), .B1(new_n675), .B2(new_n705), .ZN(G1326gat));
  NAND2_X1  g505(.A1(new_n675), .A2(new_n491), .ZN(new_n707));
  XNOR2_X1  g506(.A(KEYINPUT43), .B(G22gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(G1327gat));
  INV_X1    g508(.A(new_n586), .ZN(new_n710));
  INV_X1    g509(.A(new_n633), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n710), .A2(new_n711), .A3(new_n670), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n532), .A2(new_n232), .A3(new_n676), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT45), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n586), .B(KEYINPUT105), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n657), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n669), .B1(new_n269), .B2(new_n271), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n488), .A2(new_n490), .A3(new_n348), .A4(new_n355), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n528), .B1(new_n461), .B2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n510), .A2(new_n361), .A3(new_n362), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n525), .A2(KEYINPUT35), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n725), .B1(new_n493), .B2(new_n523), .ZN(new_n726));
  NOR2_X1   g525(.A1(KEYINPUT106), .A2(KEYINPUT44), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT106), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI22_X1  g529(.A1(new_n726), .A2(new_n711), .B1(new_n727), .B2(new_n730), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n686), .B(new_n633), .C1(new_n728), .C2(new_n729), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n720), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n733), .A2(new_n676), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n714), .B1(new_n734), .B2(new_n232), .ZN(G1328gat));
  NAND4_X1  g534(.A1(new_n532), .A2(new_n231), .A3(new_n459), .A4(new_n712), .ZN(new_n736));
  XOR2_X1   g535(.A(KEYINPUT107), .B(KEYINPUT46), .Z(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n733), .A2(new_n459), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n739), .B2(new_n231), .ZN(G1329gat));
  INV_X1    g539(.A(KEYINPUT47), .ZN(new_n741));
  INV_X1    g540(.A(new_n223), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n742), .B1(new_n733), .B2(new_n703), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n532), .A2(new_n526), .A3(new_n742), .A4(new_n712), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n741), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n726), .A2(new_n711), .A3(new_n730), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n730), .A2(new_n727), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n748), .B1(new_n686), .B2(new_n633), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n719), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n223), .B1(new_n750), .B2(new_n364), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n751), .A2(KEYINPUT47), .A3(new_n744), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n746), .A2(new_n752), .ZN(G1330gat));
  INV_X1    g552(.A(KEYINPUT48), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n216), .B1(new_n733), .B2(new_n491), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n510), .A2(G50gat), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n756), .A2(KEYINPUT108), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(KEYINPUT108), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n712), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n533), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n754), .B1(new_n755), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(G50gat), .B1(new_n750), .B2(new_n510), .ZN(new_n762));
  INV_X1    g561(.A(new_n760), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n762), .A2(KEYINPUT48), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n761), .A2(new_n764), .ZN(G1331gat));
  NAND3_X1  g564(.A1(new_n634), .A2(new_n272), .A3(new_n670), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n726), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n676), .ZN(new_n768));
  XOR2_X1   g567(.A(KEYINPUT109), .B(G57gat), .Z(new_n769));
  XNOR2_X1  g568(.A(new_n768), .B(new_n769), .ZN(G1332gat));
  NAND2_X1  g569(.A1(new_n767), .A2(new_n459), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n772));
  XOR2_X1   g571(.A(KEYINPUT49), .B(G64gat), .Z(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n771), .B2(new_n773), .ZN(G1333gat));
  XOR2_X1   g573(.A(new_n356), .B(KEYINPUT110), .Z(new_n775));
  AOI21_X1  g574(.A(G71gat), .B1(new_n767), .B2(new_n775), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n703), .A2(G71gat), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n776), .B1(new_n767), .B2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n778), .B(new_n779), .ZN(G1334gat));
  NAND2_X1  g579(.A1(new_n767), .A2(new_n491), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g581(.A1(new_n586), .A2(new_n272), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(KEYINPUT111), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n784), .A2(new_n671), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n786), .B1(new_n731), .B2(new_n732), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n787), .A2(new_n676), .ZN(new_n788));
  INV_X1    g587(.A(new_n784), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n686), .A2(new_n633), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n686), .A2(KEYINPUT51), .A3(new_n633), .A4(new_n789), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n676), .A2(new_n418), .A3(new_n670), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(KEYINPUT112), .ZN(new_n798));
  OAI22_X1  g597(.A1(new_n788), .A2(new_n418), .B1(new_n796), .B2(new_n798), .ZN(G1336gat));
  AOI21_X1  g598(.A(new_n601), .B1(new_n787), .B2(new_n459), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n460), .A2(G92gat), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  AOI211_X1 g601(.A(new_n671), .B(new_n802), .C1(new_n792), .C2(new_n794), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT52), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n601), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n785), .B1(new_n747), .B2(new_n749), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n805), .B1(new_n806), .B2(new_n460), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n670), .B(new_n801), .C1(new_n793), .C2(new_n795), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n804), .A2(new_n810), .ZN(G1337gat));
  OAI21_X1  g610(.A(G99gat), .B1(new_n806), .B2(new_n364), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n670), .B1(new_n793), .B2(new_n795), .ZN(new_n813));
  INV_X1    g612(.A(G99gat), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n526), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n812), .B1(new_n813), .B2(new_n815), .ZN(G1338gat));
  INV_X1    g615(.A(G106gat), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n817), .B1(new_n787), .B2(new_n491), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n510), .A2(G106gat), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  AOI211_X1 g619(.A(new_n671), .B(new_n820), .C1(new_n792), .C2(new_n794), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT53), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(G106gat), .B1(new_n806), .B2(new_n510), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n670), .B(new_n819), .C1(new_n793), .C2(new_n795), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n822), .A2(new_n826), .ZN(G1339gat));
  NAND3_X1  g626(.A1(new_n650), .A2(new_n653), .A3(new_n641), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n828), .A2(new_n667), .A3(KEYINPUT54), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n654), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n829), .A2(new_n831), .A3(KEYINPUT55), .A4(new_n639), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n270), .A2(new_n214), .A3(new_n263), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n256), .B1(new_n255), .B2(new_n259), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n259), .A2(new_n266), .A3(new_n265), .ZN(new_n835));
  INV_X1    g634(.A(new_n211), .ZN(new_n836));
  OAI22_X1  g635(.A1(new_n834), .A2(new_n835), .B1(new_n836), .B2(new_n209), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n654), .A2(new_n656), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n838), .B1(new_n839), .B2(new_n638), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n828), .A2(new_n667), .A3(KEYINPUT54), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n639), .B1(new_n667), .B2(KEYINPUT54), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n633), .A2(new_n832), .A3(new_n840), .A4(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n838), .B1(new_n657), .B2(new_n669), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n829), .A2(new_n831), .A3(new_n639), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n718), .B1(new_n841), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n846), .B1(new_n848), .B2(new_n832), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n845), .B1(new_n849), .B2(new_n633), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n715), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n634), .A2(new_n272), .A3(new_n671), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n426), .A2(new_n459), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n853), .A2(new_n510), .A3(new_n526), .A4(new_n854), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n855), .A2(new_n276), .A3(new_n272), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n426), .B1(new_n851), .B2(new_n852), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n857), .A2(new_n529), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n858), .A2(new_n460), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n687), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n856), .B1(new_n860), .B2(new_n276), .ZN(G1340gat));
  NOR3_X1   g660(.A1(new_n855), .A2(new_n277), .A3(new_n671), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n859), .A2(new_n670), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n863), .B2(new_n277), .ZN(G1341gat));
  NOR3_X1   g663(.A1(new_n855), .A2(new_n282), .A3(new_n715), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n859), .A2(new_n710), .ZN(new_n866));
  XOR2_X1   g665(.A(new_n866), .B(KEYINPUT113), .Z(new_n867));
  AOI21_X1  g666(.A(new_n865), .B1(new_n867), .B2(new_n282), .ZN(G1342gat));
  NAND2_X1  g667(.A1(new_n460), .A2(new_n633), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(KEYINPUT114), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n858), .A2(new_n281), .A3(new_n871), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n872), .A2(KEYINPUT56), .ZN(new_n873));
  OAI21_X1  g672(.A(G134gat), .B1(new_n855), .B2(new_n711), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(KEYINPUT56), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(G1343gat));
  AND3_X1   g675(.A1(new_n364), .A2(KEYINPUT115), .A3(new_n854), .ZN(new_n877));
  AOI21_X1  g676(.A(KEYINPUT115), .B1(new_n364), .B2(new_n854), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n850), .A2(new_n586), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n880), .A2(new_n852), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n491), .A2(KEYINPUT57), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n510), .B1(new_n851), .B2(new_n852), .ZN(new_n883));
  OAI22_X1  g682(.A1(new_n881), .A2(new_n882), .B1(new_n883), .B2(KEYINPUT57), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n879), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(G141gat), .B1(new_n885), .B2(new_n272), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n703), .A2(new_n510), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(new_n857), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n888), .A2(new_n459), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n372), .A3(new_n687), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT58), .ZN(G1344gat));
  OAI21_X1  g691(.A(new_n380), .B1(new_n885), .B2(new_n671), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n671), .A2(new_n380), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n889), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n879), .A2(new_n670), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n262), .A2(new_n263), .A3(new_n268), .ZN(new_n901));
  INV_X1    g700(.A(new_n214), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI22_X1  g702(.A1(new_n839), .A2(new_n638), .B1(new_n903), .B2(new_n833), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n844), .A2(new_n904), .A3(new_n832), .ZN(new_n905));
  INV_X1    g704(.A(new_n846), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n633), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AND4_X1   g706(.A1(new_n633), .A2(new_n832), .A3(new_n840), .A4(new_n844), .ZN(new_n908));
  OAI21_X1  g707(.A(KEYINPUT116), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT116), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n910), .B(new_n845), .C1(new_n849), .C2(new_n633), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n909), .A2(new_n911), .A3(new_n586), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT117), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n272), .B1(new_n672), .B2(new_n673), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n491), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n913), .B1(new_n912), .B2(new_n914), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n900), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n853), .A2(KEYINPUT57), .A3(new_n491), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n899), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(KEYINPUT118), .B1(new_n898), .B2(new_n922), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n920), .A2(new_n921), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT118), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n924), .A2(new_n925), .A3(new_n895), .A4(new_n897), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n923), .A2(new_n926), .ZN(G1345gat));
  OAI21_X1  g726(.A(G155gat), .B1(new_n885), .B2(new_n715), .ZN(new_n928));
  INV_X1    g727(.A(G155gat), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n889), .A2(new_n929), .A3(new_n710), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1346gat));
  OAI21_X1  g730(.A(G162gat), .B1(new_n885), .B2(new_n711), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n870), .A2(G162gat), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n888), .B2(new_n933), .ZN(G1347gat));
  NOR2_X1   g733(.A1(new_n676), .A2(new_n460), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n853), .A2(new_n529), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(G169gat), .B1(new_n936), .B2(new_n687), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n853), .A2(new_n935), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n938), .A2(new_n510), .A3(new_n775), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n272), .A2(new_n206), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  XOR2_X1   g740(.A(new_n941), .B(KEYINPUT119), .Z(G1348gat));
  NAND3_X1  g741(.A1(new_n936), .A2(new_n298), .A3(new_n670), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n939), .A2(new_n670), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n944), .B2(new_n298), .ZN(G1349gat));
  INV_X1    g744(.A(KEYINPUT120), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n939), .A2(new_n716), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n586), .A2(new_n313), .ZN(new_n948));
  AOI22_X1  g747(.A1(new_n947), .A2(G183gat), .B1(new_n936), .B2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT121), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n946), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(KEYINPUT60), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT60), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n953), .B1(new_n949), .B2(new_n946), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n952), .B1(new_n951), .B2(new_n954), .ZN(G1350gat));
  INV_X1    g754(.A(G190gat), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n936), .A2(new_n956), .A3(new_n633), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n939), .A2(new_n633), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(G190gat), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(KEYINPUT122), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT61), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT122), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n958), .A2(new_n962), .A3(G190gat), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n960), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n961), .B1(new_n960), .B2(new_n963), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n957), .B1(new_n964), .B2(new_n965), .ZN(G1351gat));
  AND2_X1   g765(.A1(new_n887), .A2(new_n938), .ZN(new_n967));
  XNOR2_X1  g766(.A(KEYINPUT123), .B(G197gat), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n967), .A2(new_n687), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n918), .A2(new_n919), .ZN(new_n970));
  XNOR2_X1  g769(.A(new_n970), .B(KEYINPUT124), .ZN(new_n971));
  INV_X1    g770(.A(new_n935), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n703), .A2(new_n972), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n971), .A2(new_n687), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n969), .B1(new_n974), .B2(new_n968), .ZN(G1352gat));
  XOR2_X1   g774(.A(KEYINPUT125), .B(G204gat), .Z(new_n976));
  NAND3_X1  g775(.A1(new_n967), .A2(new_n670), .A3(new_n976), .ZN(new_n977));
  XOR2_X1   g776(.A(new_n977), .B(KEYINPUT62), .Z(new_n978));
  AND3_X1   g777(.A1(new_n971), .A2(new_n670), .A3(new_n973), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n978), .B1(new_n979), .B2(new_n976), .ZN(G1353gat));
  INV_X1    g779(.A(G211gat), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n967), .A2(new_n981), .A3(new_n710), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n973), .A2(new_n710), .ZN(new_n983));
  INV_X1    g782(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n970), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g784(.A(KEYINPUT63), .B1(new_n985), .B2(G211gat), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n983), .B1(new_n918), .B2(new_n919), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT63), .ZN(new_n988));
  NOR3_X1   g787(.A1(new_n987), .A2(new_n988), .A3(new_n981), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n982), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT126), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI211_X1 g791(.A(KEYINPUT126), .B(new_n982), .C1(new_n986), .C2(new_n989), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n992), .A2(new_n993), .ZN(G1354gat));
  AOI21_X1  g793(.A(G218gat), .B1(new_n967), .B2(new_n633), .ZN(new_n995));
  XNOR2_X1  g794(.A(new_n995), .B(KEYINPUT127), .ZN(new_n996));
  AND3_X1   g795(.A1(new_n973), .A2(G218gat), .A3(new_n633), .ZN(new_n997));
  AOI21_X1  g796(.A(new_n996), .B1(new_n971), .B2(new_n997), .ZN(G1355gat));
endmodule


