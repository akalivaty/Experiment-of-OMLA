//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 0 1 1 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 0 0 0 0 0 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n823, new_n824, new_n825, new_n827, new_n828,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953;
  INV_X1    g000(.A(G64gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(G57gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(G57gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(KEYINPUT96), .B2(KEYINPUT9), .ZN(new_n206));
  NAND2_X1  g005(.A1(G71gat), .A2(G78gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT96), .ZN(new_n208));
  OR2_X1    g007(.A1(G71gat), .A2(G78gat), .ZN(new_n209));
  AND2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n206), .B(new_n210), .C1(KEYINPUT96), .C2(new_n207), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT97), .B(G57gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n204), .B1(new_n212), .B2(new_n202), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT9), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n207), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT21), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G231gat), .A2(G233gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n219), .B(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n221), .B(G127gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(G15gat), .B(G22gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G1gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G8gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT90), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n228), .B1(new_n223), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G22gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G15gat), .ZN(new_n232));
  INV_X1    g031(.A(G15gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G22gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n234), .A3(new_n229), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n235), .A2(G8gat), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n227), .B1(new_n230), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(G8gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n223), .A2(new_n229), .A3(new_n228), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n238), .A2(new_n239), .A3(new_n226), .A4(new_n225), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(new_n217), .B2(new_n218), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n222), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n244));
  INV_X1    g043(.A(G155gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(G183gat), .B(G211gat), .Z(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  OR2_X1    g048(.A1(new_n243), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n243), .A2(new_n249), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G190gat), .B(G218gat), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT7), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT98), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT98), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT7), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(G85gat), .A2(G92gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G99gat), .A2(G106gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT99), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT99), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n263), .A2(G99gat), .A3(G106gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n262), .A2(new_n264), .A3(KEYINPUT8), .ZN(new_n265));
  NOR2_X1   g064(.A1(G85gat), .A2(G92gat), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G85gat), .ZN(new_n268));
  INV_X1    g067(.A(G92gat), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n270), .A2(new_n255), .A3(new_n257), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n260), .A2(new_n265), .A3(new_n267), .A4(new_n271), .ZN(new_n272));
  XOR2_X1   g071(.A(G99gat), .B(G106gat), .Z(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT98), .B(KEYINPUT7), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n266), .B1(new_n275), .B2(new_n270), .ZN(new_n276));
  INV_X1    g075(.A(new_n273), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n276), .A2(new_n277), .A3(new_n265), .A4(new_n260), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT15), .ZN(new_n281));
  OR2_X1    g080(.A1(G43gat), .A2(G50gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(G43gat), .A2(G50gat), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G29gat), .ZN(new_n285));
  INV_X1    g084(.A(G36gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(new_n286), .A3(KEYINPUT14), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT14), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n288), .B1(G29gat), .B2(G36gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT89), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G29gat), .A2(G36gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n290), .B1(new_n287), .B2(new_n289), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n284), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n284), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n287), .A2(new_n289), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n282), .A2(new_n281), .A3(new_n283), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n296), .A2(new_n297), .A3(new_n292), .A4(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT17), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT17), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n295), .A2(new_n302), .A3(new_n299), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n280), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G232gat), .A2(G233gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT41), .ZN(new_n307));
  AND2_X1   g106(.A1(new_n295), .A2(new_n299), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n307), .B1(new_n308), .B2(new_n279), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n253), .B1(new_n304), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT100), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n306), .A2(KEYINPUT41), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n312), .B(G134gat), .ZN(new_n313));
  INV_X1    g112(.A(G162gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n313), .B(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  OR3_X1    g115(.A1(new_n304), .A2(new_n253), .A3(new_n309), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(new_n310), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n316), .A2(new_n318), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G230gat), .A2(G233gat), .ZN(new_n323));
  AND2_X1   g122(.A1(new_n211), .A2(new_n216), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n277), .B1(new_n272), .B2(KEYINPUT101), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT102), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT101), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n276), .A2(new_n327), .A3(new_n265), .A4(new_n260), .ZN(new_n328));
  AND3_X1   g127(.A1(new_n325), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n325), .A2(new_n328), .B1(new_n326), .B2(new_n278), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n324), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n280), .A2(new_n217), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT10), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT10), .ZN(new_n334));
  NOR3_X1   g133(.A1(new_n217), .A2(new_n279), .A3(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n323), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G120gat), .B(G148gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(G176gat), .B(G204gat), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n337), .B(new_n338), .Z(new_n339));
  INV_X1    g138(.A(new_n323), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n331), .A2(new_n340), .A3(new_n332), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT103), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n331), .A2(KEYINPUT103), .A3(new_n340), .A4(new_n332), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n336), .A2(new_n339), .A3(new_n343), .A4(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT104), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AND2_X1   g146(.A1(new_n343), .A2(new_n344), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n348), .A2(KEYINPUT104), .A3(new_n339), .A4(new_n336), .ZN(new_n349));
  INV_X1    g148(.A(new_n339), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n336), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n347), .A2(new_n349), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n252), .A2(new_n322), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(G228gat), .A2(G233gat), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT3), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n356));
  OR2_X1    g155(.A1(G197gat), .A2(G204gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(G197gat), .A2(G204gat), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  XOR2_X1   g160(.A(G211gat), .B(G218gat), .Z(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n359), .A2(new_n360), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n362), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n355), .B1(new_n368), .B2(KEYINPUT29), .ZN(new_n369));
  XOR2_X1   g168(.A(G141gat), .B(G148gat), .Z(new_n370));
  OAI21_X1  g169(.A(KEYINPUT2), .B1(new_n245), .B2(new_n314), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(G155gat), .B(G162gat), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n370), .A2(new_n373), .A3(new_n371), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n354), .B1(new_n369), .B2(new_n377), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n375), .A2(new_n376), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(new_n355), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT77), .B(KEYINPUT29), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(KEYINPUT81), .A3(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n381), .B1(new_n377), .B2(KEYINPUT3), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT81), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n382), .A2(new_n368), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT82), .ZN(new_n387));
  AND2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n386), .A2(new_n387), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n378), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n367), .A2(new_n381), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n379), .B1(new_n391), .B2(new_n355), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n367), .B1(new_n380), .B2(new_n381), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n354), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n390), .A2(new_n231), .A3(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n231), .B1(new_n390), .B2(new_n394), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT83), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n390), .A2(new_n394), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(G22gat), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT83), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n400), .A2(new_n401), .A3(new_n395), .ZN(new_n402));
  XNOR2_X1  g201(.A(G78gat), .B(G106gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT31), .B(G50gat), .ZN(new_n404));
  XOR2_X1   g203(.A(new_n403), .B(new_n404), .Z(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n398), .A2(new_n402), .A3(new_n406), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n400), .A2(new_n401), .A3(new_n395), .A4(new_n405), .ZN(new_n408));
  AND2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT78), .ZN(new_n410));
  NAND2_X1  g209(.A1(G169gat), .A2(G176gat), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT26), .ZN(new_n412));
  NOR2_X1   g211(.A1(G169gat), .A2(G176gat), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n413), .A2(KEYINPUT70), .A3(new_n412), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT70), .B1(new_n413), .B2(new_n412), .ZN(new_n415));
  OAI221_X1 g214(.A(new_n411), .B1(new_n412), .B2(new_n413), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(G183gat), .A2(G190gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT71), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n416), .A2(KEYINPUT71), .A3(new_n417), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT27), .B(G183gat), .ZN(new_n422));
  INV_X1    g221(.A(G190gat), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(KEYINPUT28), .A3(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT69), .B(G183gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT27), .ZN(new_n426));
  OR2_X1    g225(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n427));
  AOI21_X1  g226(.A(G190gat), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n424), .B1(new_n428), .B2(KEYINPUT28), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n420), .A2(new_n421), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n413), .A2(KEYINPUT23), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n411), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT66), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n432), .B(new_n433), .ZN(new_n434));
  AND2_X1   g233(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n435));
  NOR2_X1   g234(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n436));
  OAI22_X1  g235(.A1(new_n435), .A2(new_n436), .B1(G169gat), .B2(G176gat), .ZN(new_n437));
  XOR2_X1   g236(.A(KEYINPUT69), .B(G183gat), .Z(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n423), .ZN(new_n439));
  XOR2_X1   g238(.A(KEYINPUT67), .B(KEYINPUT24), .Z(new_n440));
  AOI22_X1  g239(.A1(new_n439), .A2(new_n440), .B1(G183gat), .B2(G190gat), .ZN(new_n441));
  NAND3_X1  g240(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n442));
  XOR2_X1   g241(.A(new_n442), .B(KEYINPUT68), .Z(new_n443));
  OAI211_X1 g242(.A(new_n434), .B(new_n437), .C1(new_n441), .C2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT25), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT64), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n431), .A2(new_n446), .ZN(new_n447));
  AOI211_X1 g246(.A(KEYINPUT25), .B(new_n447), .C1(G169gat), .C2(G176gat), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT24), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n417), .A2(new_n449), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n450), .B(new_n442), .C1(G183gat), .C2(G190gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n431), .A2(new_n446), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n448), .A2(new_n451), .A3(new_n437), .A4(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n430), .A2(new_n445), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(G226gat), .A2(G233gat), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT29), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n457), .B(new_n367), .C1(new_n459), .C2(new_n456), .ZN(new_n460));
  INV_X1    g259(.A(new_n457), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n456), .B1(new_n454), .B2(new_n381), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n368), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(G8gat), .B(G36gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(G64gat), .B(G92gat), .ZN(new_n466));
  XOR2_X1   g265(.A(new_n465), .B(new_n466), .Z(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n410), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  AOI211_X1 g268(.A(KEYINPUT78), .B(new_n467), .C1(new_n460), .C2(new_n463), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n464), .A2(new_n468), .ZN(new_n471));
  OAI22_X1  g270(.A1(new_n469), .A2(new_n470), .B1(new_n471), .B2(KEYINPUT30), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n460), .A2(new_n463), .A3(KEYINPUT30), .A4(new_n467), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(KEYINPUT79), .ZN(new_n474));
  XOR2_X1   g273(.A(G1gat), .B(G29gat), .Z(new_n475));
  XNOR2_X1  g274(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n475), .B(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G57gat), .B(G85gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n477), .B(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(G127gat), .ZN(new_n480));
  INV_X1    g279(.A(G134gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(G113gat), .B(G120gat), .ZN(new_n483));
  XOR2_X1   g282(.A(KEYINPUT72), .B(G127gat), .Z(new_n484));
  OAI221_X1 g283(.A(new_n482), .B1(new_n483), .B2(KEYINPUT1), .C1(new_n484), .C2(new_n481), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(KEYINPUT73), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT1), .ZN(new_n487));
  XNOR2_X1  g286(.A(G127gat), .B(G134gat), .ZN(new_n488));
  INV_X1    g287(.A(G113gat), .ZN(new_n489));
  OR3_X1    g288(.A1(new_n489), .A2(KEYINPUT73), .A3(G120gat), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n486), .A2(new_n487), .A3(new_n488), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n485), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n379), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n493), .A2(KEYINPUT4), .A3(new_n379), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(G225gat), .A2(G233gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n377), .A2(KEYINPUT3), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n380), .A2(new_n492), .A3(new_n500), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n498), .A2(KEYINPUT5), .A3(new_n499), .A4(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n496), .A2(new_n501), .A3(new_n497), .ZN(new_n503));
  INV_X1    g302(.A(new_n499), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n492), .A2(new_n377), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n499), .B1(new_n494), .B2(new_n506), .ZN(new_n507));
  OAI22_X1  g306(.A1(new_n503), .A2(new_n504), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n479), .B1(new_n502), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT6), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n502), .A2(new_n508), .A3(new_n479), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n512), .A2(new_n511), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR3_X1   g314(.A1(new_n472), .A2(new_n474), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n454), .A2(new_n493), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n430), .A2(new_n445), .A3(new_n492), .A4(new_n453), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n517), .A2(G227gat), .A3(G233gat), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT32), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT33), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  XOR2_X1   g321(.A(G15gat), .B(G43gat), .Z(new_n523));
  XNOR2_X1  g322(.A(G71gat), .B(G99gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n520), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n525), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n519), .B(KEYINPUT32), .C1(new_n521), .C2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n517), .A2(new_n518), .ZN(new_n530));
  NAND2_X1  g329(.A1(G227gat), .A2(G233gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT34), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT74), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n533), .B1(new_n531), .B2(new_n534), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n532), .A2(new_n535), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n529), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n526), .A2(new_n536), .A3(new_n537), .A4(new_n528), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n409), .A2(new_n516), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT35), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n512), .A2(new_n511), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT85), .B1(new_n545), .B2(new_n509), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT85), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n510), .A2(new_n547), .A3(new_n511), .A4(new_n512), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n546), .A2(new_n548), .A3(new_n514), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT35), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR3_X1   g350(.A1(new_n551), .A2(new_n472), .A3(new_n474), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n539), .A2(KEYINPUT75), .A3(new_n540), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT75), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n529), .A2(new_n538), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT87), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT87), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n553), .A2(new_n558), .A3(new_n555), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n552), .A2(new_n557), .A3(new_n409), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n461), .A2(new_n462), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(new_n367), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n456), .B1(new_n454), .B2(new_n458), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n368), .B1(new_n461), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n565), .A3(KEYINPUT86), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT37), .ZN(new_n567));
  NOR3_X1   g366(.A1(new_n461), .A2(new_n462), .A3(new_n368), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT86), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT38), .B1(new_n566), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n468), .B1(new_n464), .B2(KEYINPUT37), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n471), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n549), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n567), .B1(new_n460), .B2(new_n463), .ZN(new_n576));
  OAI21_X1  g375(.A(KEYINPUT38), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n574), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n503), .A2(new_n504), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n494), .A2(new_n499), .A3(new_n506), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(KEYINPUT39), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n479), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n581), .B(new_n582), .C1(KEYINPUT39), .C2(new_n579), .ZN(new_n583));
  NOR2_X1   g382(.A1(KEYINPUT84), .A2(KEYINPUT40), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n584), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n585), .A2(new_n512), .A3(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n587), .B1(new_n472), .B2(new_n474), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n409), .A2(new_n578), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n474), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n469), .A2(new_n470), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n513), .A2(new_n514), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n471), .A2(KEYINPUT30), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n590), .A2(new_n591), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n407), .A2(new_n408), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n542), .A2(KEYINPUT36), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT36), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n553), .A2(new_n598), .A3(new_n555), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n589), .A2(new_n596), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n561), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G113gat), .B(G141gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(G169gat), .B(G197gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(KEYINPUT88), .B(KEYINPUT11), .Z(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT12), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT91), .ZN(new_n610));
  AND3_X1   g409(.A1(new_n295), .A2(new_n302), .A3(new_n299), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n302), .B1(new_n295), .B2(new_n299), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n610), .B(new_n241), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n237), .A2(new_n240), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n614), .B1(new_n301), .B2(new_n303), .ZN(new_n615));
  OAI21_X1  g414(.A(KEYINPUT91), .B1(new_n308), .B2(new_n241), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n613), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT92), .ZN(new_n618));
  NAND2_X1  g417(.A1(G229gat), .A2(G233gat), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n617), .A2(new_n618), .A3(KEYINPUT18), .A4(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n308), .B(new_n241), .ZN(new_n621));
  XNOR2_X1  g420(.A(KEYINPUT93), .B(KEYINPUT13), .ZN(new_n622));
  INV_X1    g421(.A(new_n619), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n241), .B1(new_n611), .B2(new_n612), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n610), .B1(new_n614), .B2(new_n300), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n623), .B1(new_n628), .B2(new_n613), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n620), .B(new_n625), .C1(KEYINPUT18), .C2(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n618), .B1(new_n629), .B2(KEYINPUT18), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n609), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT94), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n619), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT18), .ZN(new_n635));
  AOI22_X1  g434(.A1(new_n634), .A2(new_n635), .B1(new_n621), .B2(new_n624), .ZN(new_n636));
  OAI21_X1  g435(.A(KEYINPUT92), .B1(new_n634), .B2(new_n635), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n636), .A2(new_n637), .A3(new_n620), .A4(new_n608), .ZN(new_n638));
  AND3_X1   g437(.A1(new_n632), .A2(new_n633), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n633), .B1(new_n632), .B2(new_n638), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n602), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT95), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT95), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n602), .A2(new_n644), .A3(new_n641), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n353), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n515), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g447(.A1(new_n472), .A2(new_n474), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g450(.A(KEYINPUT16), .B(G8gat), .Z(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n228), .B1(new_n646), .B2(new_n650), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT42), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n656), .B1(KEYINPUT42), .B2(new_n654), .ZN(G1325gat));
  AND2_X1   g456(.A1(new_n557), .A2(new_n559), .ZN(new_n658));
  AOI21_X1  g457(.A(G15gat), .B1(new_n646), .B2(new_n658), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n659), .A2(KEYINPUT105), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(KEYINPUT105), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n600), .A2(new_n233), .ZN(new_n662));
  AOI22_X1  g461(.A1(new_n660), .A2(new_n661), .B1(new_n646), .B2(new_n662), .ZN(G1326gat));
  NAND2_X1  g462(.A1(new_n646), .A2(new_n595), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT43), .B(G22gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(G1327gat));
  INV_X1    g465(.A(KEYINPUT45), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n347), .A2(new_n349), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n351), .A2(new_n350), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n252), .A2(new_n322), .A3(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n672), .B1(new_n643), .B2(new_n645), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n515), .A2(new_n285), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n667), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n673), .A2(KEYINPUT45), .A3(new_n285), .A4(new_n515), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n321), .A2(KEYINPUT44), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n650), .A2(new_n595), .A3(new_n551), .ZN(new_n679));
  AOI22_X1  g478(.A1(new_n658), .A2(new_n679), .B1(new_n543), .B2(KEYINPUT35), .ZN(new_n680));
  INV_X1    g479(.A(new_n601), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n678), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n632), .A2(new_n638), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n252), .A2(new_n684), .A3(new_n670), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT106), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n686), .B1(new_n409), .B2(new_n516), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n594), .A2(new_n595), .A3(KEYINPUT106), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n687), .A2(new_n589), .A3(new_n688), .A4(new_n600), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n322), .B1(new_n561), .B2(new_n689), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n682), .B(new_n685), .C1(new_n690), .C2(KEYINPUT44), .ZN(new_n691));
  OAI21_X1  g490(.A(G29gat), .B1(new_n691), .B2(new_n592), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n676), .A2(new_n677), .A3(new_n692), .ZN(G1328gat));
  NOR2_X1   g492(.A1(new_n649), .A2(G36gat), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  OR3_X1    g494(.A1(new_n674), .A2(KEYINPUT46), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(G36gat), .B1(new_n691), .B2(new_n649), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT46), .B1(new_n674), .B2(new_n695), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(G1329gat));
  NOR2_X1   g498(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n700));
  INV_X1    g499(.A(new_n658), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n701), .A2(G43gat), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n700), .B1(new_n673), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(G43gat), .B1(new_n691), .B2(new_n600), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1330gat));
  OAI21_X1  g506(.A(G50gat), .B1(new_n691), .B2(new_n409), .ZN(new_n708));
  INV_X1    g507(.A(G50gat), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n595), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n708), .B1(new_n674), .B2(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT108), .B(KEYINPUT48), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1331gat));
  NAND4_X1  g512(.A1(new_n252), .A2(new_n684), .A3(new_n322), .A4(new_n670), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n714), .B1(new_n561), .B2(new_n689), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n515), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(new_n212), .ZN(G1332gat));
  AOI21_X1  g516(.A(new_n649), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g518(.A(new_n719), .B(KEYINPUT109), .Z(new_n720));
  NOR2_X1   g519(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1333gat));
  XOR2_X1   g521(.A(new_n658), .B(KEYINPUT110), .Z(new_n723));
  AOI21_X1  g522(.A(G71gat), .B1(new_n723), .B2(new_n715), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n597), .A2(new_n599), .A3(G71gat), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n724), .B1(new_n715), .B2(new_n725), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n726), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g526(.A1(new_n715), .A2(new_n595), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g528(.A1(new_n252), .A2(new_n683), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n731), .A2(new_n352), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n682), .B(new_n732), .C1(new_n690), .C2(KEYINPUT44), .ZN(new_n733));
  OAI21_X1  g532(.A(G85gat), .B1(new_n733), .B2(new_n592), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n690), .A2(KEYINPUT51), .A3(new_n730), .ZN(new_n735));
  AOI21_X1  g534(.A(KEYINPUT51), .B1(new_n690), .B2(new_n730), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n670), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n515), .A2(new_n268), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n734), .B1(new_n737), .B2(new_n738), .ZN(G1336gat));
  OAI21_X1  g538(.A(G92gat), .B1(new_n733), .B2(new_n649), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n650), .A2(new_n269), .A3(new_n670), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT111), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n735), .B2(new_n736), .ZN(new_n743));
  XNOR2_X1  g542(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n740), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT51), .ZN(new_n746));
  AOI211_X1 g545(.A(new_n322), .B(new_n731), .C1(new_n561), .C2(new_n689), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n746), .B1(new_n747), .B2(KEYINPUT112), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n690), .A2(new_n730), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n749), .A2(new_n750), .A3(KEYINPUT51), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n748), .A2(new_n751), .A3(new_n742), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n752), .A2(new_n740), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754));
  OAI211_X1 g553(.A(KEYINPUT114), .B(new_n745), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT114), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n740), .A2(new_n743), .A3(new_n744), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n754), .B1(new_n752), .B2(new_n740), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n755), .A2(new_n759), .ZN(G1337gat));
  OAI21_X1  g559(.A(G99gat), .B1(new_n733), .B2(new_n600), .ZN(new_n761));
  OR2_X1    g560(.A1(new_n701), .A2(G99gat), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n761), .B1(new_n737), .B2(new_n762), .ZN(G1338gat));
  OAI21_X1  g562(.A(G106gat), .B1(new_n733), .B2(new_n409), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n751), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n409), .A2(G106gat), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n670), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n764), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(KEYINPUT53), .ZN(new_n769));
  XNOR2_X1  g568(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n770));
  INV_X1    g569(.A(new_n766), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n764), .B(new_n770), .C1(new_n737), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n769), .A2(new_n772), .ZN(G1339gat));
  INV_X1    g572(.A(new_n252), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n272), .A2(KEYINPUT101), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n775), .A2(new_n273), .A3(new_n328), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n278), .A2(new_n326), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n325), .A2(new_n326), .A3(new_n328), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n217), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n324), .A2(new_n279), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n334), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n335), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n782), .A2(new_n340), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT116), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT116), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n782), .A2(new_n786), .A3(new_n340), .A4(new_n783), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n785), .A2(KEYINPUT54), .A3(new_n336), .A4(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n340), .B1(new_n782), .B2(new_n783), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT54), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n339), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n788), .A2(KEYINPUT55), .A3(new_n791), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n668), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n788), .A2(new_n791), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT117), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT117), .ZN(new_n797));
  AOI211_X1 g596(.A(new_n797), .B(KEYINPUT55), .C1(new_n788), .C2(new_n791), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n793), .B(new_n683), .C1(new_n796), .C2(new_n798), .ZN(new_n799));
  OAI22_X1  g598(.A1(new_n617), .A2(new_n619), .B1(new_n621), .B2(new_n624), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n607), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n638), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n670), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n321), .B1(new_n799), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n322), .A2(new_n802), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n793), .B(new_n806), .C1(new_n796), .C2(new_n798), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n774), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n353), .A2(new_n683), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n592), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n409), .A2(new_n542), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n812), .A2(new_n650), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(G113gat), .B1(new_n815), .B2(new_n683), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n595), .B1(new_n809), .B2(new_n810), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n650), .A2(new_n592), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n817), .A2(new_n658), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n641), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n819), .A2(new_n489), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n816), .A2(new_n821), .ZN(G1340gat));
  AOI21_X1  g621(.A(G120gat), .B1(new_n815), .B2(new_n670), .ZN(new_n823));
  INV_X1    g622(.A(G120gat), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n819), .A2(new_n824), .A3(new_n352), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n823), .A2(new_n825), .ZN(G1341gat));
  NAND3_X1  g625(.A1(new_n815), .A2(new_n484), .A3(new_n252), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n819), .A2(new_n774), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n827), .B1(new_n484), .B2(new_n828), .ZN(G1342gat));
  NOR3_X1   g628(.A1(new_n814), .A2(G134gat), .A3(new_n322), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  OR2_X1    g630(.A1(new_n831), .A2(KEYINPUT56), .ZN(new_n832));
  OAI21_X1  g631(.A(G134gat), .B1(new_n819), .B2(new_n322), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(KEYINPUT56), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(G1343gat));
  INV_X1    g634(.A(KEYINPUT58), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n600), .A2(new_n595), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n837), .A2(new_n650), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n811), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(G141gat), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n839), .A2(new_n840), .A3(new_n641), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n818), .A2(new_n600), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n595), .A2(KEYINPUT57), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n794), .A2(new_n795), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n844), .B1(new_n639), .B2(new_n640), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n668), .A2(new_n792), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n670), .A2(new_n848), .A3(new_n803), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT118), .B1(new_n352), .B2(new_n802), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n322), .B1(new_n847), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n252), .B1(new_n852), .B2(new_n807), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n843), .B1(new_n854), .B2(new_n810), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n809), .A2(new_n810), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT57), .B1(new_n856), .B2(new_n595), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n842), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(KEYINPUT119), .B1(new_n858), .B2(new_n820), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(G141gat), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n858), .A2(KEYINPUT119), .A3(new_n820), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n836), .B(new_n841), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(G141gat), .B1(new_n858), .B2(new_n684), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n841), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(KEYINPUT58), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n862), .A2(new_n865), .ZN(G1344gat));
  INV_X1    g665(.A(G148gat), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n867), .A2(KEYINPUT59), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n868), .B1(new_n858), .B2(new_n352), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n843), .B1(new_n809), .B2(new_n810), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n353), .A2(new_n641), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n595), .B1(new_n853), .B2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n870), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n842), .A2(new_n670), .ZN(new_n875));
  OAI21_X1  g674(.A(G148gat), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n877));
  XOR2_X1   g676(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n878));
  AND3_X1   g677(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n877), .B1(new_n876), .B2(new_n878), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n869), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n839), .A2(new_n867), .A3(new_n670), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(G1345gat));
  OAI21_X1  g682(.A(G155gat), .B1(new_n858), .B2(new_n774), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n839), .A2(new_n245), .A3(new_n252), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(G1346gat));
  OAI21_X1  g685(.A(G162gat), .B1(new_n858), .B2(new_n322), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n839), .A2(new_n314), .A3(new_n321), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(G1347gat));
  NAND2_X1  g688(.A1(new_n650), .A2(new_n592), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n890), .B(KEYINPUT122), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n723), .A2(new_n817), .A3(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(G169gat), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n892), .A2(new_n893), .A3(new_n820), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n515), .B1(new_n809), .B2(new_n810), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n812), .A2(new_n649), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(G169gat), .B1(new_n898), .B2(new_n683), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n894), .A2(new_n899), .ZN(G1348gat));
  OAI21_X1  g699(.A(G176gat), .B1(new_n892), .B2(new_n352), .ZN(new_n901));
  OR2_X1    g700(.A1(new_n352), .A2(G176gat), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n897), .B2(new_n902), .ZN(G1349gat));
  OAI21_X1  g702(.A(new_n425), .B1(new_n892), .B2(new_n774), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n898), .A2(new_n422), .A3(new_n252), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g706(.A1(new_n898), .A2(new_n423), .A3(new_n321), .ZN(new_n908));
  OAI21_X1  g707(.A(G190gat), .B1(new_n892), .B2(new_n322), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n909), .A2(KEYINPUT61), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n909), .A2(KEYINPUT61), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(G1351gat));
  NOR2_X1   g711(.A1(new_n837), .A2(new_n649), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n895), .A2(new_n913), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n914), .A2(G197gat), .A3(new_n684), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n891), .A2(new_n600), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n874), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n641), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n915), .B1(new_n918), .B2(G197gat), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT123), .ZN(G1352gat));
  NOR3_X1   g719(.A1(new_n914), .A2(G204gat), .A3(new_n352), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT62), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n917), .A2(new_n670), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(G204gat), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT124), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n922), .A2(new_n924), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n928), .ZN(G1353gat));
  OR3_X1    g728(.A1(new_n914), .A2(G211gat), .A3(new_n774), .ZN(new_n930));
  INV_X1    g729(.A(new_n916), .ZN(new_n931));
  OAI211_X1 g730(.A(new_n850), .B(new_n849), .C1(new_n845), .C2(new_n846), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n808), .B1(new_n322), .B2(new_n932), .ZN(new_n933));
  OAI22_X1  g732(.A1(new_n933), .A2(new_n252), .B1(new_n641), .B2(new_n353), .ZN(new_n934));
  AOI21_X1  g733(.A(KEYINPUT57), .B1(new_n934), .B2(new_n595), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n252), .B(new_n931), .C1(new_n935), .C2(new_n870), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n936), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n937));
  AOI21_X1  g736(.A(KEYINPUT63), .B1(new_n936), .B2(G211gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n930), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT125), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI211_X1 g740(.A(KEYINPUT125), .B(new_n930), .C1(new_n937), .C2(new_n938), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(G1354gat));
  INV_X1    g742(.A(KEYINPUT127), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT126), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n945), .B1(new_n874), .B2(new_n916), .ZN(new_n946));
  OAI211_X1 g745(.A(KEYINPUT126), .B(new_n931), .C1(new_n935), .C2(new_n870), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n946), .A2(new_n321), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(G218gat), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n914), .A2(G218gat), .A3(new_n322), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n944), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  AOI211_X1 g751(.A(KEYINPUT127), .B(new_n950), .C1(new_n948), .C2(G218gat), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n952), .A2(new_n953), .ZN(G1355gat));
endmodule


