//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 1 1 0 0 0 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0 0 0 0 1 1 0 0 1 1 1 1 0 0 1 0 0 1 0 0 0 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n188));
  INV_X1    g002(.A(G140), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G125), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(G125), .ZN(new_n191));
  INV_X1    g005(.A(G125), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G140), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n190), .B1(new_n194), .B2(new_n188), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n195), .B(G146), .ZN(new_n196));
  NOR2_X1   g010(.A1(G237), .A2(G953), .ZN(new_n197));
  AND3_X1   g011(.A1(new_n197), .A2(G143), .A3(G214), .ZN(new_n198));
  AOI21_X1  g012(.A(G143), .B1(new_n197), .B2(G214), .ZN(new_n199));
  OAI211_X1 g013(.A(KEYINPUT17), .B(G131), .C1(new_n198), .C2(new_n199), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n198), .A2(new_n199), .ZN(new_n201));
  INV_X1    g015(.A(G131), .ZN(new_n202));
  XNOR2_X1  g016(.A(new_n201), .B(new_n202), .ZN(new_n203));
  OAI211_X1 g017(.A(new_n196), .B(new_n200), .C1(new_n203), .C2(KEYINPUT17), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT18), .A2(G131), .ZN(new_n205));
  XOR2_X1   g019(.A(new_n201), .B(new_n205), .Z(new_n206));
  NAND2_X1  g020(.A1(new_n194), .A2(KEYINPUT73), .ZN(new_n207));
  XNOR2_X1  g021(.A(G125), .B(G140), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT73), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n207), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n212), .B1(new_n211), .B2(new_n208), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n206), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(G113), .B(G122), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT89), .B(G104), .ZN(new_n216));
  XOR2_X1   g030(.A(new_n215), .B(new_n216), .Z(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n204), .A2(new_n214), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n218), .B1(new_n204), .B2(new_n214), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n187), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT90), .B(G475), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT20), .ZN(new_n225));
  NOR2_X1   g039(.A1(G475), .A2(G902), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT19), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n207), .A2(new_n210), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n194), .A2(KEYINPUT19), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(new_n211), .A3(new_n229), .ZN(new_n230));
  OAI211_X1 g044(.A(G146), .B(new_n190), .C1(new_n194), .C2(new_n188), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT88), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT88), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n230), .A2(new_n234), .A3(new_n231), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n233), .A2(new_n203), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n218), .B1(new_n236), .B2(new_n214), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n225), .B(new_n226), .C1(new_n237), .C2(new_n220), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n201), .B(G131), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n240), .B1(new_n232), .B2(KEYINPUT88), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n241), .A2(new_n235), .B1(new_n213), .B2(new_n206), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n219), .B1(new_n242), .B2(new_n218), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n225), .B1(new_n243), .B2(new_n226), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n224), .B1(new_n239), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT91), .ZN(new_n246));
  INV_X1    g060(.A(G116), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n246), .B1(new_n247), .B2(G122), .ZN(new_n248));
  INV_X1    g062(.A(G122), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(KEYINPUT91), .A3(G116), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT92), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n247), .A2(G122), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n252), .B1(new_n251), .B2(new_n253), .ZN(new_n256));
  INV_X1    g070(.A(G107), .ZN(new_n257));
  NOR3_X1   g071(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n251), .A2(new_n253), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT92), .ZN(new_n260));
  AOI21_X1  g074(.A(G107), .B1(new_n260), .B2(new_n254), .ZN(new_n261));
  OAI21_X1  g075(.A(KEYINPUT93), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n257), .B1(new_n255), .B2(new_n256), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n260), .A2(G107), .A3(new_n254), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT93), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(G128), .B(G143), .ZN(new_n267));
  INV_X1    g081(.A(G134), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n269), .B(KEYINPUT94), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n267), .A2(KEYINPUT13), .ZN(new_n271));
  INV_X1    g085(.A(G128), .ZN(new_n272));
  NOR3_X1   g086(.A1(new_n272), .A2(KEYINPUT13), .A3(G143), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(new_n268), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n270), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n262), .A2(new_n266), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n253), .A2(KEYINPUT14), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n251), .A2(KEYINPUT95), .A3(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n278), .B1(KEYINPUT14), .B2(new_n253), .ZN(new_n279));
  AOI21_X1  g093(.A(KEYINPUT95), .B1(new_n251), .B2(new_n277), .ZN(new_n280));
  OAI21_X1  g094(.A(G107), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n267), .B(new_n268), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n263), .A3(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT9), .B(G234), .ZN(new_n284));
  INV_X1    g098(.A(G217), .ZN(new_n285));
  NOR3_X1   g099(.A1(new_n284), .A2(new_n285), .A3(G953), .ZN(new_n286));
  AND3_X1   g100(.A1(new_n276), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n286), .B1(new_n276), .B2(new_n283), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n187), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G478), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n290), .A2(KEYINPUT15), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  OAI221_X1 g106(.A(new_n187), .B1(KEYINPUT15), .B2(new_n290), .C1(new_n287), .C2(new_n288), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(G234), .A2(G237), .ZN(new_n295));
  INV_X1    g109(.A(G953), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n295), .A2(G952), .A3(new_n296), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n295), .A2(G902), .A3(G953), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT21), .B(G898), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n245), .A2(new_n294), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(G214), .B1(G237), .B2(G902), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT86), .ZN(new_n303));
  XNOR2_X1  g117(.A(G116), .B(G119), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT2), .B(G113), .ZN(new_n305));
  XOR2_X1   g119(.A(new_n304), .B(new_n305), .Z(new_n306));
  INV_X1    g120(.A(KEYINPUT3), .ZN(new_n307));
  INV_X1    g121(.A(G104), .ZN(new_n308));
  AOI22_X1  g122(.A1(KEYINPUT76), .A2(new_n307), .B1(new_n308), .B2(G107), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT76), .ZN(new_n310));
  AND4_X1   g124(.A1(new_n310), .A2(new_n257), .A3(KEYINPUT3), .A4(G104), .ZN(new_n311));
  AOI22_X1  g125(.A1(new_n310), .A2(KEYINPUT3), .B1(new_n257), .B2(G104), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n309), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT4), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n314), .A3(G101), .ZN(new_n315));
  OAI22_X1  g129(.A1(new_n310), .A2(KEYINPUT3), .B1(new_n257), .B2(G104), .ZN(new_n316));
  OAI22_X1  g130(.A1(KEYINPUT76), .A2(new_n307), .B1(new_n308), .B2(G107), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n310), .A2(new_n257), .A3(KEYINPUT3), .A4(G104), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G101), .ZN(new_n320));
  OAI21_X1  g134(.A(KEYINPUT4), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n320), .B(new_n309), .C1(new_n311), .C2(new_n312), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n306), .B(new_n315), .C1(new_n321), .C2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n257), .A2(G104), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n308), .A2(G107), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n320), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n327), .B1(new_n319), .B2(new_n320), .ZN(new_n328));
  INV_X1    g142(.A(new_n304), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n329), .A2(new_n305), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT5), .ZN(new_n332));
  INV_X1    g146(.A(G119), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(new_n333), .A3(G116), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT82), .ZN(new_n335));
  OR2_X1    g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n304), .A2(KEYINPUT5), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n334), .A2(new_n335), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n336), .A2(new_n337), .A3(G113), .A4(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n328), .A2(new_n331), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n324), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(G110), .B(G122), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n324), .A2(new_n340), .A3(new_n342), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(KEYINPUT6), .A3(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n272), .A2(KEYINPUT1), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n211), .A2(G143), .ZN(new_n348));
  INV_X1    g162(.A(G143), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G146), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n347), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n348), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(KEYINPUT64), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT64), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(new_n349), .A3(G146), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n352), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n272), .B1(new_n348), .B2(KEYINPUT1), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n192), .B(new_n351), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n354), .B1(new_n349), .B2(G146), .ZN(new_n359));
  NOR3_X1   g173(.A1(new_n211), .A2(KEYINPUT64), .A3(G143), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n348), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AND2_X1   g175(.A1(KEYINPUT0), .A2(G128), .ZN(new_n362));
  NOR2_X1   g176(.A1(KEYINPUT0), .A2(G128), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(G143), .B(G146), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n361), .A2(new_n364), .B1(new_n365), .B2(new_n362), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n358), .B(KEYINPUT83), .C1(new_n366), .C2(new_n192), .ZN(new_n367));
  INV_X1    g181(.A(G224), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(G953), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n369), .B(KEYINPUT84), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n365), .A2(new_n362), .ZN(new_n371));
  INV_X1    g185(.A(new_n364), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n371), .B1(new_n356), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT83), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(G125), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n367), .A2(new_n370), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n370), .B1(new_n367), .B2(new_n375), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT6), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n341), .A2(new_n379), .A3(new_n343), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n346), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n327), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n322), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(new_n331), .A3(new_n339), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n342), .B(KEYINPUT8), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT85), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n386), .B1(new_n304), .B2(KEYINPUT5), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n333), .A2(G116), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n247), .A2(G119), .ZN(new_n389));
  AND4_X1   g203(.A1(new_n386), .A2(new_n388), .A3(new_n389), .A4(KEYINPUT5), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(G113), .B1(new_n334), .B2(new_n335), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n392), .B1(new_n335), .B2(new_n334), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n330), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n384), .B(new_n385), .C1(new_n394), .C2(new_n383), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n358), .B1(new_n366), .B2(new_n192), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT7), .B1(new_n368), .B2(G953), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n345), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n397), .B1(new_n367), .B2(new_n375), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n187), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n303), .B1(new_n381), .B2(new_n401), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n345), .A2(new_n395), .A3(new_n398), .ZN(new_n403));
  INV_X1    g217(.A(new_n400), .ZN(new_n404));
  AOI21_X1  g218(.A(G902), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n346), .A2(new_n378), .A3(new_n380), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT86), .ZN(new_n407));
  OAI21_X1  g221(.A(G210), .B1(G237), .B2(G902), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n402), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n405), .A2(new_n406), .A3(new_n408), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT87), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n402), .A2(KEYINPUT87), .A3(new_n407), .A4(new_n409), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n301), .A2(new_n302), .A3(new_n415), .A4(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT81), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n351), .B1(new_n357), .B2(new_n365), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n322), .A2(new_n419), .A3(new_n382), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT10), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT77), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n366), .B(new_n315), .C1(new_n321), .C2(new_n323), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n351), .B1(new_n356), .B2(new_n357), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n328), .A2(new_n426), .A3(KEYINPUT10), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n420), .A2(KEYINPUT77), .A3(new_n421), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n424), .A2(new_n425), .A3(new_n427), .A4(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT66), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT65), .ZN(new_n431));
  INV_X1    g245(.A(G137), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AND2_X1   g247(.A1(KEYINPUT11), .A2(G134), .ZN(new_n434));
  NAND2_X1  g248(.A1(KEYINPUT65), .A2(G137), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(KEYINPUT11), .A2(G134), .ZN(new_n437));
  NOR2_X1   g251(.A1(KEYINPUT11), .A2(G134), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n437), .B1(new_n438), .B2(G137), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n436), .A2(new_n202), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n202), .B1(new_n436), .B2(new_n439), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n430), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n436), .A2(new_n439), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(G131), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n436), .A2(new_n439), .A3(new_n202), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(KEYINPUT66), .A3(new_n445), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n429), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT79), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n429), .A2(new_n450), .A3(new_n447), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n450), .B1(new_n429), .B2(new_n447), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n449), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(G110), .B(G140), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n296), .A2(G227), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n420), .B1(new_n328), .B2(new_n426), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n444), .A2(new_n445), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(KEYINPUT12), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT78), .ZN(new_n461));
  AOI211_X1 g275(.A(new_n461), .B(KEYINPUT12), .C1(new_n447), .C2(new_n458), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n458), .A2(new_n446), .A3(new_n442), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT12), .ZN(new_n464));
  AOI21_X1  g278(.A(KEYINPUT78), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n460), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n456), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n467), .B1(new_n429), .B2(new_n447), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(G902), .B1(new_n457), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT80), .B(G469), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n467), .B1(new_n466), .B2(new_n449), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n429), .A2(new_n447), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT79), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n429), .A2(new_n450), .A3(new_n447), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n468), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n187), .B1(new_n474), .B2(new_n478), .ZN(new_n479));
  AOI22_X1  g293(.A1(new_n471), .A2(new_n473), .B1(new_n479), .B2(G469), .ZN(new_n480));
  INV_X1    g294(.A(G221), .ZN(new_n481));
  INV_X1    g295(.A(new_n284), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n481), .B1(new_n482), .B2(new_n187), .ZN(new_n483));
  XOR2_X1   g297(.A(new_n483), .B(KEYINPUT75), .Z(new_n484));
  OAI21_X1  g298(.A(new_n418), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n484), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n479), .A2(G469), .ZN(new_n487));
  AOI22_X1  g301(.A1(new_n453), .A2(new_n456), .B1(new_n466), .B2(new_n469), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n488), .A2(G902), .A3(new_n472), .ZN(new_n489));
  OAI211_X1 g303(.A(KEYINPUT81), .B(new_n486), .C1(new_n487), .C2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n417), .B1(new_n485), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT70), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n442), .A2(new_n446), .A3(new_n366), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n433), .A2(new_n268), .A3(new_n435), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n202), .B1(G134), .B2(G137), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n445), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n426), .ZN(new_n498));
  INV_X1    g312(.A(new_n306), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n493), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT28), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT28), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n493), .A2(new_n502), .A3(new_n498), .A4(new_n499), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n440), .A2(new_n441), .ZN(new_n505));
  INV_X1    g319(.A(new_n357), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n361), .A2(new_n506), .B1(new_n365), .B2(new_n347), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n445), .A2(new_n496), .ZN(new_n508));
  OAI22_X1  g322(.A1(new_n505), .A2(new_n373), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n306), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  XOR2_X1   g325(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n512));
  NAND2_X1  g326(.A1(new_n197), .A2(G210), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT26), .B(G101), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n514), .B(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n516), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n500), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT31), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT30), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n499), .B1(new_n509), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT67), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n493), .A2(KEYINPUT30), .A3(new_n498), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n524), .B1(new_n523), .B2(new_n525), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n520), .B(new_n521), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n517), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT69), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n493), .A2(KEYINPUT30), .A3(new_n498), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n366), .A2(new_n459), .B1(new_n497), .B2(new_n426), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n306), .B1(new_n532), .B2(KEYINPUT30), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT67), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n519), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n530), .B1(new_n536), .B2(new_n521), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n520), .B1(new_n526), .B2(new_n527), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n538), .A2(KEYINPUT69), .A3(KEYINPUT31), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n529), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(G472), .A2(G902), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT32), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n493), .A2(new_n498), .ZN(new_n546));
  AOI22_X1  g360(.A1(new_n501), .A2(new_n503), .B1(new_n546), .B2(new_n306), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT29), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n516), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(G902), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n500), .B1(new_n526), .B2(new_n527), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n516), .ZN(new_n553));
  AOI22_X1  g367(.A1(new_n501), .A2(new_n503), .B1(new_n306), .B2(new_n509), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT29), .B1(new_n554), .B2(new_n518), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n551), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(G472), .ZN(new_n557));
  OAI22_X1  g371(.A1(new_n540), .A2(new_n545), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n536), .A2(new_n521), .B1(new_n516), .B2(new_n511), .ZN(new_n559));
  NOR3_X1   g373(.A1(new_n536), .A2(new_n530), .A3(new_n521), .ZN(new_n560));
  AOI21_X1  g374(.A(KEYINPUT69), .B1(new_n538), .B2(KEYINPUT31), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(KEYINPUT32), .B1(new_n562), .B2(new_n541), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n492), .B1(new_n558), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n534), .A2(new_n535), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n518), .B1(new_n565), .B2(new_n500), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n548), .B1(new_n511), .B2(new_n516), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n550), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n562), .A2(new_n544), .B1(G472), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n543), .B1(new_n540), .B2(new_n542), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(KEYINPUT70), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n564), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n285), .B1(G234), .B2(new_n187), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  XOR2_X1   g388(.A(G119), .B(G128), .Z(new_n575));
  XNOR2_X1  g389(.A(KEYINPUT24), .B(G110), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT71), .ZN(new_n578));
  OAI211_X1 g392(.A(G119), .B(new_n272), .C1(new_n578), .C2(KEYINPUT23), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT23), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n580), .B1(new_n333), .B2(G128), .ZN(new_n581));
  OAI21_X1  g395(.A(KEYINPUT71), .B1(new_n333), .B2(G128), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n579), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n577), .B1(new_n583), .B2(G110), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(new_n231), .A3(new_n212), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT74), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n585), .B(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n575), .A2(new_n576), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n196), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n583), .A2(G110), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(KEYINPUT72), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n587), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(KEYINPUT22), .B(G137), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n296), .A2(G221), .A3(G234), .ZN(new_n595));
  XOR2_X1   g409(.A(new_n594), .B(new_n595), .Z(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n587), .A2(new_n592), .A3(new_n596), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(new_n187), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT25), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n598), .A2(KEYINPUT25), .A3(new_n187), .A4(new_n599), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n574), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n598), .A2(new_n599), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n605), .A2(G902), .A3(new_n573), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n491), .A2(new_n572), .A3(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(G101), .ZN(G3));
  OAI21_X1  g423(.A(G472), .B1(new_n540), .B2(G902), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n562), .A2(new_n541), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n612), .B1(new_n485), .B2(new_n490), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n613), .A2(new_n607), .ZN(new_n614));
  INV_X1    g428(.A(new_n302), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n409), .B1(new_n381), .B2(new_n401), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n615), .B1(new_n616), .B2(new_n411), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(new_n300), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT33), .B1(new_n286), .B2(KEYINPUT96), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n287), .A2(new_n288), .A3(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n620), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n276), .A2(new_n283), .ZN(new_n623));
  INV_X1    g437(.A(new_n286), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n276), .A2(new_n283), .A3(new_n286), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n622), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(G478), .B1(new_n621), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n290), .A2(new_n187), .ZN(new_n629));
  AOI21_X1  g443(.A(G902), .B1(new_n625), .B2(new_n626), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n629), .B1(new_n630), .B2(new_n290), .ZN(new_n631));
  AOI21_X1  g445(.A(KEYINPUT97), .B1(new_n628), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n620), .B1(new_n287), .B2(new_n288), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n625), .A2(new_n626), .A3(new_n622), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n290), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n290), .B(new_n187), .C1(new_n287), .C2(new_n288), .ZN(new_n636));
  INV_X1    g450(.A(new_n629), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT97), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n635), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n245), .B1(new_n632), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(KEYINPUT98), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n628), .A2(KEYINPUT97), .A3(new_n631), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n639), .B1(new_n635), .B2(new_n638), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT98), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n645), .A2(new_n646), .A3(new_n245), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n614), .A2(new_n619), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT34), .B(G104), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G6));
  NOR2_X1   g465(.A1(new_n237), .A2(new_n220), .ZN(new_n652));
  INV_X1    g466(.A(new_n226), .ZN(new_n653));
  OAI21_X1  g467(.A(KEYINPUT20), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  AOI22_X1  g468(.A1(new_n654), .A2(new_n238), .B1(new_n222), .B2(new_n223), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n294), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n618), .A2(new_n656), .A3(new_n300), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n614), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT99), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT35), .B(G107), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G9));
  NAND2_X1  g475(.A1(new_n602), .A2(new_n603), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n573), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT100), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n587), .A2(new_n664), .A3(new_n592), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n664), .B1(new_n587), .B2(new_n592), .ZN(new_n667));
  OAI22_X1  g481(.A1(new_n666), .A2(new_n667), .B1(KEYINPUT36), .B2(new_n597), .ZN(new_n668));
  INV_X1    g482(.A(new_n667), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n597), .A2(KEYINPUT36), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n669), .A2(new_n670), .A3(new_n665), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n573), .A2(G902), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n668), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n663), .A2(new_n674), .A3(KEYINPUT101), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT101), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n676), .B1(new_n604), .B2(new_n673), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n417), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n613), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT37), .B(G110), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G12));
  AOI211_X1 g496(.A(new_n618), .B(new_n678), .C1(new_n485), .C2(new_n490), .ZN(new_n683));
  INV_X1    g497(.A(G900), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n298), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n297), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n655), .A2(new_n294), .A3(new_n687), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n688), .B(KEYINPUT102), .Z(new_n689));
  NAND3_X1  g503(.A1(new_n683), .A2(new_n572), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G128), .ZN(G30));
  NAND2_X1  g505(.A1(new_n485), .A2(new_n490), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  XOR2_X1   g507(.A(new_n687), .B(KEYINPUT39), .Z(new_n694));
  OR2_X1    g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g509(.A1(new_n695), .A2(KEYINPUT40), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(KEYINPUT40), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n604), .A2(new_n673), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT86), .ZN(new_n699));
  AOI21_X1  g513(.A(KEYINPUT86), .B1(new_n405), .B2(new_n406), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n699), .A2(new_n700), .A3(new_n408), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n416), .B1(new_n701), .B2(new_n413), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n703));
  XOR2_X1   g517(.A(new_n702), .B(new_n703), .Z(new_n704));
  NAND2_X1  g518(.A1(new_n552), .A2(new_n518), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n546), .A2(new_n306), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n500), .A2(new_n516), .ZN(new_n708));
  AOI211_X1 g522(.A(G902), .B(new_n706), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  OAI221_X1 g523(.A(new_n570), .B1(new_n557), .B2(new_n709), .C1(new_n540), .C2(new_n545), .ZN(new_n710));
  INV_X1    g524(.A(new_n294), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n711), .A2(new_n655), .A3(new_n615), .ZN(new_n712));
  AND4_X1   g526(.A1(new_n698), .A2(new_n704), .A3(new_n710), .A4(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n696), .A2(new_n697), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G143), .ZN(G45));
  INV_X1    g529(.A(new_n687), .ZN(new_n716));
  AOI211_X1 g530(.A(new_n655), .B(new_n716), .C1(new_n643), .C2(new_n644), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n683), .A2(new_n572), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G146), .ZN(G48));
  OAI21_X1  g533(.A(G469), .B1(new_n488), .B2(G902), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n476), .A2(new_n477), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n467), .B1(new_n721), .B2(new_n449), .ZN(new_n722));
  INV_X1    g536(.A(new_n470), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n187), .B(new_n473), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n483), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n725), .A2(new_n607), .A3(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n572), .A2(new_n648), .A3(new_n619), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(KEYINPUT41), .B(G113), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(G15));
  AND3_X1   g544(.A1(new_n569), .A2(KEYINPUT70), .A3(new_n570), .ZN(new_n731));
  AOI21_X1  g545(.A(KEYINPUT70), .B1(new_n569), .B2(new_n570), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n727), .B(new_n657), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G116), .ZN(G18));
  NAND4_X1  g548(.A1(new_n720), .A2(new_n724), .A3(new_n617), .A4(new_n726), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n300), .ZN(new_n736));
  AND4_X1   g550(.A1(new_n711), .A2(new_n675), .A3(new_n655), .A4(new_n677), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n736), .B(new_n737), .C1(new_n731), .C2(new_n732), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G119), .ZN(G21));
  AOI21_X1  g553(.A(new_n557), .B1(new_n562), .B2(new_n187), .ZN(new_n740));
  INV_X1    g554(.A(new_n607), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n547), .A2(new_n518), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n742), .B1(new_n521), .B2(new_n536), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n538), .A2(KEYINPUT31), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n542), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n740), .A2(new_n741), .A3(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n746), .A2(new_n736), .A3(new_n294), .A4(new_n245), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G122), .ZN(G24));
  NOR3_X1   g562(.A1(new_n740), .A2(new_n698), .A3(new_n745), .ZN(new_n749));
  INV_X1    g563(.A(new_n735), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n717), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G125), .ZN(G27));
  AOI21_X1  g566(.A(new_n615), .B1(new_n415), .B2(new_n416), .ZN(new_n753));
  NAND2_X1  g567(.A1(G469), .A2(G902), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(KEYINPUT104), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n474), .A2(new_n478), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n755), .B1(new_n756), .B2(G469), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n483), .B1(new_n757), .B2(new_n724), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n717), .A2(KEYINPUT42), .A3(new_n753), .A4(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(KEYINPUT105), .B1(new_n540), .B2(new_n545), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT105), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n562), .A2(new_n761), .A3(new_n544), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n568), .A2(G472), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n570), .A2(new_n760), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n607), .ZN(new_n765));
  OAI21_X1  g579(.A(KEYINPUT106), .B1(new_n759), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n758), .A2(new_n302), .A3(new_n702), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n645), .A2(KEYINPUT42), .A3(new_n245), .A4(new_n687), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT106), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n769), .A2(new_n770), .A3(new_n607), .A4(new_n764), .ZN(new_n771));
  INV_X1    g585(.A(new_n767), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n572), .A2(new_n607), .A3(new_n717), .A4(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT42), .ZN(new_n774));
  AOI22_X1  g588(.A1(new_n766), .A2(new_n771), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(new_n202), .ZN(G33));
  NAND4_X1  g590(.A1(new_n572), .A2(new_n689), .A3(new_n607), .A4(new_n772), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  AOI21_X1  g592(.A(new_n245), .B1(new_n645), .B2(KEYINPUT108), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n779), .B1(KEYINPUT108), .B2(new_n645), .ZN(new_n780));
  XNOR2_X1  g594(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT109), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n655), .B(KEYINPUT110), .ZN(new_n784));
  INV_X1    g598(.A(new_n645), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT43), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n698), .B1(new_n610), .B2(new_n611), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT44), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n788), .A2(KEYINPUT44), .A3(new_n789), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n756), .A2(KEYINPUT45), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n756), .A2(KEYINPUT45), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(G469), .A3(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n755), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT46), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n489), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n800), .B1(new_n799), .B2(new_n798), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n726), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n802), .A2(new_n694), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n792), .A2(new_n753), .A3(new_n793), .A4(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G137), .ZN(G39));
  NAND3_X1  g619(.A1(new_n717), .A2(new_n741), .A3(new_n753), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n572), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n801), .A2(KEYINPUT47), .A3(new_n726), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT47), .B1(new_n801), .B2(new_n726), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n807), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT111), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(KEYINPUT111), .B(new_n807), .C1(new_n809), .C2(new_n810), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G140), .ZN(G42));
  AND3_X1   g630(.A1(new_n690), .A2(new_n718), .A3(new_n751), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n616), .A2(new_n411), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n712), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n698), .A2(new_n726), .A3(new_n687), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n821), .B1(new_n724), .B2(new_n757), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n710), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n817), .A2(new_n818), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n690), .A2(new_n718), .A3(new_n751), .A4(new_n823), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT52), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n300), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n415), .A2(new_n302), .A3(new_n416), .A4(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n829), .B1(new_n641), .B2(new_n656), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n613), .A2(new_n607), .A3(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n608), .A2(new_n680), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT112), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n741), .B1(new_n564), .B2(new_n571), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n834), .A2(new_n491), .B1(new_n613), .B2(new_n679), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT112), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n835), .A2(new_n836), .A3(new_n831), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n766), .A2(new_n771), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n773), .A2(new_n774), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n728), .A2(new_n733), .A3(new_n738), .A4(new_n747), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n702), .A2(new_n302), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n843), .A2(new_n716), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n572), .A2(new_n692), .A3(new_n737), .A4(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n772), .A2(new_n717), .A3(new_n749), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n777), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n842), .A2(new_n847), .ZN(new_n848));
  AND4_X1   g662(.A1(KEYINPUT113), .A2(new_n838), .A3(new_n841), .A4(new_n848), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n775), .A2(new_n842), .A3(new_n847), .ZN(new_n850));
  AOI21_X1  g664(.A(KEYINPUT113), .B1(new_n850), .B2(new_n838), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n827), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n818), .B1(new_n690), .B2(new_n751), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n855), .A2(KEYINPUT53), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n854), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(KEYINPUT54), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n832), .A2(KEYINPUT112), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n836), .B1(new_n835), .B2(new_n831), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n727), .B1(new_n731), .B2(new_n732), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n646), .B1(new_n645), .B2(new_n245), .ZN(new_n864));
  AOI211_X1 g678(.A(KEYINPUT98), .B(new_n655), .C1(new_n643), .C2(new_n644), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n619), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n747), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n733), .A2(new_n738), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n777), .A2(new_n845), .A3(new_n846), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n841), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n862), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n855), .A2(new_n853), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n827), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n824), .A2(new_n826), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT113), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n876), .B1(new_n862), .B2(new_n871), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n850), .A2(KEYINPUT113), .A3(new_n838), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n859), .B(new_n874), .C1(new_n879), .C2(KEYINPUT53), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n858), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n686), .B1(new_n783), .B2(new_n787), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n725), .A2(new_n726), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n704), .A2(new_n302), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n882), .A2(new_n746), .A3(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT50), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n885), .B(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n810), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n486), .B1(new_n725), .B2(KEYINPUT114), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n889), .B1(KEYINPUT114), .B2(new_n725), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n888), .A2(new_n808), .A3(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n882), .A2(new_n891), .A3(new_n746), .A4(new_n753), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n883), .A2(new_n843), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n882), .A2(new_n749), .A3(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n710), .A2(new_n741), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n895), .A2(new_n297), .A3(new_n893), .ZN(new_n896));
  OR3_X1    g710(.A1(new_n896), .A2(new_n245), .A3(new_n645), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n892), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n887), .B(new_n899), .C1(KEYINPUT115), .C2(KEYINPUT51), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n887), .A2(new_n899), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n892), .A2(new_n894), .A3(KEYINPUT115), .A4(new_n897), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT51), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n648), .ZN(new_n906));
  OAI211_X1 g720(.A(G952), .B(new_n296), .C1(new_n896), .C2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n765), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n882), .A2(new_n908), .A3(new_n893), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT48), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT48), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n882), .A2(new_n911), .A3(new_n908), .A4(new_n893), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n907), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT117), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n882), .A2(new_n750), .A3(new_n746), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT116), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n882), .A2(KEYINPUT116), .A3(new_n750), .A4(new_n746), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n913), .A2(new_n914), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n914), .B1(new_n913), .B2(new_n919), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n900), .B(new_n905), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  OAI22_X1  g736(.A1(new_n881), .A2(new_n922), .B1(G952), .B2(G953), .ZN(new_n923));
  INV_X1    g737(.A(new_n704), .ZN(new_n924));
  NOR4_X1   g738(.A1(new_n784), .A2(new_n785), .A3(new_n484), .A4(new_n615), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n725), .B(KEYINPUT49), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n895), .A2(new_n924), .A3(new_n925), .A4(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n923), .A2(new_n927), .ZN(G75));
  OAI21_X1  g742(.A(new_n874), .B1(new_n879), .B2(KEYINPUT53), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n929), .A2(G210), .A3(G902), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT56), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n346), .A2(new_n380), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(new_n378), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT55), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n930), .A2(new_n931), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n934), .B1(new_n930), .B2(new_n931), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n296), .A2(G952), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(G51));
  INV_X1    g752(.A(KEYINPUT118), .ZN(new_n939));
  INV_X1    g753(.A(new_n929), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n940), .A2(new_n187), .A3(new_n796), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n755), .B(KEYINPUT57), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n859), .B1(new_n854), .B2(new_n874), .ZN(new_n943));
  INV_X1    g757(.A(new_n880), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n488), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n941), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n939), .B1(new_n947), .B2(new_n937), .ZN(new_n948));
  INV_X1    g762(.A(new_n937), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n929), .A2(KEYINPUT54), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n880), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n488), .B1(new_n951), .B2(new_n942), .ZN(new_n952));
  OAI211_X1 g766(.A(KEYINPUT118), .B(new_n949), .C1(new_n952), .C2(new_n941), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n948), .A2(new_n953), .ZN(G54));
  NAND4_X1  g768(.A1(new_n929), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n955));
  OR3_X1    g769(.A1(new_n955), .A2(KEYINPUT119), .A3(new_n652), .ZN(new_n956));
  OAI21_X1  g770(.A(KEYINPUT119), .B1(new_n955), .B2(new_n652), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n937), .B1(new_n955), .B2(new_n652), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(G60));
  NOR2_X1   g773(.A1(new_n621), .A2(new_n627), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n629), .B(KEYINPUT59), .Z(new_n961));
  AOI21_X1  g775(.A(new_n960), .B1(new_n881), .B2(new_n961), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n951), .A2(new_n960), .A3(new_n961), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n962), .A2(new_n937), .A3(new_n963), .ZN(G63));
  XOR2_X1   g778(.A(new_n605), .B(KEYINPUT120), .Z(new_n965));
  NAND2_X1  g779(.A1(G217), .A2(G902), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT60), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n965), .B1(new_n940), .B2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n967), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n929), .A2(new_n671), .A3(new_n668), .A4(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n968), .A2(new_n949), .A3(new_n970), .ZN(new_n971));
  XNOR2_X1  g785(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n971), .B(new_n972), .Z(G66));
  NAND2_X1  g787(.A1(new_n838), .A2(new_n869), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n296), .ZN(new_n975));
  OAI21_X1  g789(.A(G953), .B1(new_n299), .B2(new_n368), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n975), .A2(KEYINPUT122), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n977), .B1(KEYINPUT122), .B2(new_n975), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n932), .B1(G898), .B2(new_n296), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n978), .B(new_n979), .Z(G69));
  OAI21_X1  g794(.A(new_n525), .B1(KEYINPUT30), .B2(new_n532), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n228), .A2(new_n229), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(new_n982), .ZN(new_n983));
  AOI211_X1 g797(.A(new_n843), .B(new_n695), .C1(new_n641), .C2(new_n656), .ZN(new_n984));
  AOI22_X1  g798(.A1(new_n813), .A2(new_n814), .B1(new_n834), .B2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n714), .ZN(new_n986));
  OR2_X1    g800(.A1(new_n817), .A2(KEYINPUT123), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n817), .A2(KEYINPUT123), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT62), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n804), .B(new_n985), .C1(new_n989), .C2(new_n990), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n989), .A2(new_n990), .ZN(new_n992));
  OR2_X1    g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n983), .B1(new_n993), .B2(new_n296), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n296), .B1(G227), .B2(G900), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n987), .A2(new_n988), .ZN(new_n996));
  INV_X1    g810(.A(new_n777), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n908), .A2(new_n820), .ZN(new_n998));
  AOI211_X1 g812(.A(new_n997), .B(new_n775), .C1(new_n803), .C2(new_n998), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n804), .A2(new_n815), .A3(new_n996), .A4(new_n999), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n1000), .A2(G953), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n983), .B1(new_n684), .B2(new_n296), .ZN(new_n1002));
  OAI21_X1  g816(.A(KEYINPUT124), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  OR3_X1    g817(.A1(new_n994), .A2(new_n995), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n995), .B1(new_n994), .B2(new_n1003), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(G72));
  NOR3_X1   g820(.A1(new_n991), .A2(new_n992), .A3(new_n974), .ZN(new_n1007));
  NAND2_X1  g821(.A1(G472), .A2(G902), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT63), .Z(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT125), .Z(new_n1010));
  OAI21_X1  g824(.A(new_n706), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n536), .B1(new_n553), .B2(KEYINPUT126), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1012), .B1(KEYINPUT126), .B2(new_n553), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n857), .A2(new_n1009), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1010), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1015), .B1(new_n1000), .B2(new_n974), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n552), .A2(new_n518), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n937), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1011), .A2(new_n1014), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT127), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n1011), .A2(KEYINPUT127), .A3(new_n1014), .A4(new_n1018), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1021), .A2(new_n1022), .ZN(G57));
endmodule


