//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n854, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962;
  INV_X1    g000(.A(G8gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n204));
  AND2_X1   g003(.A1(G15gat), .A2(G22gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(G15gat), .A2(G22gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n202), .B1(new_n207), .B2(KEYINPUT91), .ZN(new_n208));
  XNOR2_X1  g007(.A(G15gat), .B(G22gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n207), .B1(new_n209), .B2(G1gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT92), .ZN(new_n212));
  OAI221_X1 g011(.A(new_n207), .B1(KEYINPUT91), .B2(new_n202), .C1(new_n209), .C2(G1gat), .ZN(new_n213));
  AND3_X1   g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n212), .B1(new_n211), .B2(new_n213), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI211_X1 g015(.A(KEYINPUT89), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(G29gat), .A2(G36gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT14), .ZN(new_n219));
  INV_X1    g018(.A(G29gat), .ZN(new_n220));
  INV_X1    g019(.A(G36gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n217), .B(new_n218), .C1(new_n224), .C2(KEYINPUT89), .ZN(new_n225));
  XNOR2_X1  g024(.A(G43gat), .B(G50gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT15), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  XOR2_X1   g028(.A(G43gat), .B(G50gat), .Z(new_n230));
  INV_X1    g029(.A(KEYINPUT15), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n232), .A2(new_n224), .A3(new_n227), .A4(new_n218), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n229), .A2(new_n233), .A3(KEYINPUT17), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT90), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n229), .A2(new_n233), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT17), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  AOI211_X1 g037(.A(KEYINPUT90), .B(KEYINPUT17), .C1(new_n229), .C2(new_n233), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n216), .B(new_n234), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G229gat), .A2(G233gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n211), .A2(new_n213), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n236), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n240), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT18), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT93), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n247), .B1(new_n236), .B2(new_n242), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(new_n243), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n241), .B(KEYINPUT13), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n240), .A2(KEYINPUT18), .A3(new_n241), .A4(new_n243), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n246), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G113gat), .B(G141gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(G169gat), .B(G197gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(KEYINPUT12), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n254), .A2(new_n261), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n246), .A2(new_n252), .A3(new_n253), .A4(new_n260), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT94), .ZN(new_n264));
  AND2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n263), .A2(new_n264), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n262), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(G228gat), .ZN(new_n269));
  INV_X1    g068(.A(G233gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT3), .ZN(new_n272));
  XNOR2_X1  g071(.A(G197gat), .B(G204gat), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT22), .ZN(new_n274));
  INV_X1    g073(.A(G211gat), .ZN(new_n275));
  INV_X1    g074(.A(G218gat), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G211gat), .B(G218gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n272), .B1(new_n280), .B2(KEYINPUT29), .ZN(new_n281));
  XNOR2_X1  g080(.A(G155gat), .B(G162gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(G155gat), .A2(G162gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT2), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT80), .ZN(new_n286));
  INV_X1    g085(.A(G141gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n286), .B1(new_n287), .B2(G148gat), .ZN(new_n288));
  INV_X1    g087(.A(G148gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n289), .A2(KEYINPUT80), .A3(G141gat), .ZN(new_n290));
  AND2_X1   g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n287), .A2(KEYINPUT79), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT79), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(G141gat), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n289), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT81), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n293), .A2(G141gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n287), .A2(KEYINPUT79), .ZN(new_n298));
  OAI21_X1  g097(.A(G148gat), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT81), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n288), .A2(new_n290), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n285), .B1(new_n296), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n282), .A2(KEYINPUT78), .ZN(new_n304));
  OR2_X1    g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT78), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(new_n306), .A3(new_n283), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G141gat), .B(G148gat), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n309), .B1(KEYINPUT2), .B2(new_n283), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n281), .B1(new_n303), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n302), .ZN(new_n313));
  INV_X1    g112(.A(new_n285), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n311), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT29), .B1(new_n315), .B2(new_n272), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n280), .B(KEYINPUT74), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n271), .B(new_n312), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT84), .ZN(new_n319));
  OR2_X1    g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n280), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n312), .B1(new_n316), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n322), .B1(new_n269), .B2(new_n270), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n318), .A2(new_n319), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n320), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT31), .B(G50gat), .ZN(new_n326));
  OR2_X1    g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  XOR2_X1   g126(.A(G78gat), .B(G106gat), .Z(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(G22gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n325), .A2(new_n326), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n327), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n329), .B1(new_n327), .B2(new_n330), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G120gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(G113gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT69), .B(G113gat), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n336), .B1(new_n337), .B2(G120gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT70), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT1), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  XOR2_X1   g139(.A(G127gat), .B(G134gat), .Z(new_n341));
  AND2_X1   g140(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n343));
  OAI21_X1  g142(.A(G120gat), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n335), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n341), .B1(new_n345), .B2(KEYINPUT70), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT68), .ZN(new_n347));
  INV_X1    g146(.A(G113gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G120gat), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n347), .B1(new_n335), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT1), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n335), .A2(new_n349), .A3(new_n347), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AOI22_X1  g153(.A1(new_n340), .A2(new_n346), .B1(new_n354), .B2(new_n341), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n315), .B(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G225gat), .A2(G233gat), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT83), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n353), .A2(new_n352), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n341), .B1(new_n361), .B2(new_n350), .ZN(new_n362));
  INV_X1    g161(.A(new_n341), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n363), .B1(new_n338), .B2(new_n339), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n352), .B1(new_n345), .B2(KEYINPUT70), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n362), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT4), .ZN(new_n367));
  NOR4_X1   g166(.A1(new_n366), .A2(new_n303), .A3(new_n367), .A4(new_n311), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT4), .B1(new_n315), .B2(new_n355), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n360), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n291), .A2(new_n295), .A3(KEYINPUT81), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n300), .B1(new_n299), .B2(new_n301), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n314), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n340), .A2(new_n346), .ZN(new_n374));
  INV_X1    g173(.A(new_n311), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n373), .A2(new_n374), .A3(new_n375), .A4(new_n362), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n367), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n315), .A2(KEYINPUT4), .A3(new_n355), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(KEYINPUT83), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n370), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT3), .B1(new_n303), .B2(new_n311), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n373), .A2(new_n272), .A3(new_n375), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n381), .A2(new_n382), .A3(new_n366), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n359), .B1(new_n384), .B2(new_n358), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT39), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT39), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n384), .A2(new_n387), .A3(new_n358), .ZN(new_n388));
  XNOR2_X1  g187(.A(KEYINPUT0), .B(G57gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n389), .B(G85gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(G1gat), .B(G29gat), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n390), .B(new_n391), .Z(new_n392));
  NAND4_X1  g191(.A1(new_n386), .A2(new_n388), .A3(KEYINPUT40), .A4(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n368), .A2(new_n369), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT82), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n394), .A2(new_n395), .A3(new_n357), .A4(new_n383), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n383), .A2(new_n377), .A3(new_n357), .A4(new_n378), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT82), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT5), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n399), .B1(new_n356), .B2(new_n358), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n396), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n380), .A2(new_n399), .A3(new_n357), .A4(new_n383), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n392), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n393), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n317), .ZN(new_n407));
  NAND2_X1  g206(.A1(G226gat), .A2(G233gat), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT66), .ZN(new_n410));
  NAND2_X1  g209(.A1(G183gat), .A2(G190gat), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n411), .A2(KEYINPUT24), .ZN(new_n412));
  AND2_X1   g211(.A1(G183gat), .A2(G190gat), .ZN(new_n413));
  NOR2_X1   g212(.A1(G183gat), .A2(G190gat), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n412), .B1(new_n415), .B2(KEYINPUT24), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT25), .B1(new_n416), .B2(KEYINPUT65), .ZN(new_n417));
  INV_X1    g216(.A(G183gat), .ZN(new_n418));
  INV_X1    g217(.A(G190gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n420), .A2(KEYINPUT24), .A3(new_n411), .ZN(new_n421));
  OR2_X1    g220(.A1(new_n411), .A2(KEYINPUT24), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(KEYINPUT65), .A3(new_n422), .ZN(new_n423));
  OR3_X1    g222(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n424), .A2(new_n425), .B1(G169gat), .B2(G176gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n410), .B1(new_n417), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT25), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n421), .A2(new_n422), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT65), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n432), .A2(KEYINPUT66), .A3(new_n423), .A4(new_n426), .ZN(new_n433));
  INV_X1    g232(.A(new_n425), .ZN(new_n434));
  NOR3_X1   g233(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n435));
  INV_X1    g234(.A(G169gat), .ZN(new_n436));
  INV_X1    g235(.A(G176gat), .ZN(new_n437));
  OAI22_X1  g236(.A1(new_n434), .A2(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n429), .B1(new_n430), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT64), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT64), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n441), .B(new_n429), .C1(new_n430), .C2(new_n438), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n428), .A2(new_n433), .A3(new_n440), .A4(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT27), .B(G183gat), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n419), .ZN(new_n445));
  NOR2_X1   g244(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  OR3_X1    g246(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n448), .B(new_n449), .C1(new_n436), .C2(new_n437), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n447), .A2(new_n411), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n443), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT75), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT75), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n443), .A2(new_n454), .A3(new_n451), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT29), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n409), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n408), .B1(new_n443), .B2(new_n451), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT76), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n459), .B(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n407), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT30), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n453), .A2(new_n409), .A3(new_n455), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n452), .A2(new_n457), .A3(new_n408), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n280), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(G64gat), .B(G92gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n468), .B(G36gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n469), .B(KEYINPUT77), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n470), .B(new_n202), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n462), .A2(new_n463), .A3(new_n467), .A4(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n471), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n443), .A2(new_n454), .A3(new_n451), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n454), .B1(new_n443), .B2(new_n451), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n457), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n408), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n459), .B(KEYINPUT76), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n317), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n473), .B1(new_n479), .B2(new_n466), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n462), .A2(new_n467), .A3(new_n471), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(new_n481), .A3(KEYINPUT30), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n386), .A2(new_n392), .A3(new_n388), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT40), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n406), .A2(new_n472), .A3(new_n482), .A4(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n401), .A2(new_n402), .A3(new_n392), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT6), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n392), .B1(new_n401), .B2(new_n402), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI211_X1 g290(.A(new_n488), .B(new_n392), .C1(new_n401), .C2(new_n402), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT38), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT37), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n495), .B1(new_n479), .B2(new_n466), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n462), .A2(KEYINPUT37), .A3(new_n467), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n471), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n493), .B(new_n481), .C1(new_n494), .C2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n477), .A2(new_n317), .A3(new_n478), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n464), .A2(new_n280), .A3(new_n465), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n500), .A2(KEYINPUT37), .A3(new_n501), .ZN(new_n502));
  AOI211_X1 g301(.A(KEYINPUT38), .B(new_n471), .C1(new_n496), .C2(new_n502), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n333), .B(new_n486), .C1(new_n499), .C2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT85), .ZN(new_n505));
  INV_X1    g304(.A(new_n492), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n405), .A2(new_n488), .A3(new_n487), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n482), .A2(new_n472), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n508), .A2(new_n333), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT71), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n510), .B1(new_n452), .B2(new_n366), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n452), .A2(new_n366), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n443), .A2(KEYINPUT71), .A3(new_n355), .A4(new_n451), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AND2_X1   g313(.A1(G227gat), .A2(G233gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT32), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT72), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G15gat), .B(G43gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(G71gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(G99gat), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT33), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n522), .B1(new_n516), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n516), .A2(KEYINPUT72), .A3(KEYINPUT32), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n519), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n516), .B(KEYINPUT32), .C1(new_n523), .C2(new_n522), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OR2_X1    g327(.A1(new_n514), .A2(new_n515), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT34), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n531), .A2(new_n526), .A3(new_n527), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT73), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT36), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g339(.A1(KEYINPUT73), .A2(KEYINPUT36), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n533), .B(new_n534), .C1(new_n538), .C2(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n509), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n498), .A2(new_n494), .ZN(new_n544));
  INV_X1    g343(.A(new_n503), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n544), .A2(new_n545), .A3(new_n493), .A4(new_n481), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT85), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n546), .A2(new_n547), .A3(new_n333), .A4(new_n486), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n505), .A2(new_n543), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT35), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT86), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT87), .B1(new_n508), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n533), .A2(new_n333), .A3(new_n534), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n550), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n533), .A2(new_n534), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n551), .B1(KEYINPUT87), .B2(KEYINPUT35), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n555), .A2(new_n508), .A3(new_n333), .A4(new_n557), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n268), .B1(new_n549), .B2(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(KEYINPUT101), .B(G204gat), .Z(new_n561));
  XNOR2_X1  g360(.A(G120gat), .B(G148gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(KEYINPUT100), .B(G176gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G99gat), .A2(G106gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT98), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT98), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n569), .A2(G99gat), .A3(G106gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n568), .A2(new_n570), .A3(KEYINPUT8), .ZN(new_n571));
  INV_X1    g370(.A(G92gat), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n572), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n573));
  OAI21_X1  g372(.A(G92gat), .B1(KEYINPUT7), .B2(G85gat), .ZN(new_n574));
  AND2_X1   g373(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G99gat), .B(G106gat), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G71gat), .A2(G78gat), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(G71gat), .A2(G78gat), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G57gat), .B(G64gat), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT9), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n581), .A2(new_n586), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT95), .ZN(new_n589));
  INV_X1    g388(.A(G64gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(G57gat), .ZN(new_n591));
  INV_X1    g390(.A(G57gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(G64gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G71gat), .B(G78gat), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT95), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n581), .A2(new_n596), .A3(new_n586), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n589), .A2(new_n594), .A3(new_n595), .A4(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n571), .A2(new_n576), .A3(new_n578), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n580), .A2(new_n587), .A3(new_n598), .A4(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n587), .ZN(new_n601));
  AND3_X1   g400(.A1(new_n571), .A2(new_n576), .A3(new_n578), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n578), .B1(new_n571), .B2(new_n576), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT10), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n600), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n602), .A2(new_n603), .ZN(new_n607));
  INV_X1    g406(.A(new_n601), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n607), .A2(new_n608), .A3(KEYINPUT10), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G230gat), .A2(G233gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT102), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT102), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n610), .A2(new_n614), .A3(new_n611), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n604), .ZN(new_n617));
  INV_X1    g416(.A(new_n611), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n566), .B1(new_n616), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT103), .ZN(new_n622));
  AND3_X1   g421(.A1(new_n606), .A2(KEYINPUT99), .A3(new_n609), .ZN(new_n623));
  AOI21_X1  g422(.A(KEYINPUT99), .B1(new_n606), .B2(new_n609), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n611), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n625), .A2(new_n619), .A3(new_n565), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n621), .A2(new_n622), .A3(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n622), .B1(new_n621), .B2(new_n626), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n560), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n242), .B1(KEYINPUT21), .B2(new_n608), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G183gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(G231gat), .A2(G233gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(G127gat), .B(G155gat), .Z(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT20), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n636), .B(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n608), .A2(KEYINPUT21), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(G211gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n640), .B(new_n642), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n639), .A2(new_n643), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  OAI221_X1 g446(.A(new_n234), .B1(new_n602), .B2(new_n603), .C1(new_n238), .C2(new_n239), .ZN(new_n648));
  AND2_X1   g447(.A1(G232gat), .A2(G233gat), .ZN(new_n649));
  AOI22_X1  g448(.A1(new_n236), .A2(new_n607), .B1(KEYINPUT41), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G134gat), .B(G162gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(G190gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n651), .B(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n649), .A2(KEYINPUT41), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT97), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G218gat), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n654), .A2(new_n657), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n647), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n632), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n493), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(new_n203), .ZN(G1324gat));
  NAND2_X1  g466(.A1(new_n482), .A2(new_n472), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n632), .A2(new_n663), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT16), .B(G8gat), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT104), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n672), .A2(KEYINPUT42), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n670), .A2(G8gat), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(KEYINPUT42), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(G1325gat));
  INV_X1    g475(.A(G15gat), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n540), .A2(new_n542), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n664), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n632), .A2(new_n663), .A3(new_n555), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n679), .B1(new_n677), .B2(new_n680), .ZN(G1326gat));
  NOR2_X1   g480(.A1(new_n664), .A2(new_n333), .ZN(new_n682));
  XOR2_X1   g481(.A(KEYINPUT43), .B(G22gat), .Z(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(G1327gat));
  NOR2_X1   g483(.A1(new_n647), .A2(new_n630), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(new_n660), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(KEYINPUT105), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n686), .A2(KEYINPUT105), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n560), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n690), .A2(new_n220), .A3(new_n493), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n692));
  OR2_X1    g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT107), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n554), .A2(new_n694), .A3(new_n558), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n694), .B1(new_n554), .B2(new_n558), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n549), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n660), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n549), .A2(new_n559), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n701), .A2(KEYINPUT44), .A3(new_n660), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n700), .A2(new_n267), .A3(new_n685), .A4(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(G29gat), .B1(new_n703), .B2(new_n665), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n691), .A2(new_n692), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n693), .A2(new_n704), .A3(new_n705), .ZN(G1328gat));
  NAND3_X1  g505(.A1(new_n690), .A2(new_n221), .A3(new_n669), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n707), .A2(KEYINPUT46), .ZN(new_n708));
  OAI21_X1  g507(.A(G36gat), .B1(new_n703), .B2(new_n668), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(KEYINPUT46), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(G1329gat));
  NOR3_X1   g510(.A1(new_n689), .A2(G43gat), .A3(new_n535), .ZN(new_n712));
  AOI21_X1  g511(.A(KEYINPUT44), .B1(new_n697), .B2(new_n660), .ZN(new_n713));
  AOI211_X1 g512(.A(new_n699), .B(new_n661), .C1(new_n549), .C2(new_n559), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n678), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n715), .A2(new_n267), .A3(new_n716), .A4(new_n685), .ZN(new_n717));
  AOI211_X1 g516(.A(KEYINPUT47), .B(new_n712), .C1(new_n717), .C2(G43gat), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT47), .ZN(new_n719));
  OAI21_X1  g518(.A(G43gat), .B1(new_n703), .B2(new_n678), .ZN(new_n720));
  INV_X1    g519(.A(new_n712), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n719), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n718), .A2(new_n722), .ZN(G1330gat));
  NOR3_X1   g522(.A1(new_n689), .A2(G50gat), .A3(new_n333), .ZN(new_n724));
  INV_X1    g523(.A(new_n333), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n715), .A2(new_n267), .A3(new_n725), .A4(new_n685), .ZN(new_n726));
  AOI211_X1 g525(.A(KEYINPUT48), .B(new_n724), .C1(new_n726), .C2(G50gat), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT48), .ZN(new_n728));
  OAI21_X1  g527(.A(G50gat), .B1(new_n703), .B2(new_n333), .ZN(new_n729));
  INV_X1    g528(.A(new_n724), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n727), .A2(new_n731), .ZN(G1331gat));
  NAND3_X1  g531(.A1(new_n647), .A2(new_n661), .A3(new_n268), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n733), .A2(new_n631), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n734), .B(KEYINPUT108), .Z(new_n735));
  NAND2_X1  g534(.A1(new_n697), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n736), .A2(new_n665), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(new_n592), .ZN(G1332gat));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(KEYINPUT109), .B1(new_n697), .B2(new_n735), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n668), .B(KEYINPUT110), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n746));
  AND2_X1   g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n745), .B2(new_n746), .ZN(G1333gat));
  NOR3_X1   g548(.A1(new_n736), .A2(G71gat), .A3(new_n535), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n716), .B1(new_n740), .B2(new_n741), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n750), .B1(new_n751), .B2(G71gat), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g552(.A1(new_n742), .A2(new_n333), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n754), .B(G78gat), .Z(G1335gat));
  NAND2_X1  g554(.A1(new_n646), .A2(new_n268), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT111), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n700), .A2(new_n630), .A3(new_n702), .A4(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(G85gat), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n759), .A2(new_n760), .A3(new_n665), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n697), .A2(new_n660), .A3(new_n758), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n697), .A2(KEYINPUT51), .A3(new_n660), .A4(new_n758), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n762), .A2(KEYINPUT112), .A3(new_n763), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n767), .A2(new_n493), .A3(new_n630), .A4(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n761), .B1(new_n760), .B2(new_n769), .ZN(G1336gat));
  NOR4_X1   g569(.A1(new_n713), .A2(new_n714), .A3(new_n631), .A4(new_n757), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n572), .B1(new_n771), .B2(new_n669), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n744), .A2(G92gat), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  AOI211_X1 g573(.A(new_n631), .B(new_n774), .C1(new_n764), .C2(new_n766), .ZN(new_n775));
  OAI21_X1  g574(.A(KEYINPUT52), .B1(new_n772), .B2(new_n775), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n767), .A2(new_n630), .A3(new_n768), .A4(new_n773), .ZN(new_n777));
  OAI21_X1  g576(.A(G92gat), .B1(new_n759), .B2(new_n744), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n776), .A2(new_n780), .ZN(G1337gat));
  OAI21_X1  g580(.A(G99gat), .B1(new_n759), .B2(new_n678), .ZN(new_n782));
  INV_X1    g581(.A(G99gat), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n767), .A2(new_n783), .A3(new_n630), .A4(new_n768), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n782), .B1(new_n784), .B2(new_n535), .ZN(G1338gat));
  INV_X1    g584(.A(G106gat), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n786), .B1(new_n771), .B2(new_n725), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n333), .A2(G106gat), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  AOI211_X1 g588(.A(new_n631), .B(new_n789), .C1(new_n764), .C2(new_n766), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT53), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n767), .A2(new_n630), .A3(new_n768), .A4(new_n788), .ZN(new_n792));
  OAI21_X1  g591(.A(G106gat), .B1(new_n759), .B2(new_n333), .ZN(new_n793));
  XNOR2_X1  g592(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n791), .A2(new_n795), .ZN(G1339gat));
  INV_X1    g595(.A(KEYINPUT117), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n733), .A2(new_n630), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n565), .B1(new_n616), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n606), .A2(new_n618), .A3(new_n609), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n802), .A2(KEYINPUT54), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n801), .B1(new_n625), .B2(new_n803), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n625), .A2(new_n801), .A3(new_n803), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n800), .B(KEYINPUT55), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n626), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT115), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT115), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n806), .A2(new_n809), .A3(new_n626), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n800), .B1(new_n805), .B2(new_n804), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n808), .A2(new_n267), .A3(new_n810), .A4(new_n813), .ZN(new_n814));
  OR2_X1    g613(.A1(new_n265), .A2(new_n266), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n240), .A2(new_n243), .ZN(new_n816));
  OAI22_X1  g615(.A1(new_n816), .A2(new_n241), .B1(new_n251), .B2(new_n249), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n259), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n815), .A2(new_n630), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n814), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT116), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n814), .A2(new_n822), .A3(new_n819), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(new_n661), .A3(new_n823), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n815), .A2(new_n818), .ZN(new_n825));
  INV_X1    g624(.A(new_n813), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n826), .B1(KEYINPUT115), .B2(new_n807), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n825), .A2(new_n660), .A3(new_n827), .A4(new_n810), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n824), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n798), .B1(new_n829), .B2(new_n646), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n797), .B1(new_n830), .B2(new_n725), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n647), .B1(new_n824), .B2(new_n828), .ZN(new_n832));
  OAI211_X1 g631(.A(KEYINPUT117), .B(new_n333), .C1(new_n832), .C2(new_n798), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n743), .A2(new_n665), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n555), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(G113gat), .B1(new_n836), .B2(new_n268), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n830), .A2(new_n665), .ZN(new_n838));
  INV_X1    g637(.A(new_n553), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n744), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n267), .A2(new_n337), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n837), .B1(new_n842), .B2(new_n843), .ZN(G1340gat));
  OAI21_X1  g643(.A(G120gat), .B1(new_n836), .B2(new_n631), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n841), .A2(new_n334), .A3(new_n744), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n845), .B1(new_n631), .B2(new_n846), .ZN(G1341gat));
  INV_X1    g646(.A(G127gat), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n836), .A2(new_n848), .A3(new_n646), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT118), .B1(new_n842), .B2(new_n646), .ZN(new_n850));
  OR4_X1    g649(.A1(KEYINPUT118), .A2(new_n840), .A3(new_n646), .A4(new_n743), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n849), .B1(new_n852), .B2(new_n848), .ZN(G1342gat));
  NOR4_X1   g652(.A1(new_n840), .A2(G134gat), .A3(new_n661), .A4(new_n669), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT56), .ZN(new_n855));
  OAI21_X1  g654(.A(G134gat), .B1(new_n836), .B2(new_n661), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1343gat));
  NAND2_X1  g656(.A1(new_n829), .A2(new_n646), .ZN(new_n858));
  INV_X1    g657(.A(new_n798), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n861), .A3(new_n725), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n835), .A2(new_n678), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n268), .A2(new_n807), .A3(new_n826), .ZN(new_n864));
  INV_X1    g663(.A(new_n819), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n661), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n647), .B1(new_n866), .B2(new_n828), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n725), .B1(new_n867), .B2(new_n798), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n863), .B1(new_n868), .B2(KEYINPUT57), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n862), .A2(new_n869), .A3(new_n267), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n297), .A2(new_n298), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT58), .B1(new_n872), .B2(KEYINPUT119), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n678), .A2(new_n725), .ZN(new_n874));
  NOR4_X1   g673(.A1(new_n830), .A2(new_n665), .A3(new_n743), .A4(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n268), .A2(G141gat), .ZN(new_n876));
  AOI22_X1  g675(.A1(new_n870), .A2(new_n871), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n873), .B(new_n877), .ZN(G1344gat));
  NAND3_X1  g677(.A1(new_n875), .A2(new_n289), .A3(new_n630), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT120), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n860), .A2(KEYINPUT57), .A3(new_n725), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n868), .A2(new_n861), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n630), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n885), .A2(new_n863), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n881), .B1(new_n886), .B2(G148gat), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n862), .A2(new_n869), .ZN(new_n888));
  AOI211_X1 g687(.A(KEYINPUT59), .B(new_n289), .C1(new_n888), .C2(new_n630), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n880), .B1(new_n887), .B2(new_n889), .ZN(G1345gat));
  AOI21_X1  g689(.A(G155gat), .B1(new_n875), .B2(new_n647), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n647), .A2(G155gat), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT121), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n891), .B1(new_n888), .B2(new_n893), .ZN(G1346gat));
  NOR3_X1   g693(.A1(new_n669), .A2(new_n661), .A3(G162gat), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n838), .A2(new_n725), .A3(new_n678), .A4(new_n895), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n888), .A2(new_n660), .ZN(new_n897));
  INV_X1    g696(.A(G162gat), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(G1347gat));
  NAND2_X1  g698(.A1(new_n669), .A2(new_n665), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n900), .A2(new_n535), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n902), .B1(new_n831), .B2(new_n833), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n436), .B1(new_n903), .B2(new_n267), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n743), .A2(new_n665), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n860), .A2(new_n839), .A3(new_n906), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n907), .A2(G169gat), .A3(new_n268), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n904), .A2(new_n908), .ZN(G1348gat));
  INV_X1    g708(.A(new_n907), .ZN(new_n910));
  AOI21_X1  g709(.A(G176gat), .B1(new_n910), .B2(new_n630), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n631), .A2(new_n437), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n911), .B1(new_n903), .B2(new_n912), .ZN(G1349gat));
  INV_X1    g712(.A(KEYINPUT122), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n647), .A2(new_n444), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n914), .B1(new_n907), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n903), .A2(new_n647), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n917), .B2(G183gat), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT60), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n918), .B(new_n919), .ZN(G1350gat));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n921));
  AOI211_X1 g720(.A(new_n661), .B(new_n902), .C1(new_n831), .C2(new_n833), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n921), .B1(new_n922), .B2(new_n419), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n834), .A2(new_n660), .A3(new_n901), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n924), .A2(KEYINPUT61), .A3(G190gat), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT123), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n910), .A2(new_n926), .A3(new_n419), .A4(new_n660), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n830), .A2(new_n905), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n928), .A2(new_n419), .A3(new_n660), .A4(new_n839), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(KEYINPUT123), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n923), .A2(new_n925), .A3(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n923), .A2(new_n925), .A3(new_n931), .A4(KEYINPUT124), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1351gat));
  NAND3_X1  g735(.A1(new_n928), .A2(new_n725), .A3(new_n678), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(G197gat), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n938), .A2(new_n939), .A3(new_n267), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n716), .A2(new_n900), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n945), .B1(new_n882), .B2(new_n883), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n946), .A2(new_n267), .ZN(new_n947));
  OAI22_X1  g746(.A1(new_n942), .A2(new_n943), .B1(new_n939), .B2(new_n947), .ZN(G1352gat));
  NOR3_X1   g747(.A1(new_n937), .A2(G204gat), .A3(new_n631), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT62), .ZN(new_n950));
  OR2_X1    g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g750(.A(G204gat), .B1(new_n885), .B2(new_n945), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n949), .A2(new_n950), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(G1353gat));
  NAND3_X1  g753(.A1(new_n938), .A2(new_n275), .A3(new_n647), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n946), .A2(new_n647), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n956), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT63), .B1(new_n956), .B2(G211gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(G1354gat));
  AOI21_X1  g758(.A(G218gat), .B1(new_n938), .B2(new_n660), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n660), .A2(G218gat), .ZN(new_n961));
  XOR2_X1   g760(.A(new_n961), .B(KEYINPUT126), .Z(new_n962));
  AOI21_X1  g761(.A(new_n960), .B1(new_n946), .B2(new_n962), .ZN(G1355gat));
endmodule


