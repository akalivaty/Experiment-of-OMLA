//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 0 1 0 0 1 1 1 0 1 1 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n562, new_n563, new_n565,
    new_n566, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n585, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n629, new_n632,
    new_n634, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1271, new_n1272, new_n1273;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  NAND2_X1  g032(.A1(G113), .A2(G2104), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT64), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n458), .B(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  AND3_X1   g039(.A1(new_n462), .A2(new_n464), .A3(G125), .ZN(new_n465));
  OAI21_X1  g040(.A(G2105), .B1(new_n460), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n461), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n462), .B1(new_n470), .B2(KEYINPUT65), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT65), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(new_n461), .A3(KEYINPUT3), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n471), .A2(G137), .A3(new_n472), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT67), .ZN(new_n480));
  AOI21_X1  g055(.A(KEYINPUT65), .B1(new_n463), .B2(G2104), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n463), .A2(G2104), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n472), .B(new_n474), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n484), .A2(KEYINPUT66), .A3(G136), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT66), .ZN(new_n486));
  INV_X1    g061(.A(G136), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n486), .B1(new_n483), .B2(new_n487), .ZN(new_n488));
  OAI211_X1 g063(.A(G2105), .B(new_n474), .C1(new_n481), .C2(new_n482), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n480), .A2(new_n485), .A3(new_n488), .A4(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT4), .B1(new_n483), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n482), .A2(new_n470), .ZN(new_n496));
  NOR3_X1   g071(.A1(new_n494), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G126), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n472), .A2(G114), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  OAI22_X1  g077(.A1(new_n489), .A2(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  XNOR2_X1  g081(.A(KEYINPUT5), .B(G543), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n509), .A2(KEYINPUT6), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G651), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n515), .A2(new_n517), .A3(new_n518), .A4(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n512), .A2(new_n513), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n510), .A2(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  INV_X1    g100(.A(G51), .ZN(new_n526));
  INV_X1    g101(.A(G89), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n512), .A2(new_n526), .B1(new_n521), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT7), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n530), .A2(new_n531), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n529), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n528), .A2(new_n534), .ZN(G168));
  AOI22_X1  g110(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n509), .ZN(new_n537));
  INV_X1    g112(.A(G52), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n512), .A2(new_n538), .B1(new_n521), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n537), .A2(new_n540), .ZN(G171));
  NAND2_X1  g116(.A1(new_n507), .A2(G56), .ZN(new_n542));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n509), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n507), .A2(new_n511), .A3(G81), .ZN(new_n546));
  NAND4_X1  g121(.A1(new_n518), .A2(new_n520), .A3(G43), .A4(G543), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n546), .A2(KEYINPUT68), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g123(.A(KEYINPUT68), .B1(new_n546), .B2(new_n547), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n545), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(KEYINPUT69), .ZN(new_n551));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n547), .B1(new_n521), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT68), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n546), .A2(KEYINPUT68), .A3(new_n547), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT69), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n557), .A2(new_n558), .A3(new_n545), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n551), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  AND3_X1   g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G36), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT70), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n562), .A2(new_n566), .ZN(G188));
  INV_X1    g142(.A(G91), .ZN(new_n568));
  OAI21_X1  g143(.A(KEYINPUT71), .B1(new_n521), .B2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT71), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n507), .A2(new_n511), .A3(new_n570), .A4(G91), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n511), .A2(G53), .A3(G543), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(KEYINPUT9), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n511), .A2(new_n575), .A3(G53), .A4(G543), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(G78), .A2(G543), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n515), .A2(new_n517), .ZN(new_n579));
  INV_X1    g154(.A(G65), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n572), .A2(new_n577), .A3(new_n582), .ZN(G299));
  INV_X1    g158(.A(G171), .ZN(G301));
  XNOR2_X1  g159(.A(G168), .B(KEYINPUT72), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G286));
  INV_X1    g161(.A(G74), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n509), .B1(new_n579), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n512), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n588), .B1(new_n589), .B2(G49), .ZN(new_n590));
  INV_X1    g165(.A(new_n521), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n591), .A2(KEYINPUT73), .A3(G87), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT73), .ZN(new_n593));
  INV_X1    g168(.A(G87), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n521), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n590), .A2(new_n592), .A3(new_n595), .ZN(G288));
  NAND3_X1  g171(.A1(new_n511), .A2(G48), .A3(G543), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT74), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n591), .A2(G86), .ZN(new_n599));
  NAND2_X1  g174(.A1(G73), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G61), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n579), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G651), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n598), .A2(new_n599), .A3(new_n603), .ZN(G305));
  AOI22_X1  g179(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n509), .B1(new_n605), .B2(KEYINPUT75), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(KEYINPUT75), .B2(new_n605), .ZN(new_n607));
  AOI22_X1  g182(.A1(G47), .A2(new_n589), .B1(new_n591), .B2(G85), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(G54), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT76), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n611), .B1(new_n512), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n511), .A2(KEYINPUT76), .A3(G543), .ZN(new_n614));
  NAND2_X1  g189(.A1(G79), .A2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G66), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n579), .B2(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n613), .A2(new_n614), .B1(G651), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n591), .A2(KEYINPUT10), .A3(G92), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT10), .ZN(new_n620));
  INV_X1    g195(.A(G92), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n521), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n610), .B1(new_n625), .B2(G868), .ZN(G284));
  OAI21_X1  g201(.A(new_n610), .B1(new_n625), .B2(G868), .ZN(G321));
  INV_X1    g202(.A(G868), .ZN(new_n628));
  NAND2_X1  g203(.A1(G299), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(new_n585), .B2(new_n628), .ZN(G297));
  OAI21_X1  g205(.A(new_n629), .B1(new_n585), .B2(new_n628), .ZN(G280));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n625), .B1(new_n632), .B2(G860), .ZN(G148));
  NOR2_X1   g208(.A1(new_n624), .A2(G559), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(G868), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(new_n560), .B2(G868), .ZN(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g213(.A1(new_n472), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT12), .Z(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(KEYINPUT13), .ZN(new_n642));
  AOI22_X1  g217(.A1(new_n641), .A2(new_n642), .B1(KEYINPUT77), .B2(G2100), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(new_n642), .B2(new_n641), .ZN(new_n644));
  NOR2_X1   g219(.A1(KEYINPUT77), .A2(G2100), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n490), .A2(G123), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n484), .A2(G135), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n472), .A2(G111), .ZN(new_n649));
  OAI21_X1  g224(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n647), .B(new_n648), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(G2096), .Z(new_n652));
  NAND2_X1  g227(.A1(new_n646), .A2(new_n652), .ZN(G156));
  INV_X1    g228(.A(G14), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2427), .B(G2430), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT80), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT79), .B(G2438), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT80), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n661), .B(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n663), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT15), .B(G2435), .Z(new_n669));
  NAND3_X1  g244(.A1(new_n664), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n670), .A2(KEYINPUT14), .ZN(new_n671));
  INV_X1    g246(.A(new_n669), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n666), .A2(new_n667), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n662), .A2(new_n663), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n660), .B1(new_n671), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n675), .A2(KEYINPUT14), .A3(new_n670), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n677), .A2(new_n659), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n658), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n671), .A2(new_n660), .A3(new_n675), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n659), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n680), .A2(new_n681), .A3(new_n657), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1341), .B(G1348), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT81), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n654), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT82), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n679), .A2(new_n682), .ZN(new_n688));
  INV_X1    g263(.A(new_n685), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  AOI211_X1 g265(.A(KEYINPUT82), .B(new_n685), .C1(new_n679), .C2(new_n682), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n686), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(G401));
  XOR2_X1   g268(.A(G2084), .B(G2090), .Z(new_n694));
  XNOR2_X1  g269(.A(G2067), .B(G2678), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G2072), .B(G2078), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n694), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n697), .B(KEYINPUT17), .Z(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(new_n696), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT83), .Z(new_n702));
  NAND3_X1  g277(.A1(new_n694), .A2(new_n695), .A3(new_n697), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT18), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n696), .A2(new_n694), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n704), .B1(new_n700), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(G2096), .B(G2100), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(G227));
  XNOR2_X1  g284(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G1996), .ZN(new_n712));
  XOR2_X1   g287(.A(G1956), .B(G2474), .Z(new_n713));
  XOR2_X1   g288(.A(G1961), .B(G1966), .Z(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(G1971), .B(G1976), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT19), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT84), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n713), .A2(new_n714), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT20), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(KEYINPUT20), .B1(new_n718), .B2(new_n721), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n716), .A2(new_n718), .A3(new_n721), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n720), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n728), .A2(G1991), .ZN(new_n729));
  INV_X1    g304(.A(G1991), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n726), .A2(new_n727), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(new_n720), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n712), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(G1981), .B(G1986), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n728), .A2(G1991), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n731), .A2(new_n730), .A3(new_n720), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n736), .A2(new_n737), .A3(G1996), .ZN(new_n738));
  AND3_X1   g313(.A1(new_n733), .A2(new_n735), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n735), .B1(new_n733), .B2(new_n738), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n711), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n733), .A2(new_n738), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(new_n734), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n733), .A2(new_n735), .A3(new_n738), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n743), .A2(new_n710), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n741), .A2(new_n745), .ZN(G229));
  NAND3_X1  g321(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT26), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n748), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n749), .A2(new_n750), .B1(G105), .B2(new_n467), .ZN(new_n751));
  INV_X1    g326(.A(G141), .ZN(new_n752));
  INV_X1    g327(.A(G129), .ZN(new_n753));
  OAI221_X1 g328(.A(new_n751), .B1(new_n483), .B2(new_n752), .C1(new_n753), .C2(new_n489), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G29), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G29), .B2(G32), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT27), .B(G1996), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT97), .Z(new_n760));
  NAND2_X1  g335(.A1(new_n467), .A2(G103), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT25), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n496), .A2(G127), .ZN(new_n763));
  INV_X1    g338(.A(G115), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(new_n461), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n762), .B1(new_n765), .B2(G2105), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n484), .A2(G139), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(G29), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G29), .B2(G33), .ZN(new_n770));
  INV_X1    g345(.A(G2072), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT95), .ZN(new_n773));
  NOR2_X1   g348(.A1(G27), .A2(G29), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G164), .B2(G29), .ZN(new_n775));
  AOI211_X1 g350(.A(new_n760), .B(new_n773), .C1(G2078), .C2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G29), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n777), .A2(G26), .ZN(new_n778));
  INV_X1    g353(.A(G128), .ZN(new_n779));
  OR3_X1    g354(.A1(new_n489), .A2(KEYINPUT94), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n484), .A2(G140), .ZN(new_n781));
  OAI21_X1  g356(.A(KEYINPUT94), .B1(new_n489), .B2(new_n779), .ZN(new_n782));
  OR2_X1    g357(.A1(G104), .A2(G2105), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n783), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n780), .A2(new_n781), .A3(new_n782), .A4(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n778), .B1(new_n786), .B2(new_n777), .ZN(new_n787));
  MUX2_X1   g362(.A(new_n778), .B(new_n787), .S(KEYINPUT28), .Z(new_n788));
  INV_X1    g363(.A(G2067), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(G5), .A2(G16), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G171), .B2(G16), .ZN(new_n792));
  INV_X1    g367(.A(G1961), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(G16), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(G21), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G168), .B2(new_n795), .ZN(new_n797));
  OAI221_X1 g372(.A(new_n794), .B1(new_n777), .B2(new_n651), .C1(G1966), .C2(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n625), .A2(new_n795), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G4), .B2(new_n795), .ZN(new_n800));
  INV_X1    g375(.A(G1348), .ZN(new_n801));
  OAI22_X1  g376(.A1(new_n800), .A2(new_n801), .B1(new_n757), .B2(new_n758), .ZN(new_n802));
  AOI211_X1 g377(.A(new_n798), .B(new_n802), .C1(new_n801), .C2(new_n800), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT24), .B(G34), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(new_n777), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT96), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n476), .B2(new_n777), .ZN(new_n807));
  INV_X1    g382(.A(G2084), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n770), .B2(new_n771), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n775), .A2(G2078), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n797), .A2(G1966), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT30), .B(G28), .ZN(new_n813));
  OR2_X1    g388(.A1(KEYINPUT31), .A2(G11), .ZN(new_n814));
  NAND2_X1  g389(.A1(KEYINPUT31), .A2(G11), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n813), .A2(new_n777), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n812), .B(new_n816), .C1(new_n807), .C2(new_n808), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n810), .A2(new_n811), .A3(new_n817), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n776), .A2(new_n790), .A3(new_n803), .A4(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(G16), .A2(G19), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(new_n560), .B2(G16), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT93), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G1341), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n777), .A2(G35), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(G162), .B2(new_n777), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT29), .Z(new_n826));
  INV_X1    g401(.A(G2090), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(G299), .ZN(new_n829));
  OAI21_X1  g404(.A(KEYINPUT23), .B1(new_n829), .B2(new_n795), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n795), .A2(G20), .ZN(new_n831));
  MUX2_X1   g406(.A(KEYINPUT23), .B(new_n830), .S(new_n831), .Z(new_n832));
  INV_X1    g407(.A(G1956), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n826), .A2(new_n827), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n828), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  OR3_X1    g411(.A1(new_n819), .A2(new_n823), .A3(new_n836), .ZN(new_n837));
  OR2_X1    g412(.A1(G95), .A2(G2105), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n838), .B(G2104), .C1(G107), .C2(new_n472), .ZN(new_n839));
  INV_X1    g414(.A(G131), .ZN(new_n840));
  INV_X1    g415(.A(G119), .ZN(new_n841));
  OAI221_X1 g416(.A(new_n839), .B1(new_n483), .B2(new_n840), .C1(new_n841), .C2(new_n489), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT85), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n843), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT86), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(G29), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(G25), .B2(G29), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT87), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(KEYINPUT35), .B(G1991), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n850), .B(KEYINPUT87), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(new_n853), .ZN(new_n857));
  NOR2_X1   g432(.A1(G16), .A2(G22), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n858), .B1(G166), .B2(G16), .ZN(new_n859));
  XOR2_X1   g434(.A(KEYINPUT91), .B(G1971), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n795), .A2(G6), .ZN(new_n862));
  INV_X1    g437(.A(G305), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n862), .B1(new_n863), .B2(new_n795), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(KEYINPUT32), .B(G1981), .Z(new_n866));
  AOI21_X1  g441(.A(new_n861), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(G288), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n868), .A2(new_n795), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n869), .B1(new_n795), .B2(G23), .ZN(new_n870));
  XNOR2_X1  g445(.A(KEYINPUT33), .B(G1976), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT90), .ZN(new_n872));
  INV_X1    g447(.A(new_n866), .ZN(new_n873));
  AOI22_X1  g448(.A1(new_n870), .A2(new_n872), .B1(new_n864), .B2(new_n873), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n867), .B(new_n874), .C1(new_n872), .C2(new_n870), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n875), .A2(KEYINPUT34), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT88), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n795), .A2(G24), .ZN(new_n878));
  AOI211_X1 g453(.A(new_n877), .B(new_n878), .C1(G290), .C2(G16), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n879), .B1(new_n877), .B2(new_n878), .ZN(new_n880));
  XNOR2_X1  g455(.A(KEYINPUT89), .B(G1986), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n880), .B(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n882), .B1(new_n875), .B2(KEYINPUT34), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n855), .A2(new_n857), .A3(new_n876), .A4(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT92), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(KEYINPUT36), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n884), .A2(new_n887), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n837), .B1(new_n888), .B2(new_n889), .ZN(G311));
  XNOR2_X1  g465(.A(new_n884), .B(new_n887), .ZN(new_n891));
  INV_X1    g466(.A(new_n837), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(G150));
  NAND2_X1  g468(.A1(new_n589), .A2(G55), .ZN(new_n894));
  NAND2_X1  g469(.A1(G80), .A2(G543), .ZN(new_n895));
  INV_X1    g470(.A(G67), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n895), .B1(new_n579), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(G651), .ZN(new_n898));
  XOR2_X1   g473(.A(KEYINPUT98), .B(G93), .Z(new_n899));
  OR2_X1    g474(.A1(new_n521), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n894), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n902), .B1(new_n551), .B2(new_n559), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT100), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n901), .A2(KEYINPUT99), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT99), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n894), .A2(new_n898), .A3(new_n900), .A4(new_n906), .ZN(new_n907));
  AOI22_X1  g482(.A1(new_n905), .A2(new_n907), .B1(new_n557), .B2(new_n545), .ZN(new_n908));
  NOR3_X1   g483(.A1(new_n903), .A2(new_n904), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n558), .B1(new_n557), .B2(new_n545), .ZN(new_n910));
  AOI211_X1 g485(.A(KEYINPUT69), .B(new_n544), .C1(new_n555), .C2(new_n556), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n901), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n905), .A2(new_n907), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n550), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT100), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n909), .A2(new_n915), .ZN(new_n916));
  XOR2_X1   g491(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n917));
  XNOR2_X1  g492(.A(new_n916), .B(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n624), .A2(new_n632), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(KEYINPUT39), .ZN(new_n921));
  AOI21_X1  g496(.A(G860), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n922), .B1(new_n921), .B2(new_n919), .ZN(new_n923));
  INV_X1    g498(.A(new_n913), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(G860), .ZN(new_n925));
  XOR2_X1   g500(.A(new_n925), .B(KEYINPUT37), .Z(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n926), .ZN(G145));
  OR2_X1    g502(.A1(G106), .A2(G2105), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n928), .B(G2104), .C1(G118), .C2(new_n472), .ZN(new_n929));
  INV_X1    g504(.A(G142), .ZN(new_n930));
  INV_X1    g505(.A(G130), .ZN(new_n931));
  OAI221_X1 g506(.A(new_n929), .B1(new_n483), .B2(new_n930), .C1(new_n931), .C2(new_n489), .ZN(new_n932));
  OR2_X1    g507(.A1(new_n932), .A2(new_n640), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n640), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OR2_X1    g510(.A1(new_n846), .A2(new_n935), .ZN(new_n936));
  AOI22_X1  g511(.A1(new_n845), .A2(new_n844), .B1(new_n933), .B2(new_n934), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n936), .A2(new_n938), .A3(KEYINPUT103), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT103), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n935), .A2(new_n846), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n940), .B1(new_n941), .B2(new_n937), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n768), .A2(G164), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n766), .A2(new_n767), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n505), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n944), .A2(new_n785), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n785), .B1(new_n944), .B2(new_n946), .ZN(new_n949));
  XOR2_X1   g524(.A(new_n754), .B(KEYINPUT102), .Z(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n948), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n944), .A2(new_n946), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n786), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n950), .B1(new_n954), .B2(new_n947), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n943), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n951), .B1(new_n948), .B2(new_n949), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n954), .A2(new_n950), .A3(new_n947), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n957), .A2(new_n958), .A3(new_n936), .A4(new_n938), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n476), .B(new_n651), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(G162), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n956), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n957), .A2(new_n958), .A3(new_n939), .A4(new_n942), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n961), .B1(new_n956), .B2(new_n963), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n962), .A2(new_n964), .A3(G37), .ZN(new_n965));
  XOR2_X1   g540(.A(new_n965), .B(KEYINPUT40), .Z(G395));
  OAI21_X1  g541(.A(new_n634), .B1(new_n909), .B2(new_n915), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT105), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT104), .ZN(new_n969));
  NAND2_X1  g544(.A1(G299), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n572), .A2(new_n577), .A3(KEYINPUT104), .A4(new_n582), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n625), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT41), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n624), .A2(new_n969), .A3(G299), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n973), .B1(new_n972), .B2(new_n974), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n968), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n904), .B1(new_n903), .B2(new_n908), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n912), .A2(KEYINPUT100), .A3(new_n914), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(new_n979), .A3(new_n635), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n972), .A2(new_n974), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT41), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT105), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n967), .A2(new_n977), .A3(new_n980), .A4(new_n983), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n978), .A2(new_n979), .A3(new_n635), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n635), .B1(new_n978), .B2(new_n979), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n981), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n988), .B(KEYINPUT42), .ZN(new_n989));
  XNOR2_X1  g564(.A(G290), .B(G305), .ZN(new_n990));
  XOR2_X1   g565(.A(G303), .B(G288), .Z(new_n991));
  XNOR2_X1  g566(.A(new_n990), .B(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n988), .A2(KEYINPUT42), .ZN(new_n994));
  INV_X1    g569(.A(new_n992), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n988), .A2(KEYINPUT42), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n993), .A2(G868), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT106), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n628), .B1(new_n989), .B2(new_n992), .ZN(new_n1001));
  AOI22_X1  g576(.A1(new_n1001), .A2(new_n997), .B1(new_n628), .B2(new_n924), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1000), .B1(new_n1002), .B2(new_n999), .ZN(G295));
  OAI21_X1  g578(.A(new_n1000), .B1(new_n1002), .B2(new_n999), .ZN(G331));
  INV_X1    g579(.A(G168), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1005), .A2(G171), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(new_n585), .B2(G301), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n978), .A2(new_n979), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1008), .B1(new_n978), .B2(new_n979), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n975), .A2(new_n976), .ZN(new_n1011));
  NOR3_X1   g586(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1008), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(new_n909), .B2(new_n915), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n978), .A2(new_n979), .A3(new_n1008), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n981), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g591(.A(KEYINPUT107), .B(new_n992), .C1(new_n1012), .C2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G37), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT105), .B1(new_n982), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n976), .A2(new_n968), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1015), .B(new_n1014), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n981), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1022), .A2(new_n995), .A3(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1017), .A2(new_n1018), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT43), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n982), .A2(new_n1019), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1014), .A2(new_n1028), .A3(new_n1015), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1024), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT107), .B1(new_n1030), .B2(new_n992), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n1026), .A2(new_n1027), .A3(new_n1031), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1025), .A2(new_n1018), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n992), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT43), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT44), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n1026), .A2(KEYINPUT43), .A3(new_n1031), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1027), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1037), .B1(new_n1040), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g616(.A(KEYINPUT113), .ZN(new_n1042));
  INV_X1    g617(.A(G1384), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n471), .A2(G138), .A3(new_n472), .A4(new_n474), .ZN(new_n1044));
  AOI22_X1  g619(.A1(new_n1044), .A2(KEYINPUT4), .B1(new_n496), .B2(new_n497), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1043), .B1(new_n1045), .B2(new_n503), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT45), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n466), .A2(G40), .A3(new_n475), .A4(new_n468), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1046), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT108), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT108), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1046), .A2(new_n1049), .A3(new_n1052), .A4(new_n1047), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1054), .A2(new_n712), .A3(new_n755), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT111), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1051), .A2(KEYINPUT110), .A3(new_n1053), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT110), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n754), .A2(G1996), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1056), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  NOR4_X1   g637(.A1(new_n1057), .A2(new_n1058), .A3(KEYINPUT111), .A4(new_n1060), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1055), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n786), .A2(new_n789), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n785), .A2(G2067), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT112), .B1(new_n1059), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT112), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1067), .ZN(new_n1070));
  NOR4_X1   g645(.A1(new_n1057), .A2(new_n1058), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1042), .B1(new_n1064), .B2(new_n1072), .ZN(new_n1073));
  OR2_X1    g648(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1074));
  OR2_X1    g649(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT111), .B1(new_n1075), .B2(new_n1060), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1063), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1074), .A2(new_n1078), .A3(KEYINPUT113), .A4(new_n1055), .ZN(new_n1079));
  XNOR2_X1  g654(.A(new_n846), .B(new_n853), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1059), .A2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(G290), .A2(G1986), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n1082), .B(KEYINPUT109), .ZN(new_n1083));
  AND2_X1   g658(.A1(G290), .A2(G1986), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1054), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AND4_X1   g660(.A1(new_n1073), .A2(new_n1079), .A3(new_n1081), .A4(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT125), .ZN(new_n1087));
  NAND2_X1  g662(.A1(G303), .A2(G8), .ZN(new_n1088));
  XNOR2_X1  g663(.A(new_n1088), .B(KEYINPUT55), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT114), .B(G1971), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1048), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n1043), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1091), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1046), .A2(KEYINPUT50), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT50), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n505), .A2(new_n1096), .A3(new_n1043), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1095), .A2(new_n1049), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(G2090), .B1(new_n1098), .B2(KEYINPUT118), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1048), .B1(new_n1046), .B2(KEYINPUT50), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1100), .A2(new_n1101), .A3(new_n1097), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1094), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1103));
  OR2_X1    g678(.A1(new_n1103), .A2(KEYINPUT119), .ZN(new_n1104));
  INV_X1    g679(.A(G8), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1105), .B1(new_n1103), .B2(KEYINPUT119), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1090), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1049), .A2(new_n505), .A3(new_n1043), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(G8), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT74), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n597), .B(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n603), .A2(new_n599), .ZN(new_n1112));
  OAI21_X1  g687(.A(G1981), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(G1981), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n598), .A2(new_n1114), .A3(new_n599), .A4(new_n603), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT49), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT116), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT116), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1116), .A2(new_n1120), .A3(new_n1117), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1109), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1113), .A2(new_n1115), .A3(KEYINPUT49), .ZN(new_n1123));
  XOR2_X1   g698(.A(new_n1123), .B(KEYINPUT117), .Z(new_n1124));
  NAND2_X1  g699(.A1(new_n868), .A2(G1976), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1125), .A2(new_n1108), .A3(G8), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT52), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n868), .B2(G1976), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT115), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1122), .A2(new_n1124), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1098), .A2(G2090), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1090), .B(G8), .C1(new_n1133), .C2(new_n1094), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1126), .A2(KEYINPUT52), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT115), .B1(new_n1135), .B2(new_n1129), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1132), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1087), .B1(new_n1107), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1094), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1139), .A2(KEYINPUT119), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(G8), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1103), .A2(KEYINPUT119), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1089), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1132), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1144), .A2(KEYINPUT125), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1138), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT53), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1149));
  INV_X1    g724(.A(G2078), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1149), .A2(new_n1150), .A3(new_n1093), .A4(new_n1049), .ZN(new_n1151));
  AOI22_X1  g726(.A1(new_n1148), .A2(new_n1151), .B1(new_n1098), .B2(new_n793), .ZN(new_n1152));
  OR2_X1    g727(.A1(new_n1151), .A2(new_n1148), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(G171), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1100), .A2(new_n808), .A3(new_n1097), .ZN(new_n1156));
  AOI21_X1  g731(.A(G1966), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1157));
  OAI21_X1  g732(.A(G8), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1005), .A2(G8), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1158), .A2(KEYINPUT51), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT51), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1149), .A2(new_n1093), .A3(new_n1049), .ZN(new_n1162));
  INV_X1    g737(.A(G1966), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1100), .A2(new_n808), .A3(new_n1097), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1161), .B(G8), .C1(new_n1166), .C2(new_n1005), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1159), .ZN(new_n1168));
  AOI21_X1  g743(.A(KEYINPUT124), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT124), .ZN(new_n1170));
  AOI211_X1 g745(.A(new_n1170), .B(new_n1159), .C1(new_n1164), .C2(new_n1165), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1160), .B(new_n1167), .C1(new_n1169), .C2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT62), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1155), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1172), .A2(KEYINPUT62), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(KEYINPUT126), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT126), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1172), .A2(new_n1178), .A3(KEYINPUT62), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1175), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT54), .ZN(new_n1181));
  AND3_X1   g756(.A1(new_n1152), .A2(new_n1153), .A3(G301), .ZN(new_n1182));
  AOI21_X1  g757(.A(G301), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1152), .A2(new_n1153), .A3(G301), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1155), .A2(KEYINPUT54), .A3(new_n1185), .ZN(new_n1186));
  AND3_X1   g761(.A1(new_n1172), .A2(new_n1184), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT61), .ZN(new_n1188));
  XNOR2_X1  g763(.A(KEYINPUT56), .B(G2072), .ZN(new_n1189));
  AND3_X1   g764(.A1(new_n1092), .A2(new_n1093), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(G1956), .B1(new_n1100), .B2(new_n1097), .ZN(new_n1191));
  XNOR2_X1  g766(.A(G299), .B(KEYINPUT57), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1192), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1098), .A2(new_n833), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1092), .A2(new_n1093), .A3(new_n1189), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1194), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1188), .B1(new_n1193), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT59), .ZN(new_n1199));
  INV_X1    g774(.A(new_n560), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1149), .A2(new_n712), .A3(new_n1093), .A4(new_n1049), .ZN(new_n1201));
  XNOR2_X1  g776(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1202), .B(G1341), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1108), .A2(new_n1203), .ZN(new_n1204));
  AOI211_X1 g779(.A(new_n1199), .B(new_n1200), .C1(new_n1201), .C2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1201), .A2(new_n1204), .ZN(new_n1206));
  AOI21_X1  g781(.A(KEYINPUT59), .B1(new_n1206), .B2(new_n560), .ZN(new_n1207));
  NOR2_X1   g782(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1192), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1195), .A2(new_n1194), .A3(new_n1196), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1209), .A2(KEYINPUT61), .A3(new_n1210), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1198), .A2(new_n1208), .A3(new_n1211), .ZN(new_n1212));
  NOR3_X1   g787(.A1(new_n1046), .A2(G2067), .A3(new_n1048), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1213), .B1(new_n1098), .B2(new_n801), .ZN(new_n1214));
  INV_X1    g789(.A(new_n1214), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT60), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g792(.A(KEYINPUT123), .ZN(new_n1218));
  OAI211_X1 g793(.A(new_n1218), .B(new_n625), .C1(new_n1215), .C2(new_n1216), .ZN(new_n1219));
  AOI211_X1 g794(.A(new_n1216), .B(new_n1213), .C1(new_n1098), .C2(new_n801), .ZN(new_n1220));
  OAI21_X1  g795(.A(KEYINPUT123), .B1(new_n1220), .B2(new_n624), .ZN(new_n1221));
  NAND3_X1  g796(.A1(new_n1214), .A2(KEYINPUT60), .A3(new_n624), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT122), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g799(.A1(new_n1220), .A2(KEYINPUT122), .A3(new_n624), .ZN(new_n1225));
  NAND4_X1  g800(.A1(new_n1219), .A2(new_n1221), .A3(new_n1224), .A4(new_n1225), .ZN(new_n1226));
  AOI21_X1  g801(.A(new_n1212), .B1(new_n1217), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1215), .A2(new_n625), .ZN(new_n1228));
  AOI21_X1  g803(.A(new_n1193), .B1(new_n1228), .B2(new_n1209), .ZN(new_n1229));
  OAI21_X1  g804(.A(new_n1187), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g805(.A(new_n1147), .B1(new_n1180), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g806(.A(KEYINPUT120), .ZN(new_n1232));
  NOR2_X1   g807(.A1(new_n1158), .A2(G286), .ZN(new_n1233));
  NAND4_X1  g808(.A1(new_n1132), .A2(new_n1233), .A3(new_n1134), .A4(new_n1136), .ZN(new_n1234));
  OAI21_X1  g809(.A(new_n1232), .B1(new_n1107), .B2(new_n1234), .ZN(new_n1235));
  INV_X1    g810(.A(new_n1234), .ZN(new_n1236));
  NAND3_X1  g811(.A1(new_n1236), .A2(new_n1144), .A3(KEYINPUT120), .ZN(new_n1237));
  INV_X1    g812(.A(KEYINPUT63), .ZN(new_n1238));
  NAND3_X1  g813(.A1(new_n1235), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  NAND2_X1  g814(.A1(new_n1132), .A2(new_n1136), .ZN(new_n1240));
  NAND2_X1  g815(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1241));
  NOR2_X1   g816(.A1(G288), .A2(G1976), .ZN(new_n1242));
  AOI22_X1  g817(.A1(new_n1241), .A2(new_n1242), .B1(new_n1114), .B2(new_n863), .ZN(new_n1243));
  OAI22_X1  g818(.A1(new_n1134), .A2(new_n1240), .B1(new_n1243), .B2(new_n1109), .ZN(new_n1244));
  OAI21_X1  g819(.A(G8), .B1(new_n1133), .B2(new_n1094), .ZN(new_n1245));
  NAND2_X1  g820(.A1(new_n1245), .A2(new_n1089), .ZN(new_n1246));
  NAND2_X1  g821(.A1(new_n1236), .A2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g822(.A(new_n1244), .B1(new_n1247), .B2(KEYINPUT63), .ZN(new_n1248));
  NAND2_X1  g823(.A1(new_n1239), .A2(new_n1248), .ZN(new_n1249));
  OAI21_X1  g824(.A(new_n1086), .B1(new_n1231), .B2(new_n1249), .ZN(new_n1250));
  AND2_X1   g825(.A1(new_n848), .A2(new_n854), .ZN(new_n1251));
  NAND3_X1  g826(.A1(new_n1079), .A2(new_n1073), .A3(new_n1251), .ZN(new_n1252));
  AOI21_X1  g827(.A(new_n1075), .B1(new_n1252), .B2(new_n1065), .ZN(new_n1253));
  NAND2_X1  g828(.A1(new_n1083), .A2(new_n1054), .ZN(new_n1254));
  XNOR2_X1  g829(.A(new_n1254), .B(KEYINPUT48), .ZN(new_n1255));
  NAND4_X1  g830(.A1(new_n1079), .A2(new_n1073), .A3(new_n1081), .A4(new_n1255), .ZN(new_n1256));
  NAND2_X1  g831(.A1(new_n1054), .A2(new_n712), .ZN(new_n1257));
  XNOR2_X1  g832(.A(new_n1257), .B(KEYINPUT46), .ZN(new_n1258));
  OAI21_X1  g833(.A(new_n1059), .B1(new_n754), .B2(new_n1067), .ZN(new_n1259));
  NAND2_X1  g834(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  XNOR2_X1  g835(.A(new_n1260), .B(KEYINPUT47), .ZN(new_n1261));
  NAND2_X1  g836(.A1(new_n1256), .A2(new_n1261), .ZN(new_n1262));
  NOR2_X1   g837(.A1(new_n1253), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g838(.A1(new_n1250), .A2(new_n1263), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g839(.A(G319), .ZN(new_n1266));
  NOR2_X1   g840(.A1(G227), .A2(new_n1266), .ZN(new_n1267));
  NAND4_X1  g841(.A1(new_n692), .A2(new_n741), .A3(new_n745), .A4(new_n1267), .ZN(new_n1268));
  NOR2_X1   g842(.A1(new_n965), .A2(new_n1268), .ZN(new_n1269));
  OAI21_X1  g843(.A(new_n1269), .B1(new_n1038), .B2(new_n1039), .ZN(G225));
  NAND2_X1  g844(.A1(G225), .A2(KEYINPUT127), .ZN(new_n1271));
  INV_X1    g845(.A(KEYINPUT127), .ZN(new_n1272));
  OAI211_X1 g846(.A(new_n1272), .B(new_n1269), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1273));
  NAND2_X1  g847(.A1(new_n1271), .A2(new_n1273), .ZN(G308));
endmodule


