

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588;

  XNOR2_X1 U321 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U322 ( .A(KEYINPUT37), .B(KEYINPUT105), .ZN(n479) );
  XOR2_X1 U323 ( .A(n346), .B(n345), .Z(n573) );
  XNOR2_X1 U324 ( .A(n451), .B(n450), .ZN(n552) );
  AND2_X1 U325 ( .A1(G227GAT), .A2(G233GAT), .ZN(n289) );
  INV_X1 U326 ( .A(KEYINPUT25), .ZN(n463) );
  AND2_X1 U327 ( .A1(n562), .A2(n405), .ZN(n406) );
  AND2_X1 U328 ( .A1(n407), .A2(n406), .ZN(n409) );
  XNOR2_X1 U329 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U330 ( .A(n350), .B(n289), .ZN(n305) );
  XNOR2_X1 U331 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U332 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U333 ( .A(n340), .B(n339), .ZN(n344) );
  XNOR2_X1 U334 ( .A(n480), .B(n479), .ZN(n524) );
  XNOR2_X1 U335 ( .A(KEYINPUT124), .B(n455), .ZN(n568) );
  XOR2_X1 U336 ( .A(n387), .B(n386), .Z(n562) );
  XNOR2_X1 U337 ( .A(n447), .B(n310), .ZN(n536) );
  XNOR2_X1 U338 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n456) );
  XNOR2_X1 U339 ( .A(n484), .B(G43GAT), .ZN(n485) );
  XNOR2_X1 U340 ( .A(n457), .B(n456), .ZN(G1351GAT) );
  XNOR2_X1 U341 ( .A(n486), .B(n485), .ZN(G1330GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT0), .B(G134GAT), .Z(n291) );
  XNOR2_X1 U343 ( .A(KEYINPUT82), .B(G127GAT), .ZN(n290) );
  XNOR2_X1 U344 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U345 ( .A(G113GAT), .B(n292), .Z(n447) );
  XOR2_X1 U346 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n294) );
  XNOR2_X1 U347 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n293) );
  XNOR2_X1 U348 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U349 ( .A(G176GAT), .B(KEYINPUT88), .Z(n296) );
  XNOR2_X1 U350 ( .A(G169GAT), .B(KEYINPUT64), .ZN(n295) );
  XNOR2_X1 U351 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U352 ( .A(n298), .B(n297), .Z(n309) );
  XNOR2_X1 U353 ( .A(KEYINPUT19), .B(KEYINPUT86), .ZN(n299) );
  XNOR2_X1 U354 ( .A(n299), .B(G183GAT), .ZN(n300) );
  XNOR2_X1 U355 ( .A(n300), .B(KEYINPUT87), .ZN(n302) );
  XNOR2_X1 U356 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n301) );
  XNOR2_X1 U357 ( .A(n302), .B(n301), .ZN(n429) );
  XOR2_X1 U358 ( .A(KEYINPUT85), .B(G190GAT), .Z(n304) );
  XNOR2_X1 U359 ( .A(G43GAT), .B(G99GAT), .ZN(n303) );
  XNOR2_X1 U360 ( .A(n304), .B(n303), .ZN(n306) );
  XOR2_X1 U361 ( .A(G120GAT), .B(G71GAT), .Z(n350) );
  XOR2_X1 U362 ( .A(n429), .B(n307), .Z(n308) );
  XNOR2_X1 U363 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U364 ( .A(KEYINPUT21), .B(KEYINPUT91), .Z(n312) );
  XNOR2_X1 U365 ( .A(G218GAT), .B(KEYINPUT90), .ZN(n311) );
  XNOR2_X1 U366 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U367 ( .A(n313), .B(G211GAT), .Z(n315) );
  XNOR2_X1 U368 ( .A(G197GAT), .B(G204GAT), .ZN(n314) );
  XNOR2_X1 U369 ( .A(n315), .B(n314), .ZN(n427) );
  XOR2_X1 U370 ( .A(KEYINPUT3), .B(KEYINPUT92), .Z(n317) );
  XNOR2_X1 U371 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n316) );
  XNOR2_X1 U372 ( .A(n317), .B(n316), .ZN(n440) );
  XOR2_X1 U373 ( .A(G22GAT), .B(G155GAT), .Z(n369) );
  XOR2_X1 U374 ( .A(n440), .B(n369), .Z(n319) );
  NAND2_X1 U375 ( .A1(G228GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U376 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U377 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n321) );
  XNOR2_X1 U378 ( .A(KEYINPUT89), .B(KEYINPUT23), .ZN(n320) );
  XNOR2_X1 U379 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U380 ( .A(n323), .B(n322), .Z(n327) );
  XNOR2_X1 U381 ( .A(G50GAT), .B(KEYINPUT76), .ZN(n324) );
  XNOR2_X1 U382 ( .A(n324), .B(G162GAT), .ZN(n401) );
  XNOR2_X1 U383 ( .A(G106GAT), .B(G78GAT), .ZN(n325) );
  XNOR2_X1 U384 ( .A(n325), .B(G148GAT), .ZN(n359) );
  XNOR2_X1 U385 ( .A(n401), .B(n359), .ZN(n326) );
  XNOR2_X1 U386 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U387 ( .A(n427), .B(n328), .Z(n472) );
  INV_X1 U388 ( .A(KEYINPUT46), .ZN(n365) );
  XOR2_X1 U389 ( .A(G22GAT), .B(G141GAT), .Z(n330) );
  XNOR2_X1 U390 ( .A(G113GAT), .B(G197GAT), .ZN(n329) );
  XNOR2_X1 U391 ( .A(n330), .B(n329), .ZN(n346) );
  XOR2_X1 U392 ( .A(KEYINPUT67), .B(KEYINPUT29), .Z(n332) );
  XNOR2_X1 U393 ( .A(KEYINPUT70), .B(KEYINPUT30), .ZN(n331) );
  XNOR2_X1 U394 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U395 ( .A(G15GAT), .B(G1GAT), .Z(n373) );
  XOR2_X1 U396 ( .A(G36GAT), .B(G50GAT), .Z(n333) );
  XNOR2_X1 U397 ( .A(n373), .B(n333), .ZN(n334) );
  XOR2_X1 U398 ( .A(G169GAT), .B(G8GAT), .Z(n424) );
  XNOR2_X1 U399 ( .A(n334), .B(n424), .ZN(n335) );
  XOR2_X1 U400 ( .A(n336), .B(n335), .Z(n340) );
  NAND2_X1 U401 ( .A1(G229GAT), .A2(G233GAT), .ZN(n338) );
  INV_X1 U402 ( .A(KEYINPUT68), .ZN(n337) );
  XOR2_X1 U403 ( .A(G29GAT), .B(G43GAT), .Z(n342) );
  XNOR2_X1 U404 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n341) );
  XNOR2_X1 U405 ( .A(n342), .B(n341), .ZN(n402) );
  XNOR2_X1 U406 ( .A(n402), .B(KEYINPUT69), .ZN(n343) );
  XNOR2_X1 U407 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U408 ( .A(KEYINPUT72), .B(KEYINPUT74), .Z(n348) );
  XNOR2_X1 U409 ( .A(KEYINPUT33), .B(KEYINPUT32), .ZN(n347) );
  XNOR2_X1 U410 ( .A(n348), .B(n347), .ZN(n363) );
  XNOR2_X1 U411 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n349) );
  XNOR2_X1 U412 ( .A(n349), .B(KEYINPUT71), .ZN(n383) );
  XOR2_X1 U413 ( .A(KEYINPUT75), .B(n383), .Z(n352) );
  XNOR2_X1 U414 ( .A(n350), .B(G204GAT), .ZN(n351) );
  XOR2_X1 U415 ( .A(n352), .B(n351), .Z(n357) );
  XNOR2_X1 U416 ( .A(G99GAT), .B(G85GAT), .ZN(n353) );
  XNOR2_X1 U417 ( .A(n353), .B(KEYINPUT73), .ZN(n394) );
  XOR2_X1 U418 ( .A(n394), .B(KEYINPUT31), .Z(n355) );
  NAND2_X1 U419 ( .A1(G230GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U420 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U421 ( .A(n357), .B(n356), .ZN(n361) );
  XNOR2_X1 U422 ( .A(G176GAT), .B(G92GAT), .ZN(n358) );
  XNOR2_X1 U423 ( .A(n358), .B(G64GAT), .ZN(n419) );
  XNOR2_X1 U424 ( .A(n359), .B(n419), .ZN(n360) );
  XNOR2_X1 U425 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U426 ( .A(n363), .B(n362), .Z(n579) );
  XNOR2_X1 U427 ( .A(KEYINPUT41), .B(n579), .ZN(n540) );
  NAND2_X1 U428 ( .A1(n573), .A2(n540), .ZN(n364) );
  XOR2_X1 U429 ( .A(n365), .B(n364), .Z(n407) );
  XOR2_X1 U430 ( .A(G64GAT), .B(G78GAT), .Z(n367) );
  XNOR2_X1 U431 ( .A(G71GAT), .B(G211GAT), .ZN(n366) );
  XNOR2_X1 U432 ( .A(n367), .B(n366), .ZN(n387) );
  INV_X1 U433 ( .A(G183GAT), .ZN(n368) );
  NAND2_X1 U434 ( .A1(n369), .A2(n368), .ZN(n372) );
  INV_X1 U435 ( .A(n369), .ZN(n370) );
  NAND2_X1 U436 ( .A1(n370), .A2(G183GAT), .ZN(n371) );
  NAND2_X1 U437 ( .A1(n372), .A2(n371), .ZN(n375) );
  XNOR2_X1 U438 ( .A(n373), .B(G127GAT), .ZN(n374) );
  XNOR2_X1 U439 ( .A(n375), .B(n374), .ZN(n381) );
  XOR2_X1 U440 ( .A(KEYINPUT12), .B(KEYINPUT79), .Z(n377) );
  XNOR2_X1 U441 ( .A(G8GAT), .B(KEYINPUT80), .ZN(n376) );
  XNOR2_X1 U442 ( .A(n377), .B(n376), .ZN(n379) );
  AND2_X1 U443 ( .A1(G231GAT), .A2(G233GAT), .ZN(n378) );
  XOR2_X1 U444 ( .A(n382), .B(KEYINPUT15), .Z(n385) );
  XNOR2_X1 U445 ( .A(n383), .B(KEYINPUT14), .ZN(n384) );
  XNOR2_X1 U446 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U447 ( .A(G36GAT), .B(G190GAT), .Z(n420) );
  XOR2_X1 U448 ( .A(KEYINPUT65), .B(G92GAT), .Z(n389) );
  XNOR2_X1 U449 ( .A(G134GAT), .B(G218GAT), .ZN(n388) );
  XNOR2_X1 U450 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U451 ( .A(n420), .B(n390), .ZN(n392) );
  AND2_X1 U452 ( .A1(G232GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U453 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U454 ( .A(n393), .B(KEYINPUT77), .ZN(n396) );
  XOR2_X1 U455 ( .A(n394), .B(KEYINPUT9), .Z(n395) );
  XNOR2_X1 U456 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U457 ( .A(KEYINPUT10), .B(KEYINPUT78), .Z(n398) );
  XNOR2_X1 U458 ( .A(G106GAT), .B(KEYINPUT11), .ZN(n397) );
  XNOR2_X1 U459 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U460 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U461 ( .A(n402), .B(n401), .Z(n403) );
  XNOR2_X1 U462 ( .A(n404), .B(n403), .ZN(n546) );
  INV_X1 U463 ( .A(n546), .ZN(n405) );
  XNOR2_X1 U464 ( .A(KEYINPUT115), .B(KEYINPUT47), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n409), .B(n408), .ZN(n417) );
  XOR2_X1 U466 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n412) );
  INV_X1 U467 ( .A(KEYINPUT36), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n546), .B(n410), .ZN(n586) );
  NOR2_X1 U469 ( .A1(n562), .A2(n586), .ZN(n411) );
  XOR2_X1 U470 ( .A(n412), .B(n411), .Z(n413) );
  NAND2_X1 U471 ( .A1(n579), .A2(n413), .ZN(n414) );
  NOR2_X1 U472 ( .A1(n573), .A2(n414), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n415), .B(KEYINPUT116), .ZN(n416) );
  NOR2_X1 U474 ( .A1(n417), .A2(n416), .ZN(n418) );
  XNOR2_X1 U475 ( .A(KEYINPUT48), .B(n418), .ZN(n535) );
  XNOR2_X1 U476 ( .A(n420), .B(n419), .ZN(n422) );
  AND2_X1 U477 ( .A1(G226GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U478 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n423), .B(KEYINPUT95), .ZN(n426) );
  XOR2_X1 U480 ( .A(n424), .B(KEYINPUT96), .Z(n425) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n428) );
  XNOR2_X1 U482 ( .A(n428), .B(n427), .ZN(n430) );
  XNOR2_X1 U483 ( .A(n430), .B(n429), .ZN(n527) );
  NOR2_X1 U484 ( .A1(n535), .A2(n527), .ZN(n433) );
  XOR2_X1 U485 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n431) );
  XNOR2_X1 U486 ( .A(KEYINPUT54), .B(n431), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n433), .B(n432), .ZN(n452) );
  XOR2_X1 U488 ( .A(KEYINPUT6), .B(KEYINPUT93), .Z(n435) );
  XNOR2_X1 U489 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n434) );
  XNOR2_X1 U490 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U491 ( .A(G155GAT), .B(G148GAT), .Z(n437) );
  XNOR2_X1 U492 ( .A(G29GAT), .B(G120GAT), .ZN(n436) );
  XNOR2_X1 U493 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U494 ( .A(n439), .B(n438), .ZN(n451) );
  XOR2_X1 U495 ( .A(G85GAT), .B(n440), .Z(n442) );
  NAND2_X1 U496 ( .A1(G225GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U498 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n444) );
  XNOR2_X1 U499 ( .A(KEYINPUT94), .B(G57GAT), .ZN(n443) );
  XNOR2_X1 U500 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U501 ( .A(n446), .B(n445), .Z(n449) );
  XNOR2_X1 U502 ( .A(n447), .B(G162GAT), .ZN(n448) );
  XNOR2_X1 U503 ( .A(n449), .B(n448), .ZN(n450) );
  NAND2_X1 U504 ( .A1(n452), .A2(n552), .ZN(n571) );
  NOR2_X1 U505 ( .A1(n472), .A2(n571), .ZN(n453) );
  XNOR2_X1 U506 ( .A(n453), .B(KEYINPUT55), .ZN(n454) );
  NOR2_X1 U507 ( .A1(n536), .A2(n454), .ZN(n455) );
  NAND2_X1 U508 ( .A1(n568), .A2(n546), .ZN(n457) );
  NAND2_X1 U509 ( .A1(n568), .A2(n540), .ZN(n460) );
  XOR2_X1 U510 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n458) );
  XNOR2_X1 U511 ( .A(n458), .B(G176GAT), .ZN(n459) );
  XNOR2_X1 U512 ( .A(n460), .B(n459), .ZN(G1349GAT) );
  NOR2_X1 U513 ( .A1(n536), .A2(n527), .ZN(n461) );
  XNOR2_X1 U514 ( .A(n461), .B(KEYINPUT98), .ZN(n462) );
  NOR2_X1 U515 ( .A1(n462), .A2(n472), .ZN(n464) );
  XNOR2_X1 U516 ( .A(n464), .B(n463), .ZN(n467) );
  XOR2_X1 U517 ( .A(KEYINPUT27), .B(n527), .Z(n473) );
  INV_X1 U518 ( .A(n473), .ZN(n466) );
  NAND2_X1 U519 ( .A1(n536), .A2(n472), .ZN(n465) );
  XNOR2_X1 U520 ( .A(n465), .B(KEYINPUT26), .ZN(n572) );
  NOR2_X1 U521 ( .A1(n466), .A2(n572), .ZN(n554) );
  NOR2_X1 U522 ( .A1(n467), .A2(n554), .ZN(n468) );
  XNOR2_X1 U523 ( .A(n468), .B(KEYINPUT99), .ZN(n469) );
  NAND2_X1 U524 ( .A1(n469), .A2(n552), .ZN(n471) );
  INV_X1 U525 ( .A(KEYINPUT100), .ZN(n470) );
  XNOR2_X1 U526 ( .A(n471), .B(n470), .ZN(n477) );
  XOR2_X1 U527 ( .A(n472), .B(KEYINPUT28), .Z(n531) );
  NAND2_X1 U528 ( .A1(n531), .A2(n473), .ZN(n474) );
  NOR2_X1 U529 ( .A1(n552), .A2(n474), .ZN(n538) );
  NAND2_X1 U530 ( .A1(n538), .A2(n536), .ZN(n475) );
  XNOR2_X1 U531 ( .A(KEYINPUT97), .B(n475), .ZN(n476) );
  NOR2_X1 U532 ( .A1(n477), .A2(n476), .ZN(n493) );
  INV_X1 U533 ( .A(n562), .ZN(n583) );
  OR2_X1 U534 ( .A1(n583), .A2(n586), .ZN(n478) );
  OR2_X1 U535 ( .A1(n493), .A2(n478), .ZN(n480) );
  NAND2_X1 U536 ( .A1(n573), .A2(n579), .ZN(n494) );
  NOR2_X1 U537 ( .A1(n524), .A2(n494), .ZN(n482) );
  INV_X1 U538 ( .A(KEYINPUT106), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U540 ( .A(n483), .B(KEYINPUT38), .ZN(n509) );
  NOR2_X1 U541 ( .A1(n509), .A2(n536), .ZN(n486) );
  INV_X1 U542 ( .A(KEYINPUT40), .ZN(n484) );
  INV_X1 U543 ( .A(G50GAT), .ZN(n489) );
  NOR2_X1 U544 ( .A1(n531), .A2(n509), .ZN(n487) );
  XNOR2_X1 U545 ( .A(KEYINPUT108), .B(n487), .ZN(n488) );
  XNOR2_X1 U546 ( .A(n489), .B(n488), .ZN(G1331GAT) );
  XNOR2_X1 U547 ( .A(KEYINPUT81), .B(KEYINPUT16), .ZN(n491) );
  NOR2_X1 U548 ( .A1(n546), .A2(n562), .ZN(n490) );
  XNOR2_X1 U549 ( .A(n491), .B(n490), .ZN(n492) );
  OR2_X1 U550 ( .A1(n493), .A2(n492), .ZN(n513) );
  NOR2_X1 U551 ( .A1(n494), .A2(n513), .ZN(n495) );
  XNOR2_X1 U552 ( .A(KEYINPUT101), .B(n495), .ZN(n503) );
  NOR2_X1 U553 ( .A1(n552), .A2(n503), .ZN(n497) );
  XNOR2_X1 U554 ( .A(KEYINPUT102), .B(KEYINPUT34), .ZN(n496) );
  XNOR2_X1 U555 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U556 ( .A(G1GAT), .B(n498), .Z(G1324GAT) );
  NOR2_X1 U557 ( .A1(n527), .A2(n503), .ZN(n499) );
  XOR2_X1 U558 ( .A(G8GAT), .B(n499), .Z(G1325GAT) );
  NOR2_X1 U559 ( .A1(n536), .A2(n503), .ZN(n501) );
  XNOR2_X1 U560 ( .A(KEYINPUT103), .B(KEYINPUT35), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U562 ( .A(G15GAT), .B(n502), .Z(G1326GAT) );
  NOR2_X1 U563 ( .A1(n531), .A2(n503), .ZN(n504) );
  XOR2_X1 U564 ( .A(KEYINPUT104), .B(n504), .Z(n505) );
  XNOR2_X1 U565 ( .A(G22GAT), .B(n505), .ZN(G1327GAT) );
  NOR2_X1 U566 ( .A1(n552), .A2(n509), .ZN(n508) );
  XOR2_X1 U567 ( .A(KEYINPUT107), .B(KEYINPUT39), .Z(n506) );
  XNOR2_X1 U568 ( .A(G29GAT), .B(n506), .ZN(n507) );
  XNOR2_X1 U569 ( .A(n508), .B(n507), .ZN(G1328GAT) );
  NOR2_X1 U570 ( .A1(n527), .A2(n509), .ZN(n510) );
  XOR2_X1 U571 ( .A(G36GAT), .B(n510), .Z(G1329GAT) );
  XOR2_X1 U572 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n512) );
  XNOR2_X1 U573 ( .A(G57GAT), .B(KEYINPUT109), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n512), .B(n511), .ZN(n515) );
  INV_X1 U575 ( .A(n573), .ZN(n555) );
  NAND2_X1 U576 ( .A1(n555), .A2(n540), .ZN(n523) );
  OR2_X1 U577 ( .A1(n513), .A2(n523), .ZN(n519) );
  NOR2_X1 U578 ( .A1(n552), .A2(n519), .ZN(n514) );
  XOR2_X1 U579 ( .A(n515), .B(n514), .Z(G1332GAT) );
  NOR2_X1 U580 ( .A1(n527), .A2(n519), .ZN(n516) );
  XOR2_X1 U581 ( .A(G64GAT), .B(n516), .Z(G1333GAT) );
  NOR2_X1 U582 ( .A1(n536), .A2(n519), .ZN(n518) );
  XNOR2_X1 U583 ( .A(G71GAT), .B(KEYINPUT111), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n518), .B(n517), .ZN(G1334GAT) );
  NOR2_X1 U585 ( .A1(n531), .A2(n519), .ZN(n521) );
  XNOR2_X1 U586 ( .A(KEYINPUT43), .B(KEYINPUT112), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U588 ( .A(G78GAT), .B(n522), .ZN(G1335GAT) );
  OR2_X1 U589 ( .A1(n524), .A2(n523), .ZN(n530) );
  NOR2_X1 U590 ( .A1(n552), .A2(n530), .ZN(n526) );
  XNOR2_X1 U591 ( .A(G85GAT), .B(KEYINPUT113), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n526), .B(n525), .ZN(G1336GAT) );
  NOR2_X1 U593 ( .A1(n527), .A2(n530), .ZN(n528) );
  XOR2_X1 U594 ( .A(G92GAT), .B(n528), .Z(G1337GAT) );
  NOR2_X1 U595 ( .A1(n536), .A2(n530), .ZN(n529) );
  XOR2_X1 U596 ( .A(G99GAT), .B(n529), .Z(G1338GAT) );
  NOR2_X1 U597 ( .A1(n531), .A2(n530), .ZN(n533) );
  XNOR2_X1 U598 ( .A(KEYINPUT44), .B(KEYINPUT114), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U600 ( .A(G106GAT), .B(n534), .Z(G1339GAT) );
  NOR2_X1 U601 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U602 ( .A1(n538), .A2(n537), .ZN(n547) );
  NOR2_X1 U603 ( .A1(n555), .A2(n547), .ZN(n539) );
  XOR2_X1 U604 ( .A(G113GAT), .B(n539), .Z(G1340GAT) );
  INV_X1 U605 ( .A(n540), .ZN(n558) );
  NOR2_X1 U606 ( .A1(n558), .A2(n547), .ZN(n542) );
  XNOR2_X1 U607 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(G1341GAT) );
  NOR2_X1 U609 ( .A1(n562), .A2(n547), .ZN(n544) );
  XNOR2_X1 U610 ( .A(KEYINPUT50), .B(KEYINPUT117), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(n545), .ZN(G1342GAT) );
  NOR2_X1 U613 ( .A1(n547), .A2(n405), .ZN(n551) );
  XOR2_X1 U614 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n549) );
  XNOR2_X1 U615 ( .A(G134GAT), .B(KEYINPUT118), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(G1343GAT) );
  NOR2_X1 U618 ( .A1(n552), .A2(n535), .ZN(n553) );
  NAND2_X1 U619 ( .A1(n554), .A2(n553), .ZN(n565) );
  NOR2_X1 U620 ( .A1(n555), .A2(n565), .ZN(n556) );
  XOR2_X1 U621 ( .A(KEYINPUT120), .B(n556), .Z(n557) );
  XNOR2_X1 U622 ( .A(G141GAT), .B(n557), .ZN(G1344GAT) );
  NOR2_X1 U623 ( .A1(n558), .A2(n565), .ZN(n560) );
  XNOR2_X1 U624 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(n561), .ZN(G1345GAT) );
  NOR2_X1 U627 ( .A1(n562), .A2(n565), .ZN(n564) );
  XNOR2_X1 U628 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(G1346GAT) );
  NOR2_X1 U630 ( .A1(n405), .A2(n565), .ZN(n566) );
  XOR2_X1 U631 ( .A(G162GAT), .B(n566), .Z(G1347GAT) );
  NAND2_X1 U632 ( .A1(n573), .A2(n568), .ZN(n567) );
  XNOR2_X1 U633 ( .A(G169GAT), .B(n567), .ZN(G1348GAT) );
  XOR2_X1 U634 ( .A(G183GAT), .B(KEYINPUT125), .Z(n570) );
  NAND2_X1 U635 ( .A1(n568), .A2(n583), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G1350GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT60), .B(KEYINPUT127), .Z(n575) );
  NOR2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n582) );
  NAND2_X1 U639 ( .A1(n582), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XOR2_X1 U641 ( .A(n576), .B(KEYINPUT59), .Z(n578) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .Z(n581) );
  INV_X1 U645 ( .A(n582), .ZN(n585) );
  OR2_X1 U646 ( .A1(n585), .A2(n579), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(G1353GAT) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n584), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U651 ( .A(KEYINPUT62), .B(n587), .Z(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

