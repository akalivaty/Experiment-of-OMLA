

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790;

  XOR2_X1 U378 ( .A(n755), .B(n754), .Z(n382) );
  XOR2_X1 U379 ( .A(n357), .B(n676), .Z(n383) );
  BUF_X1 U380 ( .A(n677), .Z(n357) );
  INV_X1 U381 ( .A(n732), .ZN(n358) );
  NAND2_X1 U382 ( .A1(n400), .A2(n632), .ZN(n465) );
  BUF_X1 U383 ( .A(n694), .Z(n436) );
  XNOR2_X1 U384 ( .A(n698), .B(n490), .ZN(n610) );
  BUF_X2 U385 ( .A(n625), .Z(n698) );
  NAND2_X1 U386 ( .A1(n691), .A2(n690), .ZN(n693) );
  INV_X1 U387 ( .A(G902), .ZN(n527) );
  XNOR2_X1 U388 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n482) );
  XNOR2_X1 U389 ( .A(n359), .B(KEYINPUT19), .ZN(n621) );
  BUF_X1 U390 ( .A(n524), .Z(n373) );
  NAND2_X2 U391 ( .A1(n421), .A2(n453), .ZN(n420) );
  XOR2_X2 U392 ( .A(n528), .B(KEYINPUT88), .Z(n372) );
  XNOR2_X2 U393 ( .A(n356), .B(G131), .ZN(n548) );
  INV_X4 U394 ( .A(KEYINPUT67), .ZN(n356) );
  NAND2_X1 U395 ( .A1(n400), .A2(n722), .ZN(n543) );
  XNOR2_X2 U396 ( .A(n489), .B(G472), .ZN(n625) );
  AND2_X1 U397 ( .A1(n370), .A2(n419), .ZN(n369) );
  XNOR2_X2 U398 ( .A(n532), .B(n531), .ZN(n708) );
  XNOR2_X2 U399 ( .A(n498), .B(KEYINPUT15), .ZN(n671) );
  XNOR2_X1 U400 ( .A(G143), .B(G104), .ZN(n551) );
  INV_X1 U401 ( .A(KEYINPUT4), .ZN(n431) );
  INV_X1 U402 ( .A(G146), .ZN(n508) );
  XNOR2_X1 U403 ( .A(G902), .B(KEYINPUT86), .ZN(n498) );
  INV_X2 U404 ( .A(G953), .ZN(n519) );
  BUF_X1 U405 ( .A(G128), .Z(n433) );
  AND2_X2 U406 ( .A1(n368), .A2(KEYINPUT53), .ZN(n367) );
  AND2_X2 U407 ( .A1(n417), .A2(n374), .ZN(n416) );
  NAND2_X2 U408 ( .A1(n688), .A2(n401), .ZN(n689) );
  AND2_X1 U409 ( .A1(n405), .A2(n459), .ZN(n363) );
  AND2_X1 U410 ( .A1(n458), .A2(n462), .ZN(n457) );
  NAND2_X2 U411 ( .A1(n400), .A2(n577), .ZN(n578) );
  AND2_X1 U412 ( .A1(n599), .A2(n600), .ZN(n738) );
  INV_X1 U413 ( .A(n547), .ZN(n778) );
  OR2_X1 U414 ( .A1(n589), .A2(n588), .ZN(n411) );
  NAND2_X1 U415 ( .A1(n363), .A2(n457), .ZN(n362) );
  NOR2_X1 U416 ( .A1(n604), .A2(n603), .ZN(n365) );
  NAND2_X2 U417 ( .A1(n464), .A2(n597), .ZN(n461) );
  XNOR2_X1 U418 ( .A(n431), .B(G137), .ZN(n430) );
  XNOR2_X1 U419 ( .A(n447), .B(G134), .ZN(n565) );
  INV_X1 U420 ( .A(KEYINPUT22), .ZN(n437) );
  XNOR2_X1 U421 ( .A(n362), .B(KEYINPUT106), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n365), .B(n415), .ZN(n789) );
  XNOR2_X1 U423 ( .A(n444), .B(KEYINPUT42), .ZN(n790) );
  AND2_X1 U424 ( .A1(n721), .A2(n639), .ZN(n444) );
  NOR2_X1 U425 ( .A1(n712), .A2(n442), .ZN(n441) );
  AND2_X1 U426 ( .A1(n436), .A2(n579), .ZN(n580) );
  XNOR2_X1 U427 ( .A(n410), .B(n409), .ZN(n760) );
  XNOR2_X1 U428 ( .A(n478), .B(n477), .ZN(n451) );
  XNOR2_X1 U429 ( .A(n508), .B(G125), .ZN(n521) );
  XNOR2_X2 U430 ( .A(KEYINPUT16), .B(G122), .ZN(n522) );
  XNOR2_X1 U431 ( .A(KEYINPUT87), .B(KEYINPUT83), .ZN(n520) );
  NOR2_X1 U432 ( .A1(n654), .A2(n359), .ZN(n614) );
  XNOR2_X2 U433 ( .A(n360), .B(KEYINPUT82), .ZN(n359) );
  NAND2_X1 U434 ( .A1(n621), .A2(n540), .ZN(n541) );
  NAND2_X2 U435 ( .A1(n371), .A2(n708), .ZN(n360) );
  NAND2_X1 U436 ( .A1(n364), .A2(n361), .ZN(n414) );
  INV_X1 U437 ( .A(n789), .ZN(n364) );
  AND2_X2 U438 ( .A1(n590), .A2(KEYINPUT44), .ZN(n375) );
  NAND2_X1 U439 ( .A1(n369), .A2(n366), .ZN(G75) );
  NAND2_X1 U440 ( .A1(n418), .A2(n367), .ZN(n366) );
  NAND2_X1 U441 ( .A1(n422), .A2(KEYINPUT122), .ZN(n368) );
  NAND2_X1 U442 ( .A1(n420), .A2(n475), .ZN(n370) );
  NAND2_X1 U443 ( .A1(n582), .A2(n580), .ZN(n732) );
  XNOR2_X2 U444 ( .A(n578), .B(n437), .ZN(n582) );
  INV_X1 U445 ( .A(n371), .ZN(n633) );
  XNOR2_X2 U446 ( .A(n529), .B(n372), .ZN(n371) );
  INV_X1 U447 ( .A(n712), .ZN(n462) );
  XNOR2_X1 U448 ( .A(n517), .B(n516), .ZN(n448) );
  INV_X1 U449 ( .A(G469), .ZN(n495) );
  INV_X1 U450 ( .A(KEYINPUT108), .ZN(n413) );
  XNOR2_X1 U451 ( .A(n509), .B(G140), .ZN(n510) );
  INV_X1 U452 ( .A(KEYINPUT10), .ZN(n509) );
  NAND2_X1 U453 ( .A1(n677), .A2(n527), .ZN(n489) );
  XNOR2_X1 U454 ( .A(n559), .B(G475), .ZN(n560) );
  XNOR2_X1 U455 ( .A(n515), .B(n514), .ZN(n690) );
  NOR2_X1 U456 ( .A1(n760), .A2(G902), .ZN(n515) );
  XNOR2_X1 U457 ( .A(KEYINPUT92), .B(KEYINPUT93), .ZN(n505) );
  XOR2_X1 U458 ( .A(G110), .B(G137), .Z(n504) );
  XNOR2_X1 U459 ( .A(G119), .B(n433), .ZN(n503) );
  XNOR2_X1 U460 ( .A(n408), .B(n406), .ZN(n566) );
  XNOR2_X1 U461 ( .A(KEYINPUT66), .B(KEYINPUT8), .ZN(n408) );
  NOR2_X1 U462 ( .A1(n407), .A2(G953), .ZN(n406) );
  INV_X1 U463 ( .A(G234), .ZN(n407) );
  INV_X1 U464 ( .A(n725), .ZN(n455) );
  BUF_X1 U465 ( .A(n690), .Z(n434) );
  NAND2_X1 U466 ( .A1(n389), .A2(n388), .ZN(n387) );
  AND2_X1 U467 ( .A1(n652), .A2(n377), .ZN(n388) );
  XNOR2_X1 U468 ( .A(n499), .B(n435), .ZN(n512) );
  XNOR2_X1 U469 ( .A(n500), .B(KEYINPUT94), .ZN(n435) );
  XOR2_X1 U470 ( .A(KEYINPUT95), .B(KEYINPUT20), .Z(n500) );
  XNOR2_X1 U471 ( .A(n480), .B(KEYINPUT18), .ZN(n479) );
  INV_X1 U472 ( .A(KEYINPUT45), .ZN(n449) );
  NAND2_X1 U473 ( .A1(n416), .A2(n412), .ZN(n450) );
  XNOR2_X1 U474 ( .A(n414), .B(n413), .ZN(n412) );
  XNOR2_X1 U475 ( .A(G116), .B(G107), .ZN(n562) );
  XOR2_X1 U476 ( .A(KEYINPUT105), .B(G122), .Z(n563) );
  XNOR2_X1 U477 ( .A(n492), .B(G140), .ZN(n428) );
  INV_X1 U478 ( .A(n710), .ZN(n439) );
  NOR2_X1 U479 ( .A1(n584), .A2(n610), .ZN(n484) );
  INV_X1 U480 ( .A(KEYINPUT31), .ZN(n466) );
  XNOR2_X1 U481 ( .A(n493), .B(n390), .ZN(n677) );
  XNOR2_X1 U482 ( .A(n487), .B(n391), .ZN(n390) );
  XNOR2_X1 U483 ( .A(n376), .B(n511), .ZN(n410) );
  XNOR2_X1 U484 ( .A(n778), .B(n507), .ZN(n409) );
  AND2_X1 U485 ( .A1(n454), .A2(n519), .ZN(n453) );
  NAND2_X1 U486 ( .A1(n455), .A2(KEYINPUT122), .ZN(n454) );
  INV_X1 U487 ( .A(KEYINPUT40), .ZN(n385) );
  INV_X1 U488 ( .A(KEYINPUT107), .ZN(n415) );
  INV_X1 U489 ( .A(KEYINPUT60), .ZN(n468) );
  NAND2_X1 U490 ( .A1(n471), .A2(n470), .ZN(n469) );
  XNOR2_X1 U491 ( .A(n472), .B(n382), .ZN(n471) );
  INV_X1 U492 ( .A(KEYINPUT56), .ZN(n396) );
  NAND2_X1 U493 ( .A1(n398), .A2(n470), .ZN(n397) );
  XNOR2_X1 U494 ( .A(n399), .B(n381), .ZN(n398) );
  AND2_X1 U495 ( .A1(n594), .A2(n593), .ZN(n374) );
  AND2_X1 U496 ( .A1(n566), .A2(G221), .ZN(n376) );
  AND2_X1 U497 ( .A1(n744), .A2(n624), .ZN(n377) );
  AND2_X1 U498 ( .A1(n725), .A2(n476), .ZN(n378) );
  AND2_X1 U499 ( .A1(n597), .A2(n463), .ZN(n379) );
  XOR2_X1 U500 ( .A(n585), .B(KEYINPUT32), .Z(n380) );
  XOR2_X1 U501 ( .A(n727), .B(n726), .Z(n381) );
  INV_X1 U502 ( .A(n763), .ZN(n470) );
  INV_X1 U503 ( .A(KEYINPUT53), .ZN(n475) );
  AND2_X1 U504 ( .A1(KEYINPUT122), .A2(n475), .ZN(n384) );
  XNOR2_X1 U505 ( .A(n640), .B(G131), .ZN(G33) );
  XNOR2_X1 U506 ( .A(n636), .B(n385), .ZN(n640) );
  NAND2_X1 U507 ( .A1(n386), .A2(n663), .ZN(n667) );
  XNOR2_X1 U508 ( .A(n387), .B(n653), .ZN(n386) );
  INV_X1 U509 ( .A(n642), .ZN(n389) );
  XNOR2_X1 U510 ( .A(n373), .B(n486), .ZN(n391) );
  BUF_X1 U511 ( .A(n491), .Z(n392) );
  BUF_X1 U512 ( .A(n682), .Z(n393) );
  BUF_X1 U513 ( .A(n438), .Z(n394) );
  XNOR2_X1 U514 ( .A(n575), .B(n574), .ZN(n438) );
  BUF_X1 U515 ( .A(n426), .Z(n395) );
  XNOR2_X2 U516 ( .A(n689), .B(KEYINPUT78), .ZN(n456) );
  XNOR2_X1 U517 ( .A(n397), .B(n396), .ZN(G51) );
  NAND2_X1 U518 ( .A1(n759), .A2(G210), .ZN(n399) );
  INV_X2 U519 ( .A(n595), .ZN(n400) );
  AND2_X2 U520 ( .A1(n675), .A2(n401), .ZN(n759) );
  XNOR2_X1 U521 ( .A(n666), .B(KEYINPUT73), .ZN(n401) );
  NAND2_X1 U522 ( .A1(n456), .A2(n378), .ZN(n421) );
  XNOR2_X2 U523 ( .A(n465), .B(KEYINPUT97), .ZN(n464) );
  NAND2_X1 U524 ( .A1(n375), .A2(n402), .ZN(n404) );
  NAND2_X1 U525 ( .A1(n403), .A2(KEYINPUT64), .ZN(n402) );
  INV_X1 U526 ( .A(n592), .ZN(n403) );
  NOR2_X2 U527 ( .A1(n682), .A2(n358), .ZN(n592) );
  NAND2_X1 U528 ( .A1(n404), .A2(n411), .ZN(n417) );
  NAND2_X1 U529 ( .A1(n460), .A2(n461), .ZN(n405) );
  XNOR2_X2 U530 ( .A(n483), .B(n380), .ZN(n682) );
  INV_X1 U531 ( .A(n420), .ZN(n418) );
  NAND2_X1 U532 ( .A1(n422), .A2(n384), .ZN(n419) );
  INV_X1 U533 ( .A(n456), .ZN(n422) );
  XNOR2_X2 U534 ( .A(n765), .B(n525), .ZN(n452) );
  XNOR2_X2 U535 ( .A(n423), .B(n764), .ZN(n525) );
  XNOR2_X2 U536 ( .A(n491), .B(KEYINPUT69), .ZN(n423) );
  XNOR2_X2 U537 ( .A(n474), .B(G101), .ZN(n491) );
  XNOR2_X2 U538 ( .A(n524), .B(n523), .ZN(n765) );
  XNOR2_X2 U539 ( .A(n425), .B(n424), .ZN(n524) );
  XNOR2_X2 U540 ( .A(G119), .B(G116), .ZN(n424) );
  XNOR2_X2 U541 ( .A(n488), .B(G113), .ZN(n425) );
  NOR2_X1 U542 ( .A1(n426), .A2(n463), .ZN(n460) );
  NAND2_X1 U543 ( .A1(n426), .A2(n463), .ZN(n458) );
  NAND2_X1 U544 ( .A1(n395), .A2(n740), .ZN(n741) );
  NAND2_X1 U545 ( .A1(n395), .A2(n738), .ZN(n739) );
  XNOR2_X1 U546 ( .A(n467), .B(n466), .ZN(n426) );
  NAND2_X1 U547 ( .A1(n464), .A2(n379), .ZN(n459) );
  INV_X1 U548 ( .A(n461), .ZN(n427) );
  NAND2_X1 U549 ( .A1(n427), .A2(n740), .ZN(n729) );
  NAND2_X1 U550 ( .A1(n427), .A2(n738), .ZN(n728) );
  XNOR2_X1 U551 ( .A(n525), .B(n428), .ZN(n494) );
  XNOR2_X2 U552 ( .A(n473), .B(G107), .ZN(n764) );
  XNOR2_X2 U553 ( .A(n565), .B(n429), .ZN(n779) );
  XNOR2_X2 U554 ( .A(n548), .B(n430), .ZN(n429) );
  XNOR2_X2 U555 ( .A(G143), .B(G128), .ZN(n447) );
  NOR2_X2 U556 ( .A1(n694), .A2(n693), .ZN(n517) );
  INV_X2 U557 ( .A(KEYINPUT65), .ZN(n474) );
  INV_X2 U558 ( .A(KEYINPUT3), .ZN(n488) );
  NAND2_X1 U559 ( .A1(n582), .A2(n484), .ZN(n483) );
  NAND2_X1 U560 ( .A1(n438), .A2(n732), .ZN(n586) );
  OR2_X2 U561 ( .A1(n438), .A2(KEYINPUT81), .ZN(n590) );
  NAND2_X1 U562 ( .A1(n394), .A2(KEYINPUT81), .ZN(n594) );
  XNOR2_X1 U563 ( .A(n394), .B(G122), .ZN(G24) );
  NAND2_X1 U564 ( .A1(n440), .A2(n439), .ZN(n637) );
  INV_X1 U565 ( .A(n442), .ZN(n440) );
  NAND2_X1 U566 ( .A1(n709), .A2(n708), .ZN(n442) );
  NAND2_X1 U567 ( .A1(n640), .A2(n443), .ZN(n641) );
  INV_X1 U568 ( .A(n790), .ZN(n443) );
  XNOR2_X1 U569 ( .A(n445), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U570 ( .A1(n446), .A2(n470), .ZN(n445) );
  XNOR2_X1 U571 ( .A(n678), .B(n383), .ZN(n446) );
  XNOR2_X1 U572 ( .A(n447), .B(n521), .ZN(n477) );
  NAND2_X1 U573 ( .A1(n448), .A2(n610), .ZN(n518) );
  NAND2_X1 U574 ( .A1(n448), .A2(n698), .ZN(n702) );
  XNOR2_X2 U575 ( .A(n450), .B(n449), .ZN(n769) );
  XNOR2_X2 U576 ( .A(n452), .B(n451), .ZN(n727) );
  INV_X1 U577 ( .A(KEYINPUT98), .ZN(n463) );
  NOR2_X1 U578 ( .A1(n702), .A2(n595), .ZN(n467) );
  XNOR2_X1 U579 ( .A(n469), .B(n468), .ZN(G60) );
  NAND2_X1 U580 ( .A1(n759), .A2(G475), .ZN(n472) );
  XNOR2_X2 U581 ( .A(G110), .B(G104), .ZN(n473) );
  INV_X1 U582 ( .A(KEYINPUT122), .ZN(n476) );
  XNOR2_X1 U583 ( .A(n481), .B(n479), .ZN(n478) );
  NAND2_X1 U584 ( .A1(n519), .A2(G224), .ZN(n480) );
  XNOR2_X1 U585 ( .A(n520), .B(n482), .ZN(n481) );
  NAND2_X1 U586 ( .A1(n582), .A2(n581), .ZN(n604) );
  XOR2_X1 U587 ( .A(n659), .B(KEYINPUT43), .Z(n485) );
  XNOR2_X1 U588 ( .A(n641), .B(KEYINPUT46), .ZN(n642) );
  XNOR2_X1 U589 ( .A(n545), .B(G122), .ZN(n546) );
  INV_X1 U590 ( .A(KEYINPUT2), .ZN(n685) );
  XNOR2_X1 U591 ( .A(n547), .B(n546), .ZN(n550) );
  INV_X1 U592 ( .A(KEYINPUT71), .ZN(n516) );
  INV_X1 U593 ( .A(KEYINPUT36), .ZN(n612) );
  NOR2_X1 U594 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U595 ( .A(n493), .B(n494), .ZN(n747) );
  XNOR2_X1 U596 ( .A(n612), .B(KEYINPUT113), .ZN(n613) );
  XNOR2_X1 U597 ( .A(n561), .B(n560), .ZN(n598) );
  XNOR2_X1 U598 ( .A(n614), .B(n613), .ZN(n615) );
  INV_X1 U599 ( .A(n698), .ZN(n597) );
  XNOR2_X2 U600 ( .A(n779), .B(G146), .ZN(n493) );
  XOR2_X1 U601 ( .A(n392), .B(KEYINPUT5), .Z(n487) );
  NOR2_X1 U602 ( .A1(G953), .A2(G237), .ZN(n544) );
  NAND2_X1 U603 ( .A1(n544), .A2(G210), .ZN(n486) );
  INV_X1 U604 ( .A(KEYINPUT6), .ZN(n490) );
  AND2_X1 U605 ( .A1(G227), .A2(n519), .ZN(n492) );
  NOR2_X1 U606 ( .A1(n747), .A2(G902), .ZN(n496) );
  XNOR2_X2 U607 ( .A(n496), .B(n495), .ZN(n596) );
  INV_X1 U608 ( .A(KEYINPUT1), .ZN(n497) );
  XNOR2_X2 U609 ( .A(n596), .B(n497), .ZN(n694) );
  NAND2_X1 U610 ( .A1(n671), .A2(G234), .ZN(n499) );
  AND2_X1 U611 ( .A1(n512), .A2(G221), .ZN(n502) );
  XNOR2_X1 U612 ( .A(KEYINPUT96), .B(KEYINPUT21), .ZN(n501) );
  XNOR2_X1 U613 ( .A(n502), .B(n501), .ZN(n691) );
  XNOR2_X1 U614 ( .A(n504), .B(n503), .ZN(n511) );
  XOR2_X1 U615 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n506) );
  XOR2_X1 U616 ( .A(n506), .B(n505), .Z(n507) );
  XNOR2_X1 U617 ( .A(n521), .B(n510), .ZN(n547) );
  NAND2_X1 U618 ( .A1(G217), .A2(n512), .ZN(n513) );
  XNOR2_X1 U619 ( .A(KEYINPUT25), .B(n513), .ZN(n514) );
  XNOR2_X2 U620 ( .A(n518), .B(KEYINPUT33), .ZN(n722) );
  XNOR2_X1 U621 ( .A(n522), .B(KEYINPUT70), .ZN(n523) );
  NAND2_X1 U622 ( .A1(n727), .A2(n671), .ZN(n529) );
  INV_X1 U623 ( .A(G237), .ZN(n526) );
  NAND2_X1 U624 ( .A1(n527), .A2(n526), .ZN(n530) );
  NAND2_X1 U625 ( .A1(n530), .A2(G210), .ZN(n528) );
  NAND2_X1 U626 ( .A1(n530), .A2(G214), .ZN(n532) );
  INV_X1 U627 ( .A(KEYINPUT89), .ZN(n531) );
  NAND2_X1 U628 ( .A1(G234), .A2(G237), .ZN(n533) );
  XNOR2_X1 U629 ( .A(n533), .B(KEYINPUT14), .ZN(n535) );
  NAND2_X1 U630 ( .A1(n535), .A2(G952), .ZN(n534) );
  XOR2_X1 U631 ( .A(KEYINPUT90), .B(n534), .Z(n719) );
  NAND2_X1 U632 ( .A1(n719), .A2(n519), .ZN(n608) );
  NAND2_X1 U633 ( .A1(n535), .A2(G902), .ZN(n605) );
  INV_X1 U634 ( .A(n605), .ZN(n536) );
  NOR2_X1 U635 ( .A1(G898), .A2(n519), .ZN(n768) );
  NAND2_X1 U636 ( .A1(n536), .A2(n768), .ZN(n538) );
  INV_X1 U637 ( .A(KEYINPUT91), .ZN(n537) );
  XNOR2_X1 U638 ( .A(n538), .B(n537), .ZN(n539) );
  NAND2_X1 U639 ( .A1(n608), .A2(n539), .ZN(n540) );
  XNOR2_X2 U640 ( .A(n541), .B(KEYINPUT0), .ZN(n595) );
  INV_X1 U641 ( .A(KEYINPUT34), .ZN(n542) );
  XNOR2_X1 U642 ( .A(n543), .B(n542), .ZN(n573) );
  NAND2_X1 U643 ( .A1(G214), .A2(n544), .ZN(n545) );
  XNOR2_X1 U644 ( .A(G113), .B(n548), .ZN(n549) );
  XNOR2_X1 U645 ( .A(n550), .B(n549), .ZN(n558) );
  XOR2_X1 U646 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n552) );
  XNOR2_X1 U647 ( .A(n552), .B(n551), .ZN(n556) );
  XOR2_X1 U648 ( .A(KEYINPUT12), .B(KEYINPUT99), .Z(n554) );
  XNOR2_X1 U649 ( .A(KEYINPUT102), .B(KEYINPUT11), .ZN(n553) );
  XNOR2_X1 U650 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U651 ( .A(n556), .B(n555), .Z(n557) );
  XNOR2_X1 U652 ( .A(n558), .B(n557), .ZN(n753) );
  NOR2_X1 U653 ( .A1(G902), .A2(n753), .ZN(n561) );
  XNOR2_X1 U654 ( .A(KEYINPUT13), .B(KEYINPUT103), .ZN(n559) );
  XNOR2_X1 U655 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U656 ( .A(n565), .B(n564), .Z(n568) );
  NAND2_X1 U657 ( .A1(G217), .A2(n566), .ZN(n567) );
  XNOR2_X1 U658 ( .A(n568), .B(n567), .ZN(n570) );
  XOR2_X1 U659 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n569) );
  XNOR2_X1 U660 ( .A(n570), .B(n569), .ZN(n756) );
  NOR2_X1 U661 ( .A1(G902), .A2(n756), .ZN(n571) );
  XNOR2_X1 U662 ( .A(G478), .B(n571), .ZN(n600) );
  NOR2_X1 U663 ( .A1(n598), .A2(n600), .ZN(n643) );
  XNOR2_X1 U664 ( .A(n643), .B(KEYINPUT74), .ZN(n572) );
  NAND2_X1 U665 ( .A1(n573), .A2(n572), .ZN(n575) );
  INV_X1 U666 ( .A(KEYINPUT35), .ZN(n574) );
  NAND2_X1 U667 ( .A1(n598), .A2(n600), .ZN(n710) );
  INV_X1 U668 ( .A(n691), .ZN(n576) );
  NOR2_X1 U669 ( .A1(n710), .A2(n576), .ZN(n577) );
  NOR2_X1 U670 ( .A1(n698), .A2(n434), .ZN(n579) );
  INV_X1 U671 ( .A(n610), .ZN(n581) );
  INV_X1 U672 ( .A(n436), .ZN(n658) );
  INV_X1 U673 ( .A(n434), .ZN(n583) );
  NAND2_X1 U674 ( .A1(n658), .A2(n583), .ZN(n584) );
  INV_X1 U675 ( .A(KEYINPUT75), .ZN(n585) );
  NOR2_X1 U676 ( .A1(n586), .A2(n682), .ZN(n589) );
  NOR2_X1 U677 ( .A1(KEYINPUT81), .A2(KEYINPUT44), .ZN(n587) );
  NAND2_X1 U678 ( .A1(n587), .A2(KEYINPUT64), .ZN(n588) );
  INV_X1 U679 ( .A(KEYINPUT64), .ZN(n591) );
  NAND2_X1 U680 ( .A1(n592), .A2(n591), .ZN(n593) );
  INV_X1 U681 ( .A(n596), .ZN(n618) );
  NOR2_X1 U682 ( .A1(n693), .A2(n618), .ZN(n632) );
  XOR2_X1 U683 ( .A(KEYINPUT104), .B(n598), .Z(n599) );
  INV_X1 U684 ( .A(n599), .ZN(n602) );
  INV_X1 U685 ( .A(n600), .ZN(n601) );
  NAND2_X1 U686 ( .A1(n602), .A2(n601), .ZN(n661) );
  INV_X1 U687 ( .A(n661), .ZN(n740) );
  NOR2_X1 U688 ( .A1(n738), .A2(n740), .ZN(n712) );
  NAND2_X1 U689 ( .A1(n436), .A2(n434), .ZN(n603) );
  NOR2_X1 U690 ( .A1(G900), .A2(n605), .ZN(n606) );
  NAND2_X1 U691 ( .A1(G953), .A2(n606), .ZN(n607) );
  NAND2_X1 U692 ( .A1(n608), .A2(n607), .ZN(n628) );
  NAND2_X1 U693 ( .A1(n691), .A2(n628), .ZN(n609) );
  NOR2_X1 U694 ( .A1(n434), .A2(n609), .ZN(n616) );
  AND2_X1 U695 ( .A1(n738), .A2(n616), .ZN(n611) );
  NAND2_X1 U696 ( .A1(n611), .A2(n610), .ZN(n654) );
  NAND2_X1 U697 ( .A1(n615), .A2(n658), .ZN(n744) );
  NOR2_X1 U698 ( .A1(KEYINPUT47), .A2(n712), .ZN(n623) );
  AND2_X1 U699 ( .A1(n698), .A2(n616), .ZN(n617) );
  XNOR2_X1 U700 ( .A(n617), .B(KEYINPUT28), .ZN(n620) );
  XOR2_X1 U701 ( .A(n618), .B(KEYINPUT112), .Z(n619) );
  NAND2_X1 U702 ( .A1(n620), .A2(n619), .ZN(n638) );
  INV_X1 U703 ( .A(n621), .ZN(n622) );
  NOR2_X1 U704 ( .A1(n638), .A2(n622), .ZN(n736) );
  NAND2_X1 U705 ( .A1(n623), .A2(n736), .ZN(n624) );
  NAND2_X1 U706 ( .A1(n625), .A2(n708), .ZN(n627) );
  XNOR2_X1 U707 ( .A(KEYINPUT30), .B(KEYINPUT110), .ZN(n626) );
  XNOR2_X1 U708 ( .A(n627), .B(n626), .ZN(n630) );
  INV_X1 U709 ( .A(n628), .ZN(n629) );
  AND2_X1 U710 ( .A1(n632), .A2(n631), .ZN(n644) );
  XNOR2_X1 U711 ( .A(n633), .B(KEYINPUT38), .ZN(n709) );
  AND2_X1 U712 ( .A1(n644), .A2(n709), .ZN(n634) );
  XNOR2_X1 U713 ( .A(n634), .B(KEYINPUT39), .ZN(n660) );
  INV_X1 U714 ( .A(n738), .ZN(n635) );
  NOR2_X1 U715 ( .A1(n660), .A2(n635), .ZN(n636) );
  XNOR2_X1 U716 ( .A(n637), .B(KEYINPUT41), .ZN(n721) );
  INV_X1 U717 ( .A(n638), .ZN(n639) );
  NAND2_X1 U718 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U719 ( .A1(n645), .A2(n633), .ZN(n646) );
  XNOR2_X1 U720 ( .A(n646), .B(KEYINPUT111), .ZN(n788) );
  NAND2_X1 U721 ( .A1(n712), .A2(KEYINPUT47), .ZN(n647) );
  NAND2_X1 U722 ( .A1(n788), .A2(n647), .ZN(n651) );
  INV_X1 U723 ( .A(n736), .ZN(n648) );
  NAND2_X1 U724 ( .A1(n648), .A2(KEYINPUT47), .ZN(n649) );
  XNOR2_X1 U725 ( .A(KEYINPUT77), .B(n649), .ZN(n650) );
  NOR2_X1 U726 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U727 ( .A(KEYINPUT48), .B(KEYINPUT68), .Z(n653) );
  INV_X1 U728 ( .A(n708), .ZN(n655) );
  NOR2_X1 U729 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U730 ( .A(n656), .B(KEYINPUT109), .ZN(n657) );
  NOR2_X1 U731 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U732 ( .A1(n485), .A2(n633), .ZN(n680) );
  NOR2_X1 U733 ( .A1(n661), .A2(n660), .ZN(n746) );
  INV_X1 U734 ( .A(n746), .ZN(n662) );
  AND2_X1 U735 ( .A1(n680), .A2(n662), .ZN(n663) );
  INV_X1 U736 ( .A(n667), .ZN(n664) );
  NAND2_X1 U737 ( .A1(n664), .A2(KEYINPUT2), .ZN(n665) );
  NOR2_X1 U738 ( .A1(n769), .A2(n665), .ZN(n666) );
  INV_X1 U739 ( .A(n769), .ZN(n684) );
  BUF_X1 U740 ( .A(n684), .Z(n670) );
  XNOR2_X2 U741 ( .A(n667), .B(KEYINPUT80), .ZN(n780) );
  XNOR2_X1 U742 ( .A(n780), .B(KEYINPUT72), .ZN(n668) );
  NOR2_X1 U743 ( .A1(n668), .A2(n671), .ZN(n669) );
  NAND2_X1 U744 ( .A1(n670), .A2(n669), .ZN(n674) );
  XNOR2_X1 U745 ( .A(n671), .B(KEYINPUT79), .ZN(n672) );
  NAND2_X1 U746 ( .A1(n672), .A2(KEYINPUT2), .ZN(n673) );
  NAND2_X1 U747 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U748 ( .A1(n759), .A2(G472), .ZN(n678) );
  XOR2_X1 U749 ( .A(KEYINPUT84), .B(KEYINPUT62), .Z(n676) );
  INV_X1 U750 ( .A(G952), .ZN(n679) );
  AND2_X1 U751 ( .A1(n679), .A2(G953), .ZN(n763) );
  XNOR2_X1 U752 ( .A(n680), .B(G140), .ZN(G42) );
  XNOR2_X1 U753 ( .A(G119), .B(KEYINPUT127), .ZN(n681) );
  XNOR2_X1 U754 ( .A(n393), .B(n681), .ZN(G21) );
  INV_X1 U755 ( .A(n780), .ZN(n683) );
  NAND2_X1 U756 ( .A1(n684), .A2(n683), .ZN(n686) );
  NAND2_X1 U757 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U758 ( .A(n687), .B(KEYINPUT76), .ZN(n688) );
  NOR2_X1 U759 ( .A1(n691), .A2(n434), .ZN(n692) );
  XNOR2_X1 U760 ( .A(KEYINPUT49), .B(n692), .ZN(n700) );
  XOR2_X1 U761 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n696) );
  NAND2_X1 U762 ( .A1(n436), .A2(n693), .ZN(n695) );
  XOR2_X1 U763 ( .A(n696), .B(n695), .Z(n697) );
  NOR2_X1 U764 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U765 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U766 ( .A(n701), .B(KEYINPUT118), .ZN(n703) );
  NAND2_X1 U767 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U768 ( .A(n704), .B(KEYINPUT51), .ZN(n705) );
  XNOR2_X1 U769 ( .A(n705), .B(KEYINPUT119), .ZN(n706) );
  NAND2_X1 U770 ( .A1(n706), .A2(n721), .ZN(n707) );
  XNOR2_X1 U771 ( .A(n707), .B(KEYINPUT120), .ZN(n717) );
  NOR2_X1 U772 ( .A1(n709), .A2(n708), .ZN(n711) );
  NOR2_X1 U773 ( .A1(n711), .A2(n710), .ZN(n713) );
  NOR2_X1 U774 ( .A1(n713), .A2(n441), .ZN(n714) );
  XNOR2_X1 U775 ( .A(KEYINPUT121), .B(n714), .ZN(n715) );
  NAND2_X1 U776 ( .A1(n715), .A2(n722), .ZN(n716) );
  NAND2_X1 U777 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U778 ( .A(n718), .B(KEYINPUT52), .ZN(n720) );
  NAND2_X1 U779 ( .A1(n720), .A2(n719), .ZN(n724) );
  NAND2_X1 U780 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U781 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U782 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n726) );
  XNOR2_X1 U783 ( .A(n728), .B(G104), .ZN(G6) );
  XOR2_X1 U784 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n730) );
  XNOR2_X1 U785 ( .A(n730), .B(n729), .ZN(n731) );
  XNOR2_X1 U786 ( .A(G107), .B(n731), .ZN(G9) );
  XOR2_X1 U787 ( .A(G110), .B(n358), .Z(G12) );
  XOR2_X1 U788 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n734) );
  NAND2_X1 U789 ( .A1(n740), .A2(n736), .ZN(n733) );
  XNOR2_X1 U790 ( .A(n734), .B(n733), .ZN(n735) );
  XNOR2_X1 U791 ( .A(n433), .B(n735), .ZN(G30) );
  NAND2_X1 U792 ( .A1(n736), .A2(n738), .ZN(n737) );
  XNOR2_X1 U793 ( .A(n737), .B(G146), .ZN(G48) );
  XNOR2_X1 U794 ( .A(n739), .B(G113), .ZN(G15) );
  XOR2_X1 U795 ( .A(G116), .B(KEYINPUT115), .Z(n742) );
  XNOR2_X1 U796 ( .A(n742), .B(n741), .ZN(G18) );
  XOR2_X1 U797 ( .A(KEYINPUT37), .B(KEYINPUT116), .Z(n743) );
  XNOR2_X1 U798 ( .A(n744), .B(n743), .ZN(n745) );
  XNOR2_X1 U799 ( .A(G125), .B(n745), .ZN(G27) );
  XOR2_X1 U800 ( .A(G134), .B(n746), .Z(G36) );
  XOR2_X1 U801 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n749) );
  XNOR2_X1 U802 ( .A(n747), .B(KEYINPUT123), .ZN(n748) );
  XNOR2_X1 U803 ( .A(n749), .B(n748), .ZN(n751) );
  NAND2_X1 U804 ( .A1(n759), .A2(G469), .ZN(n750) );
  XOR2_X1 U805 ( .A(n751), .B(n750), .Z(n752) );
  NOR2_X1 U806 ( .A1(n763), .A2(n752), .ZN(G54) );
  XNOR2_X1 U807 ( .A(KEYINPUT124), .B(KEYINPUT85), .ZN(n755) );
  XNOR2_X1 U808 ( .A(n753), .B(KEYINPUT59), .ZN(n754) );
  NAND2_X1 U809 ( .A1(n759), .A2(G478), .ZN(n757) );
  XNOR2_X1 U810 ( .A(n757), .B(n756), .ZN(n758) );
  NOR2_X1 U811 ( .A1(n763), .A2(n758), .ZN(G63) );
  NAND2_X1 U812 ( .A1(n759), .A2(G217), .ZN(n761) );
  XNOR2_X1 U813 ( .A(n761), .B(n760), .ZN(n762) );
  NOR2_X1 U814 ( .A1(n763), .A2(n762), .ZN(G66) );
  XNOR2_X1 U815 ( .A(n764), .B(G101), .ZN(n766) );
  XOR2_X1 U816 ( .A(n765), .B(n766), .Z(n767) );
  NOR2_X1 U817 ( .A1(n768), .A2(n767), .ZN(n777) );
  BUF_X1 U818 ( .A(n769), .Z(n770) );
  NOR2_X1 U819 ( .A1(n770), .A2(G953), .ZN(n771) );
  XNOR2_X1 U820 ( .A(n771), .B(KEYINPUT125), .ZN(n775) );
  NAND2_X1 U821 ( .A1(G953), .A2(G224), .ZN(n772) );
  XNOR2_X1 U822 ( .A(KEYINPUT61), .B(n772), .ZN(n773) );
  NAND2_X1 U823 ( .A1(n773), .A2(G898), .ZN(n774) );
  NAND2_X1 U824 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U825 ( .A(n777), .B(n776), .ZN(G69) );
  XOR2_X1 U826 ( .A(n779), .B(n778), .Z(n782) );
  XNOR2_X1 U827 ( .A(n782), .B(n780), .ZN(n781) );
  NAND2_X1 U828 ( .A1(n781), .A2(n519), .ZN(n787) );
  XNOR2_X1 U829 ( .A(n782), .B(G227), .ZN(n783) );
  XNOR2_X1 U830 ( .A(n783), .B(KEYINPUT126), .ZN(n784) );
  NAND2_X1 U831 ( .A1(n784), .A2(G900), .ZN(n785) );
  NAND2_X1 U832 ( .A1(n785), .A2(G953), .ZN(n786) );
  NAND2_X1 U833 ( .A1(n787), .A2(n786), .ZN(G72) );
  XNOR2_X1 U834 ( .A(G143), .B(n788), .ZN(G45) );
  XOR2_X1 U835 ( .A(n789), .B(G101), .Z(G3) );
  XOR2_X1 U836 ( .A(G137), .B(n790), .Z(G39) );
endmodule

