

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U550 ( .A(n690), .ZN(n668) );
  INV_X1 U551 ( .A(KEYINPUT98), .ZN(n674) );
  NOR2_X2 U552 ( .A1(G164), .A2(G1384), .ZN(n633) );
  NOR2_X1 U553 ( .A1(G651), .A2(n545), .ZN(n779) );
  XOR2_X1 U554 ( .A(n745), .B(KEYINPUT105), .Z(n514) );
  NOR2_X1 U555 ( .A1(n916), .A2(n637), .ZN(n648) );
  XNOR2_X1 U556 ( .A(KEYINPUT100), .B(KEYINPUT30), .ZN(n680) );
  XNOR2_X1 U557 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U558 ( .A(KEYINPUT31), .B(KEYINPUT101), .ZN(n686) );
  XNOR2_X1 U559 ( .A(n687), .B(n686), .ZN(n688) );
  NOR2_X2 U560 ( .A1(G2105), .A2(n517), .ZN(n857) );
  NOR2_X1 U561 ( .A1(G651), .A2(G543), .ZN(n783) );
  XOR2_X1 U562 ( .A(KEYINPUT1), .B(n524), .Z(n780) );
  XOR2_X1 U563 ( .A(KEYINPUT17), .B(n515), .Z(n856) );
  NOR2_X1 U564 ( .A1(G2105), .A2(G2104), .ZN(n515) );
  NAND2_X1 U565 ( .A1(n856), .A2(G138), .ZN(n523) );
  INV_X1 U566 ( .A(G2104), .ZN(n517) );
  NAND2_X1 U567 ( .A1(G102), .A2(n857), .ZN(n516) );
  XNOR2_X1 U568 ( .A(KEYINPUT85), .B(n516), .ZN(n521) );
  AND2_X1 U569 ( .A1(n517), .A2(G2105), .ZN(n861) );
  NAND2_X1 U570 ( .A1(G126), .A2(n861), .ZN(n519) );
  AND2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n864) );
  NAND2_X1 U572 ( .A1(G114), .A2(n864), .ZN(n518) );
  NAND2_X1 U573 ( .A1(n519), .A2(n518), .ZN(n520) );
  NOR2_X1 U574 ( .A1(n521), .A2(n520), .ZN(n522) );
  AND2_X1 U575 ( .A1(n523), .A2(n522), .ZN(G164) );
  XOR2_X1 U576 ( .A(KEYINPUT0), .B(G543), .Z(n545) );
  NAND2_X1 U577 ( .A1(n779), .A2(G51), .ZN(n526) );
  XOR2_X1 U578 ( .A(G651), .B(KEYINPUT64), .Z(n529) );
  NOR2_X1 U579 ( .A1(G543), .A2(n529), .ZN(n524) );
  NAND2_X1 U580 ( .A1(G63), .A2(n780), .ZN(n525) );
  NAND2_X1 U581 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U582 ( .A(KEYINPUT6), .B(n527), .ZN(n534) );
  NAND2_X1 U583 ( .A1(n783), .A2(G89), .ZN(n528) );
  XNOR2_X1 U584 ( .A(n528), .B(KEYINPUT4), .ZN(n531) );
  NOR2_X1 U585 ( .A1(n545), .A2(n529), .ZN(n784) );
  NAND2_X1 U586 ( .A1(G76), .A2(n784), .ZN(n530) );
  NAND2_X1 U587 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U588 ( .A(n532), .B(KEYINPUT5), .Z(n533) );
  NOR2_X1 U589 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U590 ( .A(KEYINPUT72), .B(n535), .Z(n536) );
  XNOR2_X1 U591 ( .A(KEYINPUT7), .B(n536), .ZN(G168) );
  XOR2_X1 U592 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U593 ( .A1(n779), .A2(G47), .ZN(n538) );
  NAND2_X1 U594 ( .A1(G60), .A2(n780), .ZN(n537) );
  NAND2_X1 U595 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U596 ( .A(KEYINPUT65), .B(n539), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n784), .A2(G72), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n783), .A2(G85), .ZN(n540) );
  AND2_X1 U599 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U600 ( .A1(n543), .A2(n542), .ZN(G290) );
  NAND2_X1 U601 ( .A1(G49), .A2(n779), .ZN(n544) );
  XNOR2_X1 U602 ( .A(n544), .B(KEYINPUT80), .ZN(n550) );
  NAND2_X1 U603 ( .A1(G87), .A2(n545), .ZN(n547) );
  NAND2_X1 U604 ( .A1(G74), .A2(G651), .ZN(n546) );
  NAND2_X1 U605 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U606 ( .A1(n780), .A2(n548), .ZN(n549) );
  NAND2_X1 U607 ( .A1(n550), .A2(n549), .ZN(G288) );
  NAND2_X1 U608 ( .A1(n783), .A2(G88), .ZN(n552) );
  NAND2_X1 U609 ( .A1(G62), .A2(n780), .ZN(n551) );
  NAND2_X1 U610 ( .A1(n552), .A2(n551), .ZN(n555) );
  NAND2_X1 U611 ( .A1(n779), .A2(G50), .ZN(n553) );
  XOR2_X1 U612 ( .A(KEYINPUT82), .B(n553), .Z(n554) );
  NOR2_X1 U613 ( .A1(n555), .A2(n554), .ZN(n557) );
  NAND2_X1 U614 ( .A1(G75), .A2(n784), .ZN(n556) );
  NAND2_X1 U615 ( .A1(n557), .A2(n556), .ZN(G303) );
  NAND2_X1 U616 ( .A1(G78), .A2(n784), .ZN(n559) );
  NAND2_X1 U617 ( .A1(G65), .A2(n780), .ZN(n558) );
  NAND2_X1 U618 ( .A1(n559), .A2(n558), .ZN(n562) );
  NAND2_X1 U619 ( .A1(G91), .A2(n783), .ZN(n560) );
  XNOR2_X1 U620 ( .A(KEYINPUT67), .B(n560), .ZN(n561) );
  NOR2_X1 U621 ( .A1(n562), .A2(n561), .ZN(n564) );
  NAND2_X1 U622 ( .A1(n779), .A2(G53), .ZN(n563) );
  NAND2_X1 U623 ( .A1(n564), .A2(n563), .ZN(G299) );
  NAND2_X1 U624 ( .A1(n783), .A2(G90), .ZN(n566) );
  NAND2_X1 U625 ( .A1(G77), .A2(n784), .ZN(n565) );
  NAND2_X1 U626 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U627 ( .A(KEYINPUT9), .B(n567), .ZN(n572) );
  NAND2_X1 U628 ( .A1(n779), .A2(G52), .ZN(n569) );
  NAND2_X1 U629 ( .A1(G64), .A2(n780), .ZN(n568) );
  NAND2_X1 U630 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U631 ( .A(KEYINPUT66), .B(n570), .Z(n571) );
  NAND2_X1 U632 ( .A1(n572), .A2(n571), .ZN(G301) );
  NAND2_X1 U633 ( .A1(n784), .A2(G73), .ZN(n573) );
  XOR2_X1 U634 ( .A(KEYINPUT2), .B(n573), .Z(n578) );
  NAND2_X1 U635 ( .A1(n783), .A2(G86), .ZN(n575) );
  NAND2_X1 U636 ( .A1(G61), .A2(n780), .ZN(n574) );
  NAND2_X1 U637 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U638 ( .A(KEYINPUT81), .B(n576), .Z(n577) );
  NOR2_X1 U639 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U640 ( .A1(n779), .A2(G48), .ZN(n579) );
  NAND2_X1 U641 ( .A1(n580), .A2(n579), .ZN(G305) );
  INV_X1 U642 ( .A(G303), .ZN(G166) );
  NAND2_X1 U643 ( .A1(G129), .A2(n861), .ZN(n582) );
  NAND2_X1 U644 ( .A1(G117), .A2(n864), .ZN(n581) );
  NAND2_X1 U645 ( .A1(n582), .A2(n581), .ZN(n586) );
  NAND2_X1 U646 ( .A1(G105), .A2(n857), .ZN(n583) );
  XNOR2_X1 U647 ( .A(n583), .B(KEYINPUT38), .ZN(n584) );
  XNOR2_X1 U648 ( .A(n584), .B(KEYINPUT89), .ZN(n585) );
  NOR2_X1 U649 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U650 ( .A(n587), .B(KEYINPUT90), .ZN(n589) );
  NAND2_X1 U651 ( .A1(G141), .A2(n856), .ZN(n588) );
  NAND2_X1 U652 ( .A1(n589), .A2(n588), .ZN(n869) );
  NAND2_X1 U653 ( .A1(G1996), .A2(n869), .ZN(n599) );
  NAND2_X1 U654 ( .A1(G95), .A2(n857), .ZN(n590) );
  XOR2_X1 U655 ( .A(KEYINPUT88), .B(n590), .Z(n595) );
  NAND2_X1 U656 ( .A1(G119), .A2(n861), .ZN(n592) );
  NAND2_X1 U657 ( .A1(G107), .A2(n864), .ZN(n591) );
  NAND2_X1 U658 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U659 ( .A(KEYINPUT87), .B(n593), .Z(n594) );
  NOR2_X1 U660 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U661 ( .A1(n856), .A2(G131), .ZN(n596) );
  NAND2_X1 U662 ( .A1(n597), .A2(n596), .ZN(n879) );
  NAND2_X1 U663 ( .A1(G1991), .A2(n879), .ZN(n598) );
  NAND2_X1 U664 ( .A1(n599), .A2(n598), .ZN(n939) );
  INV_X1 U665 ( .A(n939), .ZN(n600) );
  XOR2_X1 U666 ( .A(G1986), .B(G290), .Z(n911) );
  NAND2_X1 U667 ( .A1(n600), .A2(n911), .ZN(n608) );
  NAND2_X1 U668 ( .A1(n856), .A2(G137), .ZN(n603) );
  NAND2_X1 U669 ( .A1(G101), .A2(n857), .ZN(n601) );
  XOR2_X1 U670 ( .A(KEYINPUT23), .B(n601), .Z(n602) );
  NAND2_X1 U671 ( .A1(n603), .A2(n602), .ZN(n761) );
  INV_X1 U672 ( .A(G40), .ZN(n606) );
  NAND2_X1 U673 ( .A1(G125), .A2(n861), .ZN(n605) );
  NAND2_X1 U674 ( .A1(G113), .A2(n864), .ZN(n604) );
  NAND2_X1 U675 ( .A1(n605), .A2(n604), .ZN(n760) );
  OR2_X1 U676 ( .A1(n606), .A2(n760), .ZN(n607) );
  OR2_X1 U677 ( .A1(n761), .A2(n607), .ZN(n631) );
  NOR2_X1 U678 ( .A1(n633), .A2(n631), .ZN(n744) );
  NAND2_X1 U679 ( .A1(n608), .A2(n744), .ZN(n619) );
  NAND2_X1 U680 ( .A1(G140), .A2(n856), .ZN(n610) );
  NAND2_X1 U681 ( .A1(G104), .A2(n857), .ZN(n609) );
  NAND2_X1 U682 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U683 ( .A(KEYINPUT34), .B(n611), .ZN(n616) );
  NAND2_X1 U684 ( .A1(G128), .A2(n861), .ZN(n613) );
  NAND2_X1 U685 ( .A1(G116), .A2(n864), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n614) );
  XOR2_X1 U687 ( .A(n614), .B(KEYINPUT35), .Z(n615) );
  NOR2_X1 U688 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U689 ( .A(KEYINPUT36), .B(n617), .Z(n618) );
  XOR2_X1 U690 ( .A(KEYINPUT86), .B(n618), .Z(n881) );
  XNOR2_X1 U691 ( .A(G2067), .B(KEYINPUT37), .ZN(n741) );
  NOR2_X1 U692 ( .A1(n881), .A2(n741), .ZN(n950) );
  NAND2_X1 U693 ( .A1(n950), .A2(n744), .ZN(n739) );
  NAND2_X1 U694 ( .A1(n619), .A2(n739), .ZN(n732) );
  NAND2_X1 U695 ( .A1(G1976), .A2(G288), .ZN(n908) );
  NOR2_X1 U696 ( .A1(G1976), .A2(G288), .ZN(n708) );
  NOR2_X1 U697 ( .A1(G1971), .A2(G303), .ZN(n620) );
  NOR2_X1 U698 ( .A1(n708), .A2(n620), .ZN(n915) );
  NAND2_X1 U699 ( .A1(n780), .A2(G56), .ZN(n621) );
  XOR2_X1 U700 ( .A(KEYINPUT14), .B(n621), .Z(n628) );
  NAND2_X1 U701 ( .A1(G81), .A2(n783), .ZN(n622) );
  XNOR2_X1 U702 ( .A(n622), .B(KEYINPUT68), .ZN(n623) );
  XNOR2_X1 U703 ( .A(n623), .B(KEYINPUT12), .ZN(n625) );
  NAND2_X1 U704 ( .A1(G68), .A2(n784), .ZN(n624) );
  NAND2_X1 U705 ( .A1(n625), .A2(n624), .ZN(n626) );
  XOR2_X1 U706 ( .A(KEYINPUT13), .B(n626), .Z(n627) );
  NOR2_X1 U707 ( .A1(n628), .A2(n627), .ZN(n630) );
  NAND2_X1 U708 ( .A1(n779), .A2(G43), .ZN(n629) );
  NAND2_X1 U709 ( .A1(n630), .A2(n629), .ZN(n916) );
  INV_X1 U710 ( .A(n631), .ZN(n632) );
  NAND2_X2 U711 ( .A1(n633), .A2(n632), .ZN(n690) );
  AND2_X1 U712 ( .A1(n668), .A2(G1996), .ZN(n634) );
  XOR2_X1 U713 ( .A(n634), .B(KEYINPUT26), .Z(n636) );
  NAND2_X1 U714 ( .A1(n690), .A2(G1341), .ZN(n635) );
  NAND2_X1 U715 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U716 ( .A1(n779), .A2(G54), .ZN(n639) );
  NAND2_X1 U717 ( .A1(G79), .A2(n784), .ZN(n638) );
  NAND2_X1 U718 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U719 ( .A(KEYINPUT70), .B(n640), .ZN(n643) );
  NAND2_X1 U720 ( .A1(G66), .A2(n780), .ZN(n641) );
  XNOR2_X1 U721 ( .A(KEYINPUT69), .B(n641), .ZN(n642) );
  NOR2_X1 U722 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U723 ( .A1(n783), .A2(G92), .ZN(n644) );
  NAND2_X1 U724 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X2 U725 ( .A(KEYINPUT15), .B(n646), .ZN(n919) );
  NOR2_X1 U726 ( .A1(n648), .A2(n919), .ZN(n647) );
  XOR2_X1 U727 ( .A(n647), .B(KEYINPUT96), .Z(n656) );
  NAND2_X1 U728 ( .A1(n648), .A2(n919), .ZN(n654) );
  NAND2_X1 U729 ( .A1(G1348), .A2(n690), .ZN(n649) );
  XNOR2_X1 U730 ( .A(n649), .B(KEYINPUT94), .ZN(n651) );
  NAND2_X1 U731 ( .A1(n668), .A2(G2067), .ZN(n650) );
  NAND2_X1 U732 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U733 ( .A(KEYINPUT95), .B(n652), .Z(n653) );
  NAND2_X1 U734 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U735 ( .A1(n656), .A2(n655), .ZN(n662) );
  NAND2_X1 U736 ( .A1(n668), .A2(G2072), .ZN(n657) );
  XOR2_X1 U737 ( .A(KEYINPUT27), .B(n657), .Z(n659) );
  XOR2_X1 U738 ( .A(KEYINPUT93), .B(G1956), .Z(n989) );
  NAND2_X1 U739 ( .A1(n989), .A2(n690), .ZN(n658) );
  NAND2_X1 U740 ( .A1(n659), .A2(n658), .ZN(n663) );
  NOR2_X1 U741 ( .A1(G299), .A2(n663), .ZN(n660) );
  XNOR2_X1 U742 ( .A(n660), .B(KEYINPUT97), .ZN(n661) );
  NAND2_X1 U743 ( .A1(n662), .A2(n661), .ZN(n666) );
  NAND2_X1 U744 ( .A1(G299), .A2(n663), .ZN(n664) );
  XNOR2_X1 U745 ( .A(n664), .B(KEYINPUT28), .ZN(n665) );
  NAND2_X1 U746 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U747 ( .A(KEYINPUT29), .B(n667), .ZN(n673) );
  NAND2_X1 U748 ( .A1(G1961), .A2(n690), .ZN(n670) );
  XOR2_X1 U749 ( .A(G2078), .B(KEYINPUT25), .Z(n961) );
  NAND2_X1 U750 ( .A1(n668), .A2(n961), .ZN(n669) );
  NAND2_X1 U751 ( .A1(n670), .A2(n669), .ZN(n683) );
  NOR2_X1 U752 ( .A1(G301), .A2(n683), .ZN(n671) );
  XNOR2_X1 U753 ( .A(n671), .B(KEYINPUT92), .ZN(n672) );
  NOR2_X1 U754 ( .A1(n673), .A2(n672), .ZN(n675) );
  XNOR2_X1 U755 ( .A(n675), .B(n674), .ZN(n689) );
  INV_X1 U756 ( .A(KEYINPUT99), .ZN(n678) );
  NAND2_X1 U757 ( .A1(n690), .A2(G8), .ZN(n676) );
  XNOR2_X1 U758 ( .A(n676), .B(KEYINPUT91), .ZN(n726) );
  INV_X1 U759 ( .A(n726), .ZN(n711) );
  NOR2_X1 U760 ( .A1(G1966), .A2(n711), .ZN(n702) );
  NOR2_X1 U761 ( .A1(G2084), .A2(n690), .ZN(n699) );
  NOR2_X1 U762 ( .A1(n702), .A2(n699), .ZN(n677) );
  XNOR2_X1 U763 ( .A(n678), .B(n677), .ZN(n679) );
  NAND2_X1 U764 ( .A1(n679), .A2(G8), .ZN(n681) );
  NOR2_X1 U765 ( .A1(G168), .A2(n682), .ZN(n685) );
  AND2_X1 U766 ( .A1(G301), .A2(n683), .ZN(n684) );
  NOR2_X1 U767 ( .A1(n685), .A2(n684), .ZN(n687) );
  NAND2_X1 U768 ( .A1(n689), .A2(n688), .ZN(n700) );
  NAND2_X1 U769 ( .A1(n700), .A2(G286), .ZN(n696) );
  NOR2_X1 U770 ( .A1(G2090), .A2(n690), .ZN(n691) );
  XNOR2_X1 U771 ( .A(n691), .B(KEYINPUT102), .ZN(n693) );
  NOR2_X1 U772 ( .A1(n711), .A2(G1971), .ZN(n692) );
  NOR2_X1 U773 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U774 ( .A1(n694), .A2(G303), .ZN(n695) );
  NAND2_X1 U775 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U776 ( .A1(n697), .A2(G8), .ZN(n698) );
  XNOR2_X1 U777 ( .A(n698), .B(KEYINPUT32), .ZN(n706) );
  NAND2_X1 U778 ( .A1(G8), .A2(n699), .ZN(n704) );
  INV_X1 U779 ( .A(n700), .ZN(n701) );
  NOR2_X1 U780 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U781 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U782 ( .A1(n706), .A2(n705), .ZN(n720) );
  NAND2_X1 U783 ( .A1(n915), .A2(n720), .ZN(n707) );
  NAND2_X1 U784 ( .A1(n908), .A2(n707), .ZN(n713) );
  AND2_X1 U785 ( .A1(n708), .A2(KEYINPUT33), .ZN(n709) );
  AND2_X1 U786 ( .A1(n709), .A2(n726), .ZN(n710) );
  XNOR2_X1 U787 ( .A(G1981), .B(G305), .ZN(n921) );
  OR2_X1 U788 ( .A1(n710), .A2(n921), .ZN(n714) );
  OR2_X1 U789 ( .A1(n711), .A2(n714), .ZN(n712) );
  NOR2_X1 U790 ( .A1(n713), .A2(n712), .ZN(n717) );
  INV_X1 U791 ( .A(n714), .ZN(n715) );
  AND2_X1 U792 ( .A1(n715), .A2(KEYINPUT33), .ZN(n716) );
  NOR2_X1 U793 ( .A1(n717), .A2(n716), .ZN(n730) );
  NOR2_X1 U794 ( .A1(G1981), .A2(G305), .ZN(n718) );
  XNOR2_X1 U795 ( .A(n718), .B(KEYINPUT24), .ZN(n719) );
  AND2_X1 U796 ( .A1(n719), .A2(n726), .ZN(n728) );
  INV_X1 U797 ( .A(n720), .ZN(n724) );
  NAND2_X1 U798 ( .A1(G8), .A2(G166), .ZN(n721) );
  NOR2_X1 U799 ( .A1(G2090), .A2(n721), .ZN(n722) );
  XOR2_X1 U800 ( .A(KEYINPUT103), .B(n722), .Z(n723) );
  NOR2_X1 U801 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U802 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U803 ( .A1(n728), .A2(n727), .ZN(n729) );
  AND2_X1 U804 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U805 ( .A1(n732), .A2(n731), .ZN(n733) );
  INV_X1 U806 ( .A(n733), .ZN(n746) );
  NOR2_X1 U807 ( .A1(G1996), .A2(n869), .ZN(n943) );
  NOR2_X1 U808 ( .A1(G1991), .A2(n879), .ZN(n734) );
  XNOR2_X1 U809 ( .A(KEYINPUT104), .B(n734), .ZN(n938) );
  NOR2_X1 U810 ( .A1(G1986), .A2(G290), .ZN(n735) );
  NOR2_X1 U811 ( .A1(n938), .A2(n735), .ZN(n736) );
  NOR2_X1 U812 ( .A1(n939), .A2(n736), .ZN(n737) );
  NOR2_X1 U813 ( .A1(n943), .A2(n737), .ZN(n738) );
  XNOR2_X1 U814 ( .A(KEYINPUT39), .B(n738), .ZN(n740) );
  NAND2_X1 U815 ( .A1(n740), .A2(n739), .ZN(n742) );
  NAND2_X1 U816 ( .A1(n881), .A2(n741), .ZN(n947) );
  NAND2_X1 U817 ( .A1(n742), .A2(n947), .ZN(n743) );
  NAND2_X1 U818 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U819 ( .A1(n746), .A2(n514), .ZN(n747) );
  XNOR2_X1 U820 ( .A(n747), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U821 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U822 ( .A1(G123), .A2(n861), .ZN(n748) );
  XNOR2_X1 U823 ( .A(n748), .B(KEYINPUT76), .ZN(n749) );
  XNOR2_X1 U824 ( .A(n749), .B(KEYINPUT18), .ZN(n751) );
  NAND2_X1 U825 ( .A1(G135), .A2(n856), .ZN(n750) );
  NAND2_X1 U826 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U827 ( .A(n752), .B(KEYINPUT77), .ZN(n754) );
  NAND2_X1 U828 ( .A1(G99), .A2(n857), .ZN(n753) );
  NAND2_X1 U829 ( .A1(n754), .A2(n753), .ZN(n757) );
  NAND2_X1 U830 ( .A1(n864), .A2(G111), .ZN(n755) );
  XOR2_X1 U831 ( .A(KEYINPUT78), .B(n755), .Z(n756) );
  NOR2_X1 U832 ( .A1(n757), .A2(n756), .ZN(n937) );
  XNOR2_X1 U833 ( .A(n937), .B(G2096), .ZN(n758) );
  XNOR2_X1 U834 ( .A(n758), .B(KEYINPUT79), .ZN(n759) );
  OR2_X1 U835 ( .A1(G2100), .A2(n759), .ZN(G156) );
  INV_X1 U836 ( .A(G132), .ZN(G219) );
  INV_X1 U837 ( .A(G82), .ZN(G220) );
  INV_X1 U838 ( .A(G57), .ZN(G237) );
  NOR2_X1 U839 ( .A1(n761), .A2(n760), .ZN(G160) );
  NAND2_X1 U840 ( .A1(G7), .A2(G661), .ZN(n762) );
  XNOR2_X1 U841 ( .A(n762), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U842 ( .A(G223), .ZN(n815) );
  NAND2_X1 U843 ( .A1(n815), .A2(G567), .ZN(n763) );
  XOR2_X1 U844 ( .A(KEYINPUT11), .B(n763), .Z(G234) );
  INV_X1 U845 ( .A(G860), .ZN(n770) );
  OR2_X1 U846 ( .A1(n916), .A2(n770), .ZN(G153) );
  INV_X1 U847 ( .A(G301), .ZN(G171) );
  NAND2_X1 U848 ( .A1(G868), .A2(G171), .ZN(n765) );
  INV_X1 U849 ( .A(G868), .ZN(n798) );
  NAND2_X1 U850 ( .A1(n919), .A2(n798), .ZN(n764) );
  NAND2_X1 U851 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U852 ( .A(n766), .B(KEYINPUT71), .ZN(G284) );
  NOR2_X1 U853 ( .A1(G286), .A2(n798), .ZN(n767) );
  XOR2_X1 U854 ( .A(KEYINPUT73), .B(n767), .Z(n769) );
  NOR2_X1 U855 ( .A1(G868), .A2(G299), .ZN(n768) );
  NOR2_X1 U856 ( .A1(n769), .A2(n768), .ZN(G297) );
  NAND2_X1 U857 ( .A1(n770), .A2(G559), .ZN(n771) );
  NAND2_X1 U858 ( .A1(n771), .A2(n919), .ZN(n772) );
  XNOR2_X1 U859 ( .A(n772), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U860 ( .A1(n919), .A2(G868), .ZN(n773) );
  NOR2_X1 U861 ( .A1(G559), .A2(n773), .ZN(n774) );
  XNOR2_X1 U862 ( .A(n774), .B(KEYINPUT74), .ZN(n776) );
  NOR2_X1 U863 ( .A1(n916), .A2(G868), .ZN(n775) );
  NOR2_X1 U864 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U865 ( .A(KEYINPUT75), .B(n777), .Z(G282) );
  NAND2_X1 U866 ( .A1(G559), .A2(n919), .ZN(n778) );
  XNOR2_X1 U867 ( .A(n916), .B(n778), .ZN(n796) );
  NOR2_X1 U868 ( .A1(n796), .A2(G860), .ZN(n789) );
  NAND2_X1 U869 ( .A1(n779), .A2(G55), .ZN(n782) );
  NAND2_X1 U870 ( .A1(G67), .A2(n780), .ZN(n781) );
  NAND2_X1 U871 ( .A1(n782), .A2(n781), .ZN(n788) );
  NAND2_X1 U872 ( .A1(n783), .A2(G93), .ZN(n786) );
  NAND2_X1 U873 ( .A1(G80), .A2(n784), .ZN(n785) );
  NAND2_X1 U874 ( .A1(n786), .A2(n785), .ZN(n787) );
  NOR2_X1 U875 ( .A1(n788), .A2(n787), .ZN(n790) );
  XNOR2_X1 U876 ( .A(n789), .B(n790), .ZN(G145) );
  NOR2_X1 U877 ( .A1(G868), .A2(n790), .ZN(n800) );
  XNOR2_X1 U878 ( .A(G305), .B(G290), .ZN(n795) );
  XOR2_X1 U879 ( .A(KEYINPUT19), .B(n790), .Z(n791) );
  XNOR2_X1 U880 ( .A(G288), .B(n791), .ZN(n792) );
  XNOR2_X1 U881 ( .A(G166), .B(n792), .ZN(n793) );
  XNOR2_X1 U882 ( .A(n793), .B(G299), .ZN(n794) );
  XNOR2_X1 U883 ( .A(n795), .B(n794), .ZN(n887) );
  XOR2_X1 U884 ( .A(n796), .B(n887), .Z(n797) );
  NOR2_X1 U885 ( .A1(n798), .A2(n797), .ZN(n799) );
  NOR2_X1 U886 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U887 ( .A(n801), .B(KEYINPUT83), .ZN(G295) );
  NAND2_X1 U888 ( .A1(G2084), .A2(G2078), .ZN(n802) );
  XOR2_X1 U889 ( .A(KEYINPUT20), .B(n802), .Z(n803) );
  NAND2_X1 U890 ( .A1(G2090), .A2(n803), .ZN(n804) );
  XNOR2_X1 U891 ( .A(KEYINPUT21), .B(n804), .ZN(n805) );
  NAND2_X1 U892 ( .A1(n805), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U893 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U894 ( .A1(G69), .A2(G120), .ZN(n806) );
  NOR2_X1 U895 ( .A1(G237), .A2(n806), .ZN(n807) );
  NAND2_X1 U896 ( .A1(G108), .A2(n807), .ZN(n819) );
  NAND2_X1 U897 ( .A1(G567), .A2(n819), .ZN(n808) );
  XNOR2_X1 U898 ( .A(n808), .B(KEYINPUT84), .ZN(n813) );
  NOR2_X1 U899 ( .A1(G220), .A2(G219), .ZN(n809) );
  XOR2_X1 U900 ( .A(KEYINPUT22), .B(n809), .Z(n810) );
  NOR2_X1 U901 ( .A1(G218), .A2(n810), .ZN(n811) );
  NAND2_X1 U902 ( .A1(G96), .A2(n811), .ZN(n820) );
  NAND2_X1 U903 ( .A1(G2106), .A2(n820), .ZN(n812) );
  NAND2_X1 U904 ( .A1(n813), .A2(n812), .ZN(n821) );
  NAND2_X1 U905 ( .A1(G483), .A2(G661), .ZN(n814) );
  NOR2_X1 U906 ( .A1(n821), .A2(n814), .ZN(n818) );
  NAND2_X1 U907 ( .A1(n818), .A2(G36), .ZN(G176) );
  NAND2_X1 U908 ( .A1(G2106), .A2(n815), .ZN(G217) );
  AND2_X1 U909 ( .A1(G15), .A2(G2), .ZN(n816) );
  NAND2_X1 U910 ( .A1(G661), .A2(n816), .ZN(G259) );
  NAND2_X1 U911 ( .A1(G3), .A2(G1), .ZN(n817) );
  NAND2_X1 U912 ( .A1(n818), .A2(n817), .ZN(G188) );
  XOR2_X1 U913 ( .A(G96), .B(KEYINPUT106), .Z(G221) );
  INV_X1 U915 ( .A(G120), .ZN(G236) );
  INV_X1 U916 ( .A(G69), .ZN(G235) );
  NOR2_X1 U917 ( .A1(n820), .A2(n819), .ZN(G325) );
  INV_X1 U918 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U919 ( .A(KEYINPUT107), .B(n821), .ZN(G319) );
  XOR2_X1 U920 ( .A(G2100), .B(G2096), .Z(n823) );
  XNOR2_X1 U921 ( .A(KEYINPUT42), .B(G2678), .ZN(n822) );
  XNOR2_X1 U922 ( .A(n823), .B(n822), .ZN(n827) );
  XOR2_X1 U923 ( .A(KEYINPUT43), .B(G2090), .Z(n825) );
  XNOR2_X1 U924 ( .A(G2067), .B(G2072), .ZN(n824) );
  XNOR2_X1 U925 ( .A(n825), .B(n824), .ZN(n826) );
  XOR2_X1 U926 ( .A(n827), .B(n826), .Z(n829) );
  XNOR2_X1 U927 ( .A(G2084), .B(G2078), .ZN(n828) );
  XNOR2_X1 U928 ( .A(n829), .B(n828), .ZN(G227) );
  XOR2_X1 U929 ( .A(G1976), .B(G1971), .Z(n831) );
  XNOR2_X1 U930 ( .A(G1966), .B(G1961), .ZN(n830) );
  XNOR2_X1 U931 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U932 ( .A(n832), .B(G2474), .Z(n834) );
  XNOR2_X1 U933 ( .A(G1996), .B(G1991), .ZN(n833) );
  XNOR2_X1 U934 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U935 ( .A(KEYINPUT41), .B(G1986), .Z(n836) );
  XNOR2_X1 U936 ( .A(G1956), .B(G1981), .ZN(n835) );
  XNOR2_X1 U937 ( .A(n836), .B(n835), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(G229) );
  NAND2_X1 U939 ( .A1(G112), .A2(n864), .ZN(n840) );
  NAND2_X1 U940 ( .A1(G100), .A2(n857), .ZN(n839) );
  NAND2_X1 U941 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U942 ( .A(KEYINPUT108), .B(n841), .ZN(n846) );
  NAND2_X1 U943 ( .A1(n861), .A2(G124), .ZN(n842) );
  XNOR2_X1 U944 ( .A(n842), .B(KEYINPUT44), .ZN(n844) );
  NAND2_X1 U945 ( .A1(G136), .A2(n856), .ZN(n843) );
  NAND2_X1 U946 ( .A1(n844), .A2(n843), .ZN(n845) );
  NOR2_X1 U947 ( .A1(n846), .A2(n845), .ZN(G162) );
  NAND2_X1 U948 ( .A1(G127), .A2(n861), .ZN(n848) );
  NAND2_X1 U949 ( .A1(G115), .A2(n864), .ZN(n847) );
  NAND2_X1 U950 ( .A1(n848), .A2(n847), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n849), .B(KEYINPUT47), .ZN(n851) );
  NAND2_X1 U952 ( .A1(G139), .A2(n856), .ZN(n850) );
  NAND2_X1 U953 ( .A1(n851), .A2(n850), .ZN(n854) );
  NAND2_X1 U954 ( .A1(n857), .A2(G103), .ZN(n852) );
  XOR2_X1 U955 ( .A(KEYINPUT112), .B(n852), .Z(n853) );
  NOR2_X1 U956 ( .A1(n854), .A2(n853), .ZN(n855) );
  XOR2_X1 U957 ( .A(KEYINPUT113), .B(n855), .Z(n932) );
  NAND2_X1 U958 ( .A1(G142), .A2(n856), .ZN(n859) );
  NAND2_X1 U959 ( .A1(G106), .A2(n857), .ZN(n858) );
  NAND2_X1 U960 ( .A1(n859), .A2(n858), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n860), .B(KEYINPUT45), .ZN(n863) );
  NAND2_X1 U962 ( .A1(G130), .A2(n861), .ZN(n862) );
  NAND2_X1 U963 ( .A1(n863), .A2(n862), .ZN(n867) );
  NAND2_X1 U964 ( .A1(G118), .A2(n864), .ZN(n865) );
  XNOR2_X1 U965 ( .A(KEYINPUT109), .B(n865), .ZN(n866) );
  NOR2_X1 U966 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U967 ( .A(n932), .B(n868), .ZN(n871) );
  XNOR2_X1 U968 ( .A(n869), .B(n937), .ZN(n870) );
  XNOR2_X1 U969 ( .A(n871), .B(n870), .ZN(n883) );
  XOR2_X1 U970 ( .A(KEYINPUT110), .B(KEYINPUT114), .Z(n873) );
  XNOR2_X1 U971 ( .A(KEYINPUT111), .B(KEYINPUT48), .ZN(n872) );
  XNOR2_X1 U972 ( .A(n873), .B(n872), .ZN(n874) );
  XOR2_X1 U973 ( .A(n874), .B(KEYINPUT46), .Z(n876) );
  XNOR2_X1 U974 ( .A(G160), .B(G162), .ZN(n875) );
  XNOR2_X1 U975 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U976 ( .A(G164), .B(n877), .Z(n878) );
  XNOR2_X1 U977 ( .A(n879), .B(n878), .ZN(n880) );
  XNOR2_X1 U978 ( .A(n881), .B(n880), .ZN(n882) );
  XNOR2_X1 U979 ( .A(n883), .B(n882), .ZN(n884) );
  NOR2_X1 U980 ( .A1(G37), .A2(n884), .ZN(G395) );
  XNOR2_X1 U981 ( .A(n916), .B(KEYINPUT115), .ZN(n886) );
  XNOR2_X1 U982 ( .A(G171), .B(n919), .ZN(n885) );
  XNOR2_X1 U983 ( .A(n886), .B(n885), .ZN(n888) );
  XNOR2_X1 U984 ( .A(n888), .B(n887), .ZN(n889) );
  XNOR2_X1 U985 ( .A(n889), .B(G286), .ZN(n890) );
  NOR2_X1 U986 ( .A1(G37), .A2(n890), .ZN(G397) );
  XOR2_X1 U987 ( .A(G2451), .B(G2430), .Z(n892) );
  XNOR2_X1 U988 ( .A(G2438), .B(G2443), .ZN(n891) );
  XNOR2_X1 U989 ( .A(n892), .B(n891), .ZN(n898) );
  XOR2_X1 U990 ( .A(G2435), .B(G2454), .Z(n894) );
  XNOR2_X1 U991 ( .A(G1341), .B(G1348), .ZN(n893) );
  XNOR2_X1 U992 ( .A(n894), .B(n893), .ZN(n896) );
  XOR2_X1 U993 ( .A(G2446), .B(G2427), .Z(n895) );
  XNOR2_X1 U994 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U995 ( .A(n898), .B(n897), .Z(n899) );
  NAND2_X1 U996 ( .A1(G14), .A2(n899), .ZN(n905) );
  NAND2_X1 U997 ( .A1(G319), .A2(n905), .ZN(n902) );
  NOR2_X1 U998 ( .A1(G227), .A2(G229), .ZN(n900) );
  XNOR2_X1 U999 ( .A(KEYINPUT49), .B(n900), .ZN(n901) );
  NOR2_X1 U1000 ( .A1(n902), .A2(n901), .ZN(n904) );
  NOR2_X1 U1001 ( .A1(G395), .A2(G397), .ZN(n903) );
  NAND2_X1 U1002 ( .A1(n904), .A2(n903), .ZN(G225) );
  INV_X1 U1003 ( .A(G225), .ZN(G308) );
  INV_X1 U1004 ( .A(G108), .ZN(G238) );
  INV_X1 U1005 ( .A(n905), .ZN(G401) );
  XNOR2_X1 U1006 ( .A(G16), .B(KEYINPUT121), .ZN(n906) );
  XNOR2_X1 U1007 ( .A(n906), .B(KEYINPUT56), .ZN(n931) );
  NAND2_X1 U1008 ( .A1(G1971), .A2(G303), .ZN(n907) );
  NAND2_X1 U1009 ( .A1(n908), .A2(n907), .ZN(n913) );
  XOR2_X1 U1010 ( .A(G1956), .B(KEYINPUT122), .Z(n909) );
  XNOR2_X1 U1011 ( .A(G299), .B(n909), .ZN(n910) );
  NAND2_X1 U1012 ( .A1(n911), .A2(n910), .ZN(n912) );
  NOR2_X1 U1013 ( .A1(n913), .A2(n912), .ZN(n914) );
  NAND2_X1 U1014 ( .A1(n915), .A2(n914), .ZN(n928) );
  XNOR2_X1 U1015 ( .A(G301), .B(G1961), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(n916), .B(G1341), .ZN(n917) );
  NOR2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n926) );
  XOR2_X1 U1018 ( .A(n919), .B(G1348), .Z(n924) );
  XOR2_X1 U1019 ( .A(G1966), .B(G168), .Z(n920) );
  NOR2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(KEYINPUT57), .B(n922), .ZN(n923) );
  NOR2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1024 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1025 ( .A(KEYINPUT123), .B(n929), .Z(n930) );
  NOR2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n1013) );
  XNOR2_X1 U1027 ( .A(KEYINPUT117), .B(KEYINPUT52), .ZN(n955) );
  XOR2_X1 U1028 ( .A(G2072), .B(n932), .Z(n934) );
  XOR2_X1 U1029 ( .A(G164), .B(G2078), .Z(n933) );
  NOR2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1031 ( .A(KEYINPUT50), .B(n935), .ZN(n953) );
  XOR2_X1 U1032 ( .A(G2084), .B(G160), .Z(n936) );
  NOR2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n941) );
  NOR2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n946) );
  XOR2_X1 U1036 ( .A(G2090), .B(G162), .Z(n942) );
  NOR2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(n944), .B(KEYINPUT51), .ZN(n945) );
  NOR2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n948) );
  NAND2_X1 U1040 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1041 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1042 ( .A(KEYINPUT116), .B(n951), .ZN(n952) );
  NAND2_X1 U1043 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1044 ( .A(n955), .B(n954), .ZN(n956) );
  INV_X1 U1045 ( .A(KEYINPUT55), .ZN(n1005) );
  NAND2_X1 U1046 ( .A1(n956), .A2(n1005), .ZN(n957) );
  NAND2_X1 U1047 ( .A1(n957), .A2(G29), .ZN(n1011) );
  XNOR2_X1 U1048 ( .A(G2090), .B(G35), .ZN(n973) );
  XNOR2_X1 U1049 ( .A(G2067), .B(G26), .ZN(n959) );
  XNOR2_X1 U1050 ( .A(G2072), .B(G33), .ZN(n958) );
  NOR2_X1 U1051 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1052 ( .A(KEYINPUT119), .B(n960), .Z(n966) );
  XNOR2_X1 U1053 ( .A(n961), .B(G27), .ZN(n963) );
  XNOR2_X1 U1054 ( .A(G32), .B(G1996), .ZN(n962) );
  NOR2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(KEYINPUT120), .B(n964), .ZN(n965) );
  NAND2_X1 U1057 ( .A1(n966), .A2(n965), .ZN(n970) );
  XOR2_X1 U1058 ( .A(G1991), .B(G25), .Z(n967) );
  NAND2_X1 U1059 ( .A1(n967), .A2(G28), .ZN(n968) );
  XNOR2_X1 U1060 ( .A(KEYINPUT118), .B(n968), .ZN(n969) );
  NOR2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1062 ( .A(KEYINPUT53), .B(n971), .ZN(n972) );
  NOR2_X1 U1063 ( .A1(n973), .A2(n972), .ZN(n976) );
  XOR2_X1 U1064 ( .A(G2084), .B(G34), .Z(n974) );
  XNOR2_X1 U1065 ( .A(KEYINPUT54), .B(n974), .ZN(n975) );
  NAND2_X1 U1066 ( .A1(n976), .A2(n975), .ZN(n1004) );
  NOR2_X1 U1067 ( .A1(G29), .A2(KEYINPUT55), .ZN(n977) );
  NAND2_X1 U1068 ( .A1(n1004), .A2(n977), .ZN(n978) );
  NAND2_X1 U1069 ( .A1(G11), .A2(n978), .ZN(n1009) );
  XOR2_X1 U1070 ( .A(G16), .B(KEYINPUT124), .Z(n1003) );
  XNOR2_X1 U1071 ( .A(G1971), .B(G22), .ZN(n980) );
  XNOR2_X1 U1072 ( .A(G1976), .B(G23), .ZN(n979) );
  NOR2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1074 ( .A(KEYINPUT126), .B(n981), .Z(n983) );
  XNOR2_X1 U1075 ( .A(G1986), .B(G24), .ZN(n982) );
  NOR2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1077 ( .A(KEYINPUT58), .B(n984), .ZN(n988) );
  XNOR2_X1 U1078 ( .A(G1966), .B(G21), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(G1961), .B(G5), .ZN(n985) );
  NOR2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n1000) );
  XNOR2_X1 U1082 ( .A(n989), .B(G20), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(G1341), .B(G19), .ZN(n991) );
  XNOR2_X1 U1084 ( .A(G1981), .B(G6), .ZN(n990) );
  NOR2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1086 ( .A(KEYINPUT125), .B(n992), .ZN(n993) );
  NOR2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n997) );
  XNOR2_X1 U1088 ( .A(G1348), .B(KEYINPUT59), .ZN(n995) );
  XNOR2_X1 U1089 ( .A(n995), .B(G4), .ZN(n996) );
  NAND2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1091 ( .A(KEYINPUT60), .B(n998), .ZN(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1093 ( .A(n1001), .B(KEYINPUT61), .ZN(n1002) );
  NAND2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1007) );
  OR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1100 ( .A(KEYINPUT127), .B(n1014), .Z(n1015) );
  XNOR2_X1 U1101 ( .A(KEYINPUT62), .B(n1015), .ZN(G311) );
  INV_X1 U1102 ( .A(G311), .ZN(G150) );
endmodule

