//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 1 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076;
  NOR2_X1   g000(.A1(G237), .A2(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G210), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT27), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT26), .B(G101), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G116), .ZN(new_n194));
  INV_X1    g008(.A(G116), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G119), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT2), .B(G113), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT68), .ZN(new_n199));
  AND3_X1   g013(.A1(new_n197), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n198), .B1(new_n199), .B2(new_n197), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  AND2_X1   g016(.A1(KEYINPUT64), .A2(G131), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT64), .A2(G131), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT11), .ZN(new_n206));
  INV_X1    g020(.A(G134), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G137), .ZN(new_n208));
  INV_X1    g022(.A(G137), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(KEYINPUT11), .A3(G134), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n207), .A2(G137), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n205), .A2(new_n208), .A3(new_n210), .A4(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n208), .A2(new_n210), .A3(new_n211), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n213), .A2(KEYINPUT65), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT65), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n208), .A2(new_n210), .A3(new_n215), .A4(new_n211), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G131), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n212), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G143), .ZN(new_n220));
  INV_X1    g034(.A(G143), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G146), .ZN(new_n222));
  NAND2_X1  g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n220), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n220), .A2(new_n222), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  OR2_X1    g040(.A1(KEYINPUT0), .A2(G128), .ZN(new_n227));
  AND2_X1   g041(.A1(new_n227), .A2(new_n223), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n224), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n218), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G128), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n232), .A2(new_n220), .A3(new_n222), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT1), .B1(new_n221), .B2(G146), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  OAI211_X1 g050(.A(KEYINPUT67), .B(KEYINPUT1), .C1(new_n221), .C2(G146), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(G128), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n233), .B1(new_n238), .B2(new_n225), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n240), .B1(new_n207), .B2(G137), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n209), .A2(KEYINPUT66), .A3(G134), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(new_n211), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G131), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(new_n212), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT69), .B1(new_n239), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n237), .A2(G128), .ZN(new_n247));
  AOI21_X1  g061(.A(KEYINPUT67), .B1(new_n220), .B2(KEYINPUT1), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n225), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n232), .A2(new_n220), .A3(new_n222), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n208), .A2(new_n210), .A3(new_n211), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n253), .A2(new_n205), .B1(new_n243), .B2(G131), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n251), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n230), .A2(new_n246), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT30), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT30), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n251), .A2(new_n254), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n230), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n202), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n230), .A2(new_n246), .A3(new_n202), .A4(new_n255), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n192), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT28), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n212), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n216), .A2(G131), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n213), .A2(KEYINPUT65), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n229), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n259), .B(new_n202), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n265), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n230), .A2(new_n259), .ZN(new_n275));
  INV_X1    g089(.A(new_n202), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n267), .A2(new_n274), .A3(new_n277), .A4(new_n191), .ZN(new_n278));
  AOI21_X1  g092(.A(KEYINPUT71), .B1(new_n264), .B2(new_n278), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n274), .B(new_n277), .C1(new_n265), .C2(new_n262), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT71), .B1(new_n280), .B2(new_n192), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT29), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n256), .A2(new_n276), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(KEYINPUT72), .A3(new_n262), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n256), .A2(new_n287), .A3(new_n276), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n286), .A2(KEYINPUT28), .A3(new_n288), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n289), .A2(KEYINPUT29), .A3(new_n274), .A4(new_n191), .ZN(new_n290));
  INV_X1    g104(.A(G902), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(G472), .B1(new_n284), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(G472), .A2(G902), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT70), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n280), .A2(new_n296), .A3(new_n192), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n296), .B1(new_n280), .B2(new_n192), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n262), .A2(new_n191), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n230), .A2(new_n258), .A3(new_n259), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n302), .B1(KEYINPUT30), .B2(new_n256), .ZN(new_n303));
  OAI211_X1 g117(.A(KEYINPUT31), .B(new_n301), .C1(new_n303), .C2(new_n202), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT31), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n305), .B1(new_n261), .B2(new_n300), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  AOI211_X1 g121(.A(KEYINPUT32), .B(new_n295), .C1(new_n299), .C2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT32), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n274), .A2(new_n277), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n192), .B1(new_n310), .B2(new_n266), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT70), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n280), .A2(new_n296), .A3(new_n192), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n257), .A2(new_n260), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n276), .ZN(new_n315));
  AOI21_X1  g129(.A(KEYINPUT31), .B1(new_n315), .B2(new_n301), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n261), .A2(new_n305), .A3(new_n300), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n312), .B(new_n313), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n309), .B1(new_n318), .B2(new_n294), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n293), .B1(new_n308), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(G110), .B(G122), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G104), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT3), .B1(new_n323), .B2(G107), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT3), .ZN(new_n325));
  INV_X1    g139(.A(G107), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(new_n326), .A3(G104), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n323), .A2(G107), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n324), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT4), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n330), .A3(G101), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n331), .B1(new_n200), .B2(new_n201), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n329), .A2(new_n333), .A3(G101), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n333), .B1(new_n329), .B2(G101), .ZN(new_n335));
  INV_X1    g149(.A(G101), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n324), .A2(new_n327), .A3(new_n336), .A4(new_n328), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT4), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n332), .B1(new_n334), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n323), .A2(G107), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n326), .A2(G104), .ZN(new_n342));
  OAI21_X1  g156(.A(G101), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n337), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT80), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT80), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n337), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(G116), .B(G119), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT5), .ZN(new_n349));
  INV_X1    g163(.A(G113), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n195), .A2(G119), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT5), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n198), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n349), .A2(new_n353), .B1(new_n354), .B2(new_n348), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n345), .A2(new_n347), .A3(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n322), .B1(new_n340), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n345), .A2(new_n347), .A3(new_n355), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n329), .A2(new_n333), .A3(G101), .ZN(new_n359));
  NOR3_X1   g173(.A1(new_n359), .A2(new_n335), .A3(new_n338), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n358), .B(new_n321), .C1(new_n360), .C2(new_n332), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n357), .A2(KEYINPUT83), .A3(KEYINPUT6), .A4(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(KEYINPUT6), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n329), .A2(G101), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT77), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n365), .A2(KEYINPUT4), .A3(new_n337), .A4(new_n334), .ZN(new_n366));
  INV_X1    g180(.A(new_n364), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n354), .B1(KEYINPUT68), .B2(new_n348), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n197), .A2(new_n198), .A3(new_n199), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n367), .A2(new_n330), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n321), .B1(new_n371), .B2(new_n358), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n363), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT6), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n374), .B(new_n322), .C1(new_n340), .C2(new_n356), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT83), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n362), .B1(new_n373), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n229), .A2(G125), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n379), .B1(new_n239), .B2(G125), .ZN(new_n380));
  INV_X1    g194(.A(G224), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(G953), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n380), .B(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n378), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(G210), .B1(G237), .B2(G902), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(KEYINPUT88), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT7), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT87), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n389), .B1(new_n382), .B2(new_n390), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n380), .B(new_n391), .C1(new_n390), .C2(new_n382), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n382), .B1(KEYINPUT86), .B2(new_n389), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n393), .B1(KEYINPUT86), .B2(new_n389), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n379), .B(new_n394), .C1(new_n239), .C2(G125), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n392), .A2(new_n361), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n355), .A2(new_n344), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n321), .B(KEYINPUT8), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT84), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n349), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n348), .A2(KEYINPUT84), .A3(KEYINPUT5), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n353), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n354), .A2(new_n348), .ZN(new_n404));
  AOI21_X1  g218(.A(KEYINPUT85), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n405), .A2(new_n344), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n403), .A2(KEYINPUT85), .A3(new_n404), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n399), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n291), .B1(new_n396), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n385), .A2(new_n388), .A3(new_n410), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n376), .B(new_n375), .C1(new_n363), .C2(new_n372), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n383), .B1(new_n412), .B2(new_n362), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n387), .B1(new_n413), .B2(new_n409), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(G214), .B1(G237), .B2(G902), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT9), .B(G234), .ZN(new_n418));
  INV_X1    g232(.A(G217), .ZN(new_n419));
  NOR3_X1   g233(.A1(new_n418), .A2(new_n419), .A3(G953), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT91), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n231), .B2(G143), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n221), .A2(KEYINPUT91), .A3(G128), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n231), .A2(G143), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n207), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G122), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G116), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n195), .A2(G122), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n326), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n429), .A2(new_n430), .A3(G107), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n427), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT13), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n425), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n423), .A2(KEYINPUT13), .A3(new_n424), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(new_n437), .A3(new_n426), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n434), .B1(G134), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n429), .A2(KEYINPUT14), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n431), .A2(new_n440), .A3(G107), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n429), .B(new_n430), .C1(KEYINPUT14), .C2(new_n326), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n425), .A2(new_n426), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G134), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n443), .B1(new_n445), .B2(new_n427), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n439), .A2(new_n446), .A3(KEYINPUT92), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT92), .ZN(new_n448));
  INV_X1    g262(.A(new_n434), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n438), .A2(G134), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n445), .A2(new_n427), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(new_n442), .A3(new_n441), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n448), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n421), .B1(new_n447), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT92), .B1(new_n439), .B2(new_n446), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n451), .A2(new_n453), .A3(new_n448), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n457), .A3(new_n420), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n455), .A2(new_n291), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT93), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT93), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n455), .A2(new_n461), .A3(new_n291), .A4(new_n458), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT15), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(G478), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  XOR2_X1   g280(.A(KEYINPUT90), .B(G475), .Z(new_n467));
  INV_X1    g281(.A(G140), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(G125), .ZN(new_n469));
  INV_X1    g283(.A(G125), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(G140), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT75), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT75), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n469), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n473), .A2(new_n475), .A3(new_n219), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n470), .A2(KEYINPUT74), .A3(G140), .ZN(new_n477));
  OAI211_X1 g291(.A(G146), .B(new_n477), .C1(new_n472), .C2(KEYINPUT74), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n187), .A2(G214), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n221), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT18), .ZN(new_n483));
  INV_X1    g297(.A(G131), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n481), .B(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n482), .ZN(new_n486));
  AOI21_X1  g300(.A(G143), .B1(new_n187), .B2(G214), .ZN(new_n487));
  OAI211_X1 g301(.A(KEYINPUT18), .B(G131), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n479), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n481), .A2(new_n482), .ZN(new_n491));
  INV_X1    g305(.A(new_n205), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT17), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n481), .A2(new_n205), .A3(new_n482), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  OAI211_X1 g310(.A(KEYINPUT16), .B(new_n477), .C1(new_n472), .C2(KEYINPUT74), .ZN(new_n497));
  AOI21_X1  g311(.A(KEYINPUT16), .B1(new_n468), .B2(G125), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(G146), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n497), .A2(new_n219), .A3(new_n499), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n491), .A2(KEYINPUT17), .A3(new_n492), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n496), .A2(new_n501), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n490), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(G113), .B(G122), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(new_n323), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n490), .A2(new_n507), .A3(new_n504), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n467), .B1(new_n511), .B2(new_n291), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT20), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT19), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n473), .A2(new_n475), .A3(new_n514), .ZN(new_n515));
  OAI211_X1 g329(.A(KEYINPUT19), .B(new_n477), .C1(new_n472), .C2(KEYINPUT74), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n219), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT89), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT89), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n515), .A2(new_n519), .A3(new_n219), .A4(new_n516), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n500), .A2(G146), .B1(new_n493), .B2(new_n495), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n489), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n510), .B1(new_n523), .B2(new_n507), .ZN(new_n524));
  NOR2_X1   g338(.A1(G475), .A2(G902), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n513), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n524), .A2(new_n513), .A3(new_n525), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n512), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n462), .A2(new_n464), .A3(G478), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(G953), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(G952), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n533), .B1(G234), .B2(G237), .ZN(new_n534));
  AOI211_X1 g348(.A(new_n291), .B(new_n532), .C1(G234), .C2(G237), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT21), .B(G898), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n466), .A2(new_n529), .A3(new_n531), .A4(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n417), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n501), .A2(new_n502), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT23), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n193), .B2(G128), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n231), .A2(KEYINPUT23), .A3(G119), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n543), .B(new_n544), .C1(G119), .C2(new_n231), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(G110), .ZN(new_n546));
  XOR2_X1   g360(.A(KEYINPUT24), .B(G110), .Z(new_n547));
  XNOR2_X1  g361(.A(G119), .B(G128), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(KEYINPUT73), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n541), .A2(new_n546), .A3(new_n550), .ZN(new_n551));
  OAI22_X1  g365(.A1(new_n545), .A2(G110), .B1(new_n548), .B2(new_n547), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n501), .A2(new_n476), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT22), .B(G137), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n532), .A2(G221), .A3(G234), .ZN(new_n556));
  XOR2_X1   g370(.A(new_n555), .B(new_n556), .Z(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n551), .A2(new_n553), .A3(new_n557), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n291), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT25), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n559), .A2(KEYINPUT25), .A3(new_n291), .A4(new_n560), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n419), .B1(G234), .B2(new_n291), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n559), .A2(new_n560), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n566), .A2(G902), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(G221), .ZN(new_n573));
  INV_X1    g387(.A(new_n418), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n573), .B1(new_n574), .B2(new_n291), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n251), .A2(new_n345), .A3(new_n347), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT10), .ZN(new_n577));
  AOI22_X1  g391(.A1(new_n234), .A2(G128), .B1(new_n220), .B2(new_n222), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(new_n233), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT79), .B1(new_n579), .B2(new_n344), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n231), .B1(new_n220), .B2(KEYINPUT1), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n250), .B1(new_n226), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT79), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n582), .A2(new_n583), .A3(new_n337), .A4(new_n343), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT10), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n580), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n577), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT78), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n229), .A2(new_n331), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n588), .B1(new_n360), .B2(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n366), .A2(KEYINPUT78), .A3(new_n229), .A4(new_n331), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n587), .A2(new_n271), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n532), .A2(G227), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(KEYINPUT76), .ZN(new_n594));
  XNOR2_X1  g408(.A(G110), .B(G140), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT82), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT82), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n592), .A2(new_n599), .A3(new_n596), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT81), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n580), .A2(new_n584), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n239), .A2(new_n344), .ZN(new_n603));
  OAI211_X1 g417(.A(KEYINPUT12), .B(new_n218), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT12), .ZN(new_n605));
  AOI22_X1  g419(.A1(new_n580), .A2(new_n584), .B1(new_n239), .B2(new_n344), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n605), .B1(new_n606), .B2(new_n271), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n601), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n604), .A2(new_n607), .A3(new_n601), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n598), .A2(new_n600), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n587), .A2(new_n590), .A3(new_n591), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n218), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n596), .B1(new_n613), .B2(new_n592), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(G469), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n616), .A2(new_n617), .A3(new_n291), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n604), .A2(new_n607), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n592), .ZN(new_n620));
  INV_X1    g434(.A(new_n596), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n613), .A2(new_n592), .A3(new_n596), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n617), .B1(new_n624), .B2(new_n291), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n575), .B1(new_n618), .B2(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n320), .A2(new_n540), .A3(new_n572), .A4(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G101), .ZN(G3));
  AND2_X1   g443(.A1(new_n304), .A2(new_n306), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n312), .A2(new_n313), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n294), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(G902), .B1(new_n299), .B2(new_n307), .ZN(new_n633));
  INV_X1    g447(.A(G472), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(new_n571), .ZN(new_n636));
  INV_X1    g450(.A(new_n386), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n385), .A2(new_n637), .A3(new_n410), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n386), .B1(new_n413), .B2(new_n409), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n638), .A2(new_n639), .A3(new_n416), .A4(new_n538), .ZN(new_n640));
  INV_X1    g454(.A(new_n458), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n420), .B1(new_n456), .B2(new_n457), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT94), .ZN(new_n643));
  OAI22_X1  g457(.A1(new_n641), .A2(new_n642), .B1(new_n643), .B2(KEYINPUT33), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT94), .B(KEYINPUT33), .Z(new_n645));
  NAND3_X1  g459(.A1(new_n455), .A2(new_n458), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(G478), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n647), .A2(G902), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n644), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n459), .A2(new_n647), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n510), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n507), .B1(new_n490), .B2(new_n504), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n291), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n467), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n528), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n656), .B1(new_n657), .B2(new_n526), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n651), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(KEYINPUT95), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT95), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n651), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n640), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n636), .A2(new_n663), .A3(new_n627), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT34), .B(G104), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G6));
  NOR2_X1   g480(.A1(new_n656), .A2(KEYINPUT96), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT96), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n512), .A2(new_n668), .ZN(new_n669));
  OAI22_X1  g483(.A1(new_n667), .A2(new_n669), .B1(new_n526), .B2(new_n657), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n530), .B1(new_n465), .B2(new_n463), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n640), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n636), .A2(new_n672), .A3(new_n627), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT35), .B(G107), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G9));
  INV_X1    g489(.A(new_n635), .ZN(new_n676));
  OR2_X1    g490(.A1(new_n558), .A2(KEYINPUT36), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n554), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n554), .A2(new_n677), .ZN(new_n679));
  NOR4_X1   g493(.A1(new_n678), .A2(new_n679), .A3(G902), .A4(new_n566), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n680), .B1(new_n565), .B2(new_n566), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n540), .A2(new_n676), .A3(new_n627), .A4(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT37), .B(G110), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G12));
  NAND3_X1  g499(.A1(new_n638), .A2(new_n416), .A3(new_n639), .ZN(new_n686));
  INV_X1    g500(.A(G900), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n535), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n534), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NOR4_X1   g505(.A1(new_n670), .A2(new_n686), .A3(new_n671), .A4(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n692), .A2(new_n320), .A3(new_n627), .A4(new_n682), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G128), .ZN(G30));
  XNOR2_X1  g508(.A(new_n690), .B(KEYINPUT39), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n627), .A2(new_n695), .ZN(new_n696));
  OR2_X1    g510(.A1(new_n696), .A2(KEYINPUT40), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n415), .B(KEYINPUT38), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n671), .A2(new_n529), .ZN(new_n699));
  AND4_X1   g513(.A1(new_n416), .A2(new_n698), .A3(new_n681), .A4(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n696), .A2(KEYINPUT40), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n315), .A2(new_n262), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n191), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  AND2_X1   g518(.A1(new_n286), .A2(new_n288), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n291), .B1(new_n705), .B2(new_n191), .ZN(new_n706));
  OAI21_X1  g520(.A(G472), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n707), .B1(new_n308), .B2(new_n319), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n697), .A2(new_n700), .A3(new_n701), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G143), .ZN(G45));
  INV_X1    g524(.A(KEYINPUT97), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n651), .A2(new_n658), .A3(new_n690), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n638), .A2(new_n416), .A3(new_n639), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n651), .A2(new_n658), .A3(new_n690), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n715), .A2(new_n686), .A3(KEYINPUT97), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n320), .A2(new_n627), .A3(new_n682), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(new_n219), .ZN(G48));
  AOI21_X1  g535(.A(new_n617), .B1(new_n616), .B2(new_n291), .ZN(new_n722));
  AOI211_X1 g536(.A(G469), .B(G902), .C1(new_n611), .C2(new_n615), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n722), .A2(new_n723), .A3(new_n575), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n724), .A2(new_n663), .A3(new_n320), .A4(new_n572), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT41), .B(G113), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G15));
  NAND4_X1  g541(.A1(new_n724), .A2(new_n320), .A3(new_n572), .A4(new_n672), .ZN(new_n728));
  XNOR2_X1  g542(.A(KEYINPUT98), .B(G116), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(G18));
  AOI21_X1  g544(.A(new_n599), .B1(new_n592), .B2(new_n596), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n604), .A2(new_n607), .A3(new_n601), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n731), .A2(new_n732), .A3(new_n608), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n614), .B1(new_n733), .B2(new_n600), .ZN(new_n734));
  OAI21_X1  g548(.A(G469), .B1(new_n734), .B2(G902), .ZN(new_n735));
  INV_X1    g549(.A(new_n575), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n735), .A2(new_n713), .A3(new_n736), .A4(new_n618), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n539), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n738), .A2(new_n320), .A3(new_n739), .A4(new_n682), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G119), .ZN(G21));
  AOI21_X1  g555(.A(new_n634), .B1(new_n318), .B2(new_n291), .ZN(new_n742));
  XOR2_X1   g556(.A(new_n294), .B(KEYINPUT99), .Z(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n289), .A2(new_n274), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n192), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n744), .B1(new_n746), .B2(new_n307), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n742), .A2(new_n571), .A3(new_n747), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n686), .A2(new_n671), .A3(new_n529), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n724), .A2(new_n748), .A3(new_n538), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G122), .ZN(G24));
  NOR4_X1   g565(.A1(new_n742), .A2(new_n715), .A3(new_n747), .A4(new_n681), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n738), .A2(new_n752), .A3(KEYINPUT100), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT100), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n318), .A2(new_n291), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(G472), .ZN(new_n756));
  INV_X1    g570(.A(new_n747), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n756), .A2(new_n682), .A3(new_n712), .A4(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n754), .B1(new_n758), .B2(new_n737), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n753), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G125), .ZN(G27));
  NAND3_X1  g575(.A1(new_n411), .A2(new_n416), .A3(new_n414), .ZN(new_n762));
  AOI211_X1 g576(.A(new_n575), .B(new_n762), .C1(new_n618), .C2(new_n626), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n763), .A2(new_n320), .A3(new_n572), .A4(new_n712), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT42), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n632), .A2(KEYINPUT32), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n295), .B1(new_n299), .B2(new_n307), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n309), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n291), .B(new_n290), .C1(new_n279), .C2(new_n283), .ZN(new_n770));
  AOI22_X1  g584(.A1(new_n767), .A2(new_n769), .B1(G472), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(new_n571), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n772), .A2(KEYINPUT42), .A3(new_n712), .A4(new_n763), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n766), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G131), .ZN(G33));
  NOR3_X1   g589(.A1(new_n670), .A2(new_n671), .A3(new_n691), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n763), .A2(new_n320), .A3(new_n572), .A4(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  NOR2_X1   g592(.A1(new_n617), .A2(new_n291), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n617), .B1(new_n624), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n622), .A2(new_n623), .A3(KEYINPUT45), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n779), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n618), .B1(new_n783), .B2(KEYINPUT46), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n590), .A2(new_n591), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n271), .B1(new_n785), .B2(new_n587), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n597), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n596), .B1(new_n619), .B2(new_n592), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n780), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(G469), .A3(new_n782), .ZN(new_n790));
  INV_X1    g604(.A(new_n779), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n790), .A2(KEYINPUT46), .A3(new_n791), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n736), .B(new_n695), .C1(new_n784), .C2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT44), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT102), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n658), .A2(new_n795), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n656), .B(KEYINPUT102), .C1(new_n657), .C2(new_n526), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT43), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n798), .B1(new_n649), .B2(new_n650), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n796), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  XOR2_X1   g614(.A(KEYINPUT101), .B(KEYINPUT43), .Z(new_n801));
  AND2_X1   g615(.A1(new_n649), .A2(new_n650), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n801), .B1(new_n802), .B2(new_n658), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n635), .A3(new_n682), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n793), .B1(new_n794), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n804), .A2(KEYINPUT44), .A3(new_n635), .A4(new_n682), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n411), .A2(new_n416), .A3(new_n414), .ZN(new_n808));
  AOI21_X1  g622(.A(KEYINPUT103), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n807), .A2(KEYINPUT103), .A3(new_n808), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n806), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G137), .ZN(G39));
  NOR4_X1   g627(.A1(new_n320), .A2(new_n572), .A3(new_n715), .A4(new_n762), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n790), .A2(new_n791), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT46), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n723), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n783), .A2(KEYINPUT46), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n575), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n820), .ZN(new_n822));
  AOI211_X1 g636(.A(new_n575), .B(new_n822), .C1(new_n817), .C2(new_n818), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n814), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(KEYINPUT105), .B(G140), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n824), .B(new_n825), .ZN(G42));
  AOI21_X1  g640(.A(KEYINPUT112), .B1(new_n724), .B2(new_n808), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n689), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n724), .A2(KEYINPUT112), .A3(new_n808), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n828), .A2(new_n772), .A3(new_n804), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT114), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n830), .A2(KEYINPUT114), .ZN(new_n833));
  OAI211_X1 g647(.A(KEYINPUT115), .B(KEYINPUT48), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n833), .ZN(new_n835));
  XOR2_X1   g649(.A(KEYINPUT115), .B(KEYINPUT48), .Z(new_n836));
  NAND3_X1  g650(.A1(new_n835), .A2(new_n831), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n660), .A2(new_n662), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n708), .A2(new_n571), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n828), .A2(new_n838), .A3(new_n829), .A4(new_n839), .ZN(new_n840));
  XOR2_X1   g654(.A(new_n533), .B(KEYINPUT113), .Z(new_n841));
  AOI21_X1  g655(.A(new_n689), .B1(new_n800), .B2(new_n803), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n748), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n841), .B1(new_n844), .B2(new_n738), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n834), .A2(new_n837), .A3(new_n840), .A4(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n724), .ZN(new_n847));
  NOR4_X1   g661(.A1(new_n843), .A2(new_n847), .A3(new_n698), .A4(new_n416), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(KEYINPUT50), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n736), .B1(new_n784), .B2(new_n792), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(new_n822), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n819), .A2(new_n820), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n722), .A2(new_n723), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT111), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n736), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n855), .B1(new_n854), .B2(new_n853), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n851), .A2(new_n852), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(new_n808), .A3(new_n844), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n742), .A2(new_n681), .A3(new_n747), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n828), .A2(new_n859), .A3(new_n804), .A4(new_n829), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n651), .A2(new_n658), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n828), .A2(new_n829), .A3(new_n839), .A4(new_n861), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n849), .A2(new_n858), .A3(new_n860), .A4(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT51), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n864), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n846), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n868));
  AND4_X1   g682(.A1(new_n725), .A2(new_n740), .A3(new_n728), .A4(new_n750), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n774), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n659), .B1(new_n671), .B2(new_n658), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n417), .A2(new_n537), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n636), .A2(new_n627), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n873), .A2(new_n628), .A3(new_n683), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT107), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n763), .A2(new_n752), .A3(new_n876), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n808), .B(new_n736), .C1(new_n723), .C2(new_n625), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT107), .B1(new_n758), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n466), .A2(new_n531), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n670), .A2(new_n881), .A3(new_n691), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n763), .A2(new_n320), .A3(new_n682), .A4(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n875), .A2(new_n777), .A3(new_n880), .A4(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n870), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n719), .ZN(new_n886));
  AND4_X1   g700(.A1(new_n627), .A2(new_n749), .A3(new_n681), .A4(new_n690), .ZN(new_n887));
  AOI22_X1  g701(.A1(new_n886), .A2(new_n717), .B1(new_n887), .B2(new_n708), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n888), .A2(KEYINPUT52), .A3(new_n693), .A4(new_n760), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT52), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT100), .B1(new_n738), .B2(new_n752), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n758), .A2(new_n737), .A3(new_n754), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n693), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n682), .A2(new_n691), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n708), .A2(new_n627), .A3(new_n749), .A4(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n895), .B1(new_n718), .B2(new_n719), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n890), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n889), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n868), .B1(new_n885), .B2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n893), .A2(KEYINPUT108), .ZN(new_n901));
  INV_X1    g715(.A(new_n720), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT108), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n760), .A2(new_n903), .A3(new_n693), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n895), .A2(KEYINPUT52), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n897), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n907), .A2(new_n868), .A3(new_n885), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n900), .A2(new_n908), .A3(KEYINPUT54), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT109), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT110), .B1(new_n869), .B2(new_n774), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n912), .A2(new_n868), .A3(new_n884), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n869), .A2(KEYINPUT110), .A3(new_n774), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n913), .A2(new_n907), .A3(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT54), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n885), .A2(new_n898), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n868), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n900), .A2(new_n908), .A3(KEYINPUT109), .A4(KEYINPUT54), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n867), .A2(new_n911), .A3(new_n919), .A4(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n921), .B1(G952), .B2(G953), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n853), .B(KEYINPUT49), .Z(new_n923));
  NAND4_X1  g737(.A1(new_n572), .A2(new_n736), .A3(new_n416), .A4(new_n651), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n796), .A2(new_n797), .ZN(new_n925));
  OR3_X1    g739(.A1(new_n698), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n923), .A2(new_n926), .A3(new_n708), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT106), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n922), .A2(new_n928), .ZN(G75));
  INV_X1    g743(.A(KEYINPUT56), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n915), .A2(new_n918), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(G902), .ZN(new_n932));
  INV_X1    g746(.A(G210), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n378), .B(KEYINPUT116), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT117), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT55), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(new_n383), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n938), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n930), .B(new_n940), .C1(new_n932), .C2(new_n933), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n532), .A2(G952), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n939), .A2(new_n941), .A3(new_n943), .ZN(G51));
  AOI21_X1  g758(.A(new_n291), .B1(new_n915), .B2(new_n918), .ZN(new_n945));
  INV_X1    g759(.A(new_n790), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n945), .A2(KEYINPUT118), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(KEYINPUT118), .B1(new_n945), .B2(new_n946), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n779), .B(KEYINPUT57), .ZN(new_n950));
  INV_X1    g764(.A(new_n919), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n916), .B1(new_n915), .B2(new_n918), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n616), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n942), .B1(new_n949), .B2(new_n954), .ZN(G54));
  AND2_X1   g769(.A1(KEYINPUT58), .A2(G475), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n945), .A2(new_n524), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n524), .B1(new_n945), .B2(new_n956), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n957), .A2(new_n958), .A3(new_n942), .ZN(G60));
  NAND2_X1  g773(.A1(new_n644), .A2(new_n646), .ZN(new_n960));
  NAND2_X1  g774(.A1(G478), .A2(G902), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT59), .Z(new_n962));
  NOR2_X1   g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n963), .B1(new_n951), .B2(new_n952), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n943), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n911), .A2(new_n919), .A3(new_n920), .ZN(new_n966));
  INV_X1    g780(.A(new_n962), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n965), .B1(new_n968), .B2(new_n960), .ZN(G63));
  NAND2_X1  g783(.A1(KEYINPUT119), .A2(KEYINPUT61), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT120), .Z(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(G217), .A2(G902), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT60), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n974), .B1(new_n915), .B2(new_n918), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n678), .A2(new_n679), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(KEYINPUT119), .A2(KEYINPUT61), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n942), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n975), .B2(new_n568), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n972), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  OR2_X1    g796(.A1(new_n975), .A2(new_n568), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n983), .A2(new_n971), .A3(new_n977), .A4(new_n980), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n982), .A2(new_n984), .ZN(G66));
  OAI21_X1  g799(.A(G953), .B1(new_n536), .B2(new_n381), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n869), .A2(new_n875), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n986), .B1(new_n988), .B2(G953), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n935), .B1(G898), .B2(new_n532), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n989), .B(new_n990), .ZN(G69));
  NAND2_X1  g805(.A1(new_n515), .A2(new_n516), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n303), .B(new_n992), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT121), .Z(new_n994));
  NAND3_X1  g808(.A1(new_n772), .A2(new_n808), .A3(new_n871), .ZN(new_n995));
  OR2_X1    g809(.A1(new_n995), .A2(new_n696), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n812), .A2(new_n824), .A3(new_n996), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n901), .A2(new_n709), .A3(new_n902), .A4(new_n904), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT62), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n720), .B1(new_n893), .B2(KEYINPUT108), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n1001), .A2(KEYINPUT62), .A3(new_n709), .A4(new_n904), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n997), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n994), .B1(new_n1003), .B2(G953), .ZN(new_n1004));
  INV_X1    g818(.A(new_n777), .ZN(new_n1005));
  AOI211_X1 g819(.A(KEYINPUT123), .B(new_n1005), .C1(new_n766), .C2(new_n773), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT123), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1007), .B1(new_n774), .B2(new_n777), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n320), .A2(new_n572), .A3(new_n749), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n793), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n851), .A2(new_n852), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1011), .B1(new_n1012), .B2(new_n814), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n1001), .A2(new_n1013), .A3(new_n812), .A4(new_n904), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n532), .B1(new_n1009), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT124), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n532), .A2(G900), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1017), .B(KEYINPUT122), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1015), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(new_n993), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1016), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1004), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n532), .B1(G227), .B2(G900), .ZN(new_n1023));
  INV_X1    g837(.A(KEYINPUT125), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OR2_X1    g839(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1022), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1021), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1028), .A2(new_n993), .A3(new_n1019), .ZN(new_n1029));
  NAND4_X1  g843(.A1(new_n1029), .A2(new_n1024), .A3(new_n1023), .A4(new_n1004), .ZN(new_n1030));
  AND2_X1   g844(.A1(new_n1027), .A2(new_n1030), .ZN(G72));
  AND2_X1   g845(.A1(new_n877), .A2(new_n879), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n777), .A2(new_n883), .ZN(new_n1033));
  NOR3_X1   g847(.A1(new_n1032), .A2(new_n1033), .A3(new_n874), .ZN(new_n1034));
  NAND4_X1  g848(.A1(new_n1034), .A2(new_n868), .A3(new_n774), .A4(new_n869), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n1001), .A2(KEYINPUT52), .A3(new_n895), .A4(new_n904), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1035), .B1(new_n897), .B2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g851(.A1(new_n702), .A2(new_n191), .ZN(new_n1038));
  INV_X1    g852(.A(new_n1038), .ZN(new_n1039));
  NAND2_X1  g853(.A1(G472), .A2(G902), .ZN(new_n1040));
  XOR2_X1   g854(.A(new_n1040), .B(KEYINPUT63), .Z(new_n1041));
  NAND3_X1  g855(.A1(new_n1039), .A2(new_n703), .A3(new_n1041), .ZN(new_n1042));
  NOR3_X1   g856(.A1(new_n1037), .A2(new_n899), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1044));
  INV_X1    g858(.A(new_n997), .ZN(new_n1045));
  NAND3_X1  g859(.A1(new_n1044), .A2(new_n988), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1046), .A2(new_n1041), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n1043), .B1(new_n1047), .B2(new_n704), .ZN(new_n1048));
  NOR3_X1   g862(.A1(new_n1009), .A2(new_n1014), .A3(new_n987), .ZN(new_n1049));
  INV_X1    g863(.A(new_n1041), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n1038), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g865(.A(KEYINPUT126), .B1(new_n1051), .B2(new_n943), .ZN(new_n1052));
  NOR3_X1   g866(.A1(new_n771), .A2(new_n878), .A3(new_n571), .ZN(new_n1053));
  AOI21_X1  g867(.A(KEYINPUT42), .B1(new_n1053), .B2(new_n712), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n320), .A2(new_n572), .ZN(new_n1055));
  NOR4_X1   g869(.A1(new_n1055), .A2(new_n765), .A3(new_n715), .A4(new_n878), .ZN(new_n1056));
  OAI21_X1  g870(.A(new_n777), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n1057), .A2(KEYINPUT123), .ZN(new_n1058));
  NAND3_X1  g872(.A1(new_n774), .A2(new_n1007), .A3(new_n777), .ZN(new_n1059));
  NAND2_X1  g873(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  AND3_X1   g874(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(new_n1061));
  INV_X1    g875(.A(new_n1011), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n824), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g877(.A1(new_n805), .A2(new_n794), .ZN(new_n1064));
  NAND3_X1  g878(.A1(new_n1064), .A2(new_n695), .A3(new_n819), .ZN(new_n1065));
  AND3_X1   g879(.A1(new_n807), .A2(KEYINPUT103), .A3(new_n808), .ZN(new_n1066));
  NOR3_X1   g880(.A1(new_n1065), .A2(new_n1066), .A3(new_n809), .ZN(new_n1067));
  NOR2_X1   g881(.A1(new_n1063), .A2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g882(.A1(new_n1060), .A2(new_n1061), .A3(new_n988), .A4(new_n1068), .ZN(new_n1069));
  AOI21_X1  g883(.A(new_n1039), .B1(new_n1069), .B2(new_n1041), .ZN(new_n1070));
  INV_X1    g884(.A(KEYINPUT126), .ZN(new_n1071));
  NOR3_X1   g885(.A1(new_n1070), .A2(new_n1071), .A3(new_n942), .ZN(new_n1072));
  OAI21_X1  g886(.A(new_n1048), .B1(new_n1052), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g887(.A1(new_n1073), .A2(KEYINPUT127), .ZN(new_n1074));
  INV_X1    g888(.A(KEYINPUT127), .ZN(new_n1075));
  OAI211_X1 g889(.A(new_n1048), .B(new_n1075), .C1(new_n1052), .C2(new_n1072), .ZN(new_n1076));
  NAND2_X1  g890(.A1(new_n1074), .A2(new_n1076), .ZN(G57));
endmodule


