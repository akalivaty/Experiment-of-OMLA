//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 0 0 0 1 0 0 1 1 0 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n837, new_n838, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n971, new_n972;
  XNOR2_X1  g000(.A(KEYINPUT80), .B(KEYINPUT6), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g002(.A1(G225gat), .A2(G233gat), .ZN(new_n204));
  INV_X1    g003(.A(G134gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G127gat), .ZN(new_n206));
  INV_X1    g005(.A(G127gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G134gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n206), .A2(new_n208), .A3(KEYINPUT67), .ZN(new_n209));
  OR3_X1    g008(.A1(new_n207), .A2(KEYINPUT67), .A3(G134gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(G113gat), .B(G120gat), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n209), .B(new_n210), .C1(KEYINPUT1), .C2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G120gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G113gat), .ZN(new_n214));
  INV_X1    g013(.A(G113gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G120gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT68), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n214), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT1), .ZN(new_n219));
  XNOR2_X1  g018(.A(G127gat), .B(G134gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n215), .A2(KEYINPUT68), .A3(G120gat), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223));
  INV_X1    g022(.A(G155gat), .ZN(new_n224));
  INV_X1    g023(.A(G162gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G141gat), .B(G148gat), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n223), .B(new_n226), .C1(new_n227), .C2(KEYINPUT2), .ZN(new_n228));
  INV_X1    g027(.A(G141gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G148gat), .ZN(new_n230));
  INV_X1    g029(.A(G148gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G141gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n226), .A2(new_n223), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n223), .A2(KEYINPUT2), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n212), .A2(new_n222), .A3(new_n228), .A4(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT4), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n209), .A2(new_n210), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT1), .B1(new_n214), .B2(new_n216), .ZN(new_n242));
  AND3_X1   g041(.A1(new_n214), .A2(new_n216), .A3(new_n217), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n221), .A2(new_n206), .A3(new_n208), .A4(new_n219), .ZN(new_n244));
  OAI22_X1  g043(.A1(new_n241), .A2(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT76), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT76), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n212), .A2(new_n222), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n228), .A2(new_n249), .A3(new_n236), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n234), .B1(new_n235), .B2(new_n233), .ZN(new_n252));
  OAI21_X1  g051(.A(KEYINPUT3), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n246), .A2(new_n248), .A3(new_n250), .A4(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n254), .A2(KEYINPUT77), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT77), .ZN(new_n256));
  AND3_X1   g055(.A1(new_n212), .A2(new_n247), .A3(new_n222), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n247), .B1(new_n212), .B2(new_n222), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n228), .A2(new_n249), .A3(new_n236), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n249), .B1(new_n228), .B2(new_n236), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n256), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n204), .B(new_n240), .C1(new_n255), .C2(new_n263), .ZN(new_n264));
  XOR2_X1   g063(.A(KEYINPUT78), .B(KEYINPUT5), .Z(new_n265));
  NAND2_X1  g064(.A1(new_n228), .A2(new_n236), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n246), .A2(new_n248), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(new_n237), .ZN(new_n268));
  INV_X1    g067(.A(new_n204), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n265), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n264), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n254), .A2(KEYINPUT77), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n262), .A2(new_n256), .A3(new_n246), .A4(new_n248), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n239), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n274), .A2(new_n204), .A3(new_n265), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(G1gat), .B(G29gat), .Z(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G57gat), .B(G85gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n203), .B1(new_n276), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n281), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n271), .A2(new_n283), .A3(new_n275), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  AOI211_X1 g084(.A(new_n283), .B(new_n202), .C1(new_n271), .C2(new_n275), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G71gat), .B(G78gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n289), .A2(KEYINPUT92), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(G57gat), .B(G64gat), .ZN(new_n292));
  NOR3_X1   g091(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n289), .A2(KEYINPUT92), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI211_X1 g094(.A(KEYINPUT92), .B(new_n289), .C1(new_n292), .C2(new_n291), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(KEYINPUT21), .ZN(new_n298));
  NAND2_X1  g097(.A1(G231gat), .A2(G233gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n300), .B(new_n207), .ZN(new_n301));
  XNOR2_X1  g100(.A(G183gat), .B(G211gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G15gat), .B(G22gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n304), .B(KEYINPUT86), .ZN(new_n305));
  INV_X1    g104(.A(G1gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(G8gat), .B1(new_n307), .B2(KEYINPUT87), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT86), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n304), .B(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT16), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n310), .B1(new_n311), .B2(G1gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(new_n307), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n308), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n312), .B(new_n307), .C1(KEYINPUT87), .C2(G8gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n297), .A2(KEYINPUT21), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n321), .B(new_n224), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n320), .B(new_n322), .ZN(new_n323));
  OR2_X1    g122(.A1(new_n303), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n303), .A2(new_n323), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G29gat), .ZN(new_n327));
  INV_X1    g126(.A(G36gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n327), .A2(new_n328), .A3(KEYINPUT14), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT14), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n330), .B1(G29gat), .B2(G36gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(KEYINPUT85), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n327), .A2(new_n328), .ZN(new_n334));
  XNOR2_X1  g133(.A(G43gat), .B(G50gat), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n334), .B1(new_n335), .B2(KEYINPUT15), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n336), .B1(KEYINPUT15), .B2(new_n335), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  OAI211_X1 g137(.A(KEYINPUT15), .B(new_n335), .C1(new_n332), .C2(new_n334), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G85gat), .A2(G92gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n341), .B(KEYINPUT7), .ZN(new_n342));
  NAND2_X1  g141(.A1(G99gat), .A2(G106gat), .ZN(new_n343));
  INV_X1    g142(.A(G85gat), .ZN(new_n344));
  INV_X1    g143(.A(G92gat), .ZN(new_n345));
  AOI22_X1  g144(.A1(KEYINPUT8), .A2(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  XOR2_X1   g146(.A(G99gat), .B(G106gat), .Z(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n347), .B(new_n349), .ZN(new_n350));
  AND2_X1   g149(.A1(G232gat), .A2(G233gat), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n340), .A2(new_n350), .B1(KEYINPUT41), .B2(new_n351), .ZN(new_n352));
  XOR2_X1   g151(.A(new_n350), .B(KEYINPUT95), .Z(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT17), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n340), .B(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n352), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  XOR2_X1   g156(.A(G190gat), .B(G218gat), .Z(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n358), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n360), .B(new_n352), .C1(new_n356), .C2(new_n354), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n351), .A2(KEYINPUT41), .ZN(new_n363));
  XNOR2_X1  g162(.A(G134gat), .B(G162gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n359), .A2(new_n361), .A3(new_n365), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  XOR2_X1   g169(.A(G120gat), .B(G148gat), .Z(new_n371));
  XNOR2_X1  g170(.A(new_n371), .B(KEYINPUT97), .ZN(new_n372));
  XNOR2_X1  g171(.A(G176gat), .B(G204gat), .ZN(new_n373));
  XOR2_X1   g172(.A(new_n372), .B(new_n373), .Z(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(G230gat), .A2(G233gat), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  OR2_X1    g176(.A1(new_n349), .A2(KEYINPUT96), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n297), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n350), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n297), .A2(new_n350), .A3(new_n378), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n297), .A2(KEYINPUT10), .A3(new_n350), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n377), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n376), .B1(new_n381), .B2(new_n383), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT98), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n375), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI211_X1 g189(.A(KEYINPUT98), .B(new_n374), .C1(new_n386), .C2(new_n387), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NOR3_X1   g192(.A1(new_n326), .A2(new_n370), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT72), .ZN(new_n395));
  NAND2_X1  g194(.A1(G211gat), .A2(G218gat), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT22), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G211gat), .B(G218gat), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n398), .B1(new_n400), .B2(KEYINPUT73), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT73), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n396), .A2(new_n395), .A3(new_n397), .ZN(new_n404));
  XNOR2_X1  g203(.A(G197gat), .B(G204gat), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n401), .A2(new_n403), .A3(new_n404), .A4(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n404), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n402), .B(new_n399), .C1(new_n407), .C2(new_n398), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n249), .B1(new_n409), .B2(KEYINPUT29), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n266), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT29), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n250), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G78gat), .B(G106gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n416), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n411), .A2(new_n414), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT81), .B1(new_n409), .B2(new_n413), .ZN(new_n421));
  AND2_X1   g220(.A1(G228gat), .A2(G233gat), .ZN(new_n422));
  OAI21_X1  g221(.A(G22gat), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NOR3_X1   g223(.A1(new_n421), .A2(G22gat), .A3(new_n422), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT31), .B(G50gat), .ZN(new_n426));
  NOR3_X1   g225(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n426), .ZN(new_n428));
  OR3_X1    g227(.A1(new_n421), .A2(G22gat), .A3(new_n422), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n428), .B1(new_n429), .B2(new_n423), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n420), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n426), .B1(new_n424), .B2(new_n425), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n429), .A2(new_n423), .A3(new_n428), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n432), .A2(new_n419), .A3(new_n433), .A4(new_n417), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n240), .B1(new_n255), .B2(new_n263), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT39), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(new_n438), .A3(new_n269), .ZN(new_n439));
  INV_X1    g238(.A(new_n237), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n440), .B1(new_n259), .B2(new_n266), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n438), .B1(new_n441), .B2(new_n204), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n442), .B1(new_n274), .B2(new_n204), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n439), .A2(new_n443), .A3(new_n283), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT40), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n276), .A2(new_n281), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n439), .A2(new_n443), .A3(KEYINPUT40), .A4(new_n283), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n409), .ZN(new_n450));
  NAND2_X1  g249(.A1(G226gat), .A2(G233gat), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NOR2_X1   g251(.A1(G169gat), .A2(G176gat), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT26), .ZN(new_n455));
  NAND2_X1  g254(.A1(G169gat), .A2(G176gat), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AOI22_X1  g256(.A1(new_n453), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  XOR2_X1   g258(.A(KEYINPUT27), .B(G183gat), .Z(new_n460));
  INV_X1    g259(.A(KEYINPUT28), .ZN(new_n461));
  OR3_X1    g260(.A1(new_n460), .A2(new_n461), .A3(G190gat), .ZN(new_n462));
  INV_X1    g261(.A(G190gat), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT27), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n464), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n465));
  AND2_X1   g264(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n463), .B(new_n465), .C1(new_n466), .C2(new_n464), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n461), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n459), .B1(new_n462), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT24), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n471), .A2(G183gat), .A3(G190gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(G183gat), .B(G190gat), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n472), .B1(new_n473), .B2(new_n471), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n456), .A2(KEYINPUT23), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n454), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT64), .ZN(new_n477));
  INV_X1    g276(.A(G169gat), .ZN(new_n478));
  INV_X1    g277(.A(G176gat), .ZN(new_n479));
  AND4_X1   g278(.A1(new_n477), .A2(new_n478), .A3(new_n479), .A4(KEYINPUT23), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n477), .B1(new_n453), .B2(KEYINPUT23), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n476), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n474), .B1(new_n482), .B2(KEYINPUT65), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT65), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n476), .B(new_n484), .C1(new_n480), .C2(new_n481), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT25), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n478), .A2(new_n479), .A3(KEYINPUT23), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n476), .A2(KEYINPUT25), .A3(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n488), .A2(new_n474), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n470), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n452), .B1(new_n490), .B2(new_n412), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT25), .ZN(new_n492));
  INV_X1    g291(.A(new_n472), .ZN(new_n493));
  XOR2_X1   g292(.A(G183gat), .B(G190gat), .Z(new_n494));
  AOI21_X1  g293(.A(new_n493), .B1(new_n494), .B2(KEYINPUT24), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n487), .A2(KEYINPUT64), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n453), .A2(new_n477), .A3(KEYINPUT23), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n496), .A2(new_n497), .B1(new_n454), .B2(new_n475), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n495), .B1(new_n498), .B2(new_n484), .ZN(new_n499));
  INV_X1    g298(.A(new_n485), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n492), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n489), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n469), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n503), .A2(new_n451), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n450), .B1(new_n491), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n451), .B1(new_n503), .B2(KEYINPUT29), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n452), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n506), .A2(new_n409), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  XOR2_X1   g308(.A(G8gat), .B(G36gat), .Z(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT74), .ZN(new_n511));
  XNOR2_X1  g310(.A(G64gat), .B(G92gat), .ZN(new_n512));
  XOR2_X1   g311(.A(new_n511), .B(new_n512), .Z(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n509), .A2(KEYINPUT30), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n505), .A2(new_n508), .A3(new_n513), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n513), .B1(new_n505), .B2(new_n508), .ZN(new_n517));
  XOR2_X1   g316(.A(KEYINPUT75), .B(KEYINPUT30), .Z(new_n518));
  OAI211_X1 g317(.A(new_n515), .B(new_n516), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n436), .B1(new_n449), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n286), .B1(new_n282), .B2(new_n284), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT37), .ZN(new_n522));
  NOR3_X1   g321(.A1(new_n491), .A2(new_n504), .A3(new_n450), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n409), .B1(new_n506), .B2(new_n507), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n505), .A2(new_n508), .A3(KEYINPUT37), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(new_n513), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT38), .ZN(new_n528));
  INV_X1    g327(.A(new_n517), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n521), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT38), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n525), .A2(new_n531), .A3(new_n513), .A4(new_n526), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT82), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n514), .B1(new_n509), .B2(new_n522), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n535), .A2(KEYINPUT82), .A3(new_n531), .A4(new_n526), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n520), .B1(new_n530), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT70), .ZN(new_n539));
  INV_X1    g338(.A(new_n245), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n482), .A2(KEYINPUT65), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n541), .A2(new_n485), .A3(new_n495), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n489), .B1(new_n542), .B2(new_n492), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n540), .B1(new_n543), .B2(new_n469), .ZN(new_n544));
  NAND2_X1  g343(.A1(G227gat), .A2(G233gat), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n470), .B(new_n245), .C1(new_n486), .C2(new_n489), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT32), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT33), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(G15gat), .B(G43gat), .Z(new_n552));
  XNOR2_X1  g351(.A(G71gat), .B(G99gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n549), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n554), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n548), .B(KEYINPUT32), .C1(new_n550), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n544), .A2(new_n547), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT34), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n559), .A2(new_n560), .A3(new_n545), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT69), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n546), .B1(new_n544), .B2(new_n547), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n564), .A2(KEYINPUT69), .A3(new_n560), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n559), .A2(new_n545), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT34), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n563), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n558), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT69), .B1(new_n564), .B2(new_n560), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n564), .A2(new_n560), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n572), .A2(new_n565), .B1(new_n555), .B2(new_n557), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n539), .B1(new_n569), .B2(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n572), .A2(new_n555), .A3(new_n557), .A4(new_n565), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n568), .ZN(new_n576));
  AOI21_X1  g375(.A(KEYINPUT71), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n574), .B(KEYINPUT36), .C1(new_n577), .C2(new_n539), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(new_n576), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT71), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT36), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(KEYINPUT70), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n515), .A2(new_n516), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n517), .A2(new_n518), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n288), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(new_n436), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n538), .A2(new_n578), .A3(new_n583), .A4(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n575), .A2(new_n576), .A3(new_n435), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT35), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n521), .A2(new_n519), .ZN(new_n592));
  INV_X1    g391(.A(new_n579), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT35), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n592), .A2(new_n593), .A3(new_n594), .A4(new_n435), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n589), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT83), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT83), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n589), .A2(new_n599), .A3(new_n596), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT90), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n314), .A2(new_n315), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(new_n340), .ZN(new_n604));
  NAND2_X1  g403(.A1(G229gat), .A2(G233gat), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n604), .B(new_n605), .C1(new_n356), .C2(new_n603), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT18), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G113gat), .B(G141gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G169gat), .B(G197gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n608), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n340), .B(KEYINPUT17), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(new_n316), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n618), .A2(new_n604), .A3(KEYINPUT18), .A4(new_n605), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT88), .B(KEYINPUT13), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(new_n605), .ZN(new_n621));
  INV_X1    g420(.A(new_n340), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n316), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n340), .B1(new_n314), .B2(new_n315), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n621), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n619), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n602), .B1(new_n616), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n614), .B1(new_n606), .B2(new_n607), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n628), .A2(KEYINPUT90), .A3(new_n625), .A4(new_n619), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT89), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n619), .A2(new_n625), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n608), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n631), .B1(new_n619), .B2(new_n625), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n614), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(KEYINPUT91), .B1(new_n601), .B2(new_n636), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n589), .A2(new_n599), .A3(new_n596), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n599), .B1(new_n589), .B2(new_n596), .ZN(new_n639));
  OAI211_X1 g438(.A(KEYINPUT91), .B(new_n636), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n394), .B1(new_n637), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT99), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT91), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n638), .A2(new_n639), .ZN(new_n646));
  INV_X1    g445(.A(new_n636), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n640), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n649), .A2(KEYINPUT99), .A3(new_n394), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n288), .B1(new_n644), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(new_n306), .ZN(G1324gat));
  INV_X1    g451(.A(KEYINPUT101), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT16), .B(G8gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT100), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT42), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(KEYINPUT99), .B1(new_n649), .B2(new_n394), .ZN(new_n658));
  INV_X1    g457(.A(new_n394), .ZN(new_n659));
  AOI211_X1 g458(.A(new_n643), .B(new_n659), .C1(new_n648), .C2(new_n640), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n519), .B(new_n657), .C1(new_n658), .C2(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n586), .B1(new_n644), .B2(new_n650), .ZN(new_n662));
  INV_X1    g461(.A(G8gat), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n655), .ZN(new_n665));
  AOI21_X1  g464(.A(KEYINPUT42), .B1(new_n662), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n653), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n519), .B1(new_n658), .B2(new_n660), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n656), .B1(new_n668), .B2(new_n655), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(G8gat), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n669), .A2(KEYINPUT101), .A3(new_n661), .A4(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n667), .A2(new_n671), .ZN(G1325gat));
  NAND2_X1  g471(.A1(new_n578), .A2(new_n583), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(G15gat), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n674), .B1(new_n644), .B2(new_n650), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n593), .B1(new_n658), .B2(new_n660), .ZN(new_n676));
  INV_X1    g475(.A(G15gat), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT102), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n676), .A2(KEYINPUT102), .A3(new_n677), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n675), .B1(new_n680), .B2(new_n681), .ZN(G1326gat));
  AOI21_X1  g481(.A(new_n435), .B1(new_n644), .B2(new_n650), .ZN(new_n683));
  XOR2_X1   g482(.A(KEYINPUT43), .B(G22gat), .Z(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(G1327gat));
  NAND3_X1  g484(.A1(new_n601), .A2(KEYINPUT44), .A3(new_n370), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n369), .B1(new_n589), .B2(new_n596), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n687), .A2(KEYINPUT44), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n326), .A2(new_n392), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n689), .A2(new_n647), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n686), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n691), .A2(KEYINPUT103), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(KEYINPUT103), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n692), .A2(new_n693), .A3(new_n521), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(G29gat), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n689), .A2(new_n369), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n649), .A2(new_n327), .A3(new_n521), .A4(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT45), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OR2_X1    g498(.A1(new_n697), .A2(new_n698), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n695), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(KEYINPUT104), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n695), .A2(new_n703), .A3(new_n699), .A4(new_n700), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(G1328gat));
  AND2_X1   g504(.A1(new_n649), .A2(new_n696), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n706), .A2(new_n328), .A3(new_n519), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT46), .Z(new_n708));
  NAND3_X1  g507(.A1(new_n692), .A2(new_n693), .A3(new_n519), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n328), .B1(new_n709), .B2(KEYINPUT105), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n710), .B1(KEYINPUT105), .B2(new_n709), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n708), .A2(new_n711), .ZN(G1329gat));
  INV_X1    g511(.A(new_n691), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n673), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(G43gat), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n579), .A2(G43gat), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n706), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n715), .A2(new_n717), .A3(KEYINPUT47), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n692), .A2(new_n693), .A3(new_n673), .ZN(new_n719));
  AOI22_X1  g518(.A1(new_n719), .A2(G43gat), .B1(new_n706), .B2(new_n716), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n718), .B1(new_n720), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g520(.A1(new_n713), .A2(KEYINPUT106), .A3(new_n436), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n723), .B1(new_n691), .B2(new_n435), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n722), .A2(new_n724), .A3(G50gat), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n435), .A2(G50gat), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n706), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n725), .A2(KEYINPUT48), .A3(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n692), .A2(new_n693), .A3(new_n436), .ZN(new_n729));
  AOI22_X1  g528(.A1(new_n729), .A2(G50gat), .B1(new_n706), .B2(new_n726), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n728), .B1(new_n730), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR4_X1   g530(.A1(new_n326), .A2(new_n636), .A3(new_n370), .A4(new_n392), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n597), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT107), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n521), .B(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  XOR2_X1   g535(.A(KEYINPUT108), .B(G57gat), .Z(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1332gat));
  XNOR2_X1  g537(.A(new_n733), .B(KEYINPUT109), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n519), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n740), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n741));
  XOR2_X1   g540(.A(KEYINPUT49), .B(G64gat), .Z(new_n742));
  OAI21_X1  g541(.A(new_n741), .B1(new_n740), .B2(new_n742), .ZN(G1333gat));
  AOI21_X1  g542(.A(G71gat), .B1(new_n733), .B2(new_n593), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n673), .A2(G71gat), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n744), .B1(new_n739), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1334gat));
  NAND2_X1  g547(.A1(new_n739), .A2(new_n436), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G78gat), .ZN(G1335gat));
  INV_X1    g549(.A(new_n326), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n751), .A2(new_n636), .A3(new_n392), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n686), .A2(new_n688), .A3(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(G85gat), .B1(new_n753), .B2(new_n288), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n687), .A2(new_n647), .A3(new_n326), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT51), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n755), .A2(new_n756), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n288), .A2(new_n392), .A3(G85gat), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT111), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n754), .B1(new_n759), .B2(new_n761), .ZN(G1336gat));
  NOR2_X1   g561(.A1(new_n759), .A2(new_n392), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n763), .A2(new_n345), .A3(new_n519), .ZN(new_n764));
  OAI21_X1  g563(.A(G92gat), .B1(new_n753), .B2(new_n586), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT52), .ZN(G1337gat));
  INV_X1    g566(.A(G99gat), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n763), .A2(new_n768), .A3(new_n593), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n753), .B1(new_n578), .B2(new_n583), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n769), .B1(new_n770), .B2(new_n768), .ZN(G1338gat));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n686), .A2(new_n436), .A3(new_n688), .A4(new_n752), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(G106gat), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n435), .A2(G106gat), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n393), .B(new_n775), .C1(new_n757), .C2(new_n758), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n772), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(G106gat), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n778), .B1(new_n773), .B2(KEYINPUT112), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(KEYINPUT112), .B2(new_n773), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n776), .A2(new_n772), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n777), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT113), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n782), .B(new_n783), .ZN(G1339gat));
  INV_X1    g583(.A(KEYINPUT116), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n384), .A2(new_n377), .A3(new_n385), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT114), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n384), .A2(new_n789), .A3(new_n377), .A4(new_n385), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n386), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n386), .A2(new_n792), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n375), .ZN(new_n797));
  OAI211_X1 g596(.A(KEYINPUT115), .B(new_n786), .C1(new_n795), .C2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n797), .B1(new_n791), .B2(new_n793), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n799), .B1(new_n800), .B2(KEYINPUT55), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n794), .A2(KEYINPUT55), .A3(new_n375), .A4(new_n796), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n388), .A2(new_n374), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n802), .A2(new_n636), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n618), .A2(new_n604), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n808), .A2(G229gat), .A3(G233gat), .ZN(new_n809));
  OR3_X1    g608(.A1(new_n623), .A2(new_n624), .A3(new_n621), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n613), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(new_n627), .B2(new_n629), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n393), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n370), .B1(new_n807), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n812), .A2(new_n370), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n805), .B1(new_n801), .B2(new_n798), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n785), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n815), .A2(new_n816), .ZN(new_n819));
  AOI22_X1  g618(.A1(new_n816), .A2(new_n636), .B1(new_n393), .B2(new_n812), .ZN(new_n820));
  OAI211_X1 g619(.A(KEYINPUT116), .B(new_n819), .C1(new_n820), .C2(new_n370), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n818), .A2(new_n326), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n394), .A2(new_n647), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n288), .A2(new_n519), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n824), .A2(new_n593), .A3(new_n435), .A4(new_n825), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n826), .A2(new_n215), .A3(new_n647), .ZN(new_n827));
  INV_X1    g626(.A(new_n735), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n828), .B1(new_n822), .B2(new_n823), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n830), .A2(new_n519), .A3(new_n590), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n636), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n827), .B1(new_n832), .B2(new_n215), .ZN(G1340gat));
  NOR3_X1   g632(.A1(new_n826), .A2(new_n213), .A3(new_n392), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n831), .A2(new_n393), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n834), .B1(new_n835), .B2(new_n213), .ZN(G1341gat));
  NAND3_X1  g635(.A1(new_n831), .A2(new_n207), .A3(new_n751), .ZN(new_n837));
  OAI21_X1  g636(.A(G127gat), .B1(new_n826), .B2(new_n326), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(G1342gat));
  NAND2_X1  g638(.A1(new_n370), .A2(new_n586), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(KEYINPUT117), .ZN(new_n841));
  OR4_X1    g640(.A1(G134gat), .A2(new_n830), .A3(new_n590), .A4(new_n841), .ZN(new_n842));
  OR2_X1    g641(.A1(new_n842), .A2(KEYINPUT56), .ZN(new_n843));
  OAI21_X1  g642(.A(G134gat), .B1(new_n826), .B2(new_n369), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(KEYINPUT56), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(G1343gat));
  NAND2_X1  g645(.A1(new_n830), .A2(KEYINPUT119), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n673), .A2(new_n435), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n849), .B1(new_n829), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n647), .A2(G141gat), .ZN(new_n852));
  AND4_X1   g651(.A1(new_n586), .A2(new_n847), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n853), .A2(KEYINPUT58), .ZN(new_n854));
  INV_X1    g653(.A(new_n825), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n673), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT57), .B1(new_n824), .B2(new_n436), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n786), .B1(new_n795), .B2(new_n797), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n636), .A2(new_n806), .A3(new_n858), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n859), .A2(new_n813), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n819), .B1(new_n860), .B2(new_n370), .ZN(new_n861));
  AOI22_X1  g660(.A1(new_n861), .A2(new_n326), .B1(new_n647), .B2(new_n394), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n435), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n856), .B1(new_n857), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(G141gat), .B1(new_n867), .B2(new_n647), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n854), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(KEYINPUT118), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n435), .B1(new_n822), .B2(new_n823), .ZN(new_n871));
  OAI22_X1  g670(.A1(new_n871), .A2(KEYINPUT57), .B1(new_n865), .B2(new_n862), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n872), .A2(new_n873), .A3(new_n856), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n870), .A2(new_n636), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n853), .B1(new_n875), .B2(G141gat), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT58), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n869), .B1(new_n876), .B2(new_n877), .ZN(G1344gat));
  AND2_X1   g677(.A1(new_n847), .A2(new_n851), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n879), .A2(new_n586), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n231), .A3(new_n393), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT59), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(G148gat), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n872), .A2(new_n873), .A3(new_n856), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n873), .B1(new_n872), .B2(new_n856), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n883), .B1(new_n886), .B2(new_n393), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n863), .B1(new_n862), .B2(new_n435), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n822), .A2(new_n823), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n888), .B1(new_n889), .B2(new_n865), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n673), .A2(new_n392), .A3(new_n855), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI211_X1 g691(.A(KEYINPUT120), .B(KEYINPUT59), .C1(new_n892), .C2(new_n231), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT120), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n231), .B1(new_n890), .B2(new_n891), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n894), .B1(new_n895), .B2(new_n882), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n881), .B1(new_n887), .B2(new_n897), .ZN(G1345gat));
  NAND3_X1  g697(.A1(new_n880), .A2(new_n224), .A3(new_n751), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n870), .A2(new_n874), .ZN(new_n900));
  OAI21_X1  g699(.A(G155gat), .B1(new_n900), .B2(new_n326), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(G1346gat));
  OAI21_X1  g701(.A(G162gat), .B1(new_n900), .B2(new_n369), .ZN(new_n903));
  INV_X1    g702(.A(new_n841), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n879), .A2(new_n225), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(G1347gat));
  NOR2_X1   g705(.A1(new_n889), .A2(new_n521), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n590), .A2(new_n586), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT121), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(G169gat), .B1(new_n910), .B2(new_n636), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n735), .A2(new_n586), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n912), .B1(new_n914), .B2(new_n579), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n913), .A2(KEYINPUT122), .A3(new_n593), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n915), .A2(new_n435), .A3(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n889), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n647), .A2(new_n478), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n911), .B1(new_n918), .B2(new_n919), .ZN(G1348gat));
  NAND3_X1  g719(.A1(new_n910), .A2(new_n479), .A3(new_n393), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n889), .A2(new_n392), .A3(new_n917), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n921), .B1(new_n479), .B2(new_n922), .ZN(G1349gat));
  NAND2_X1  g722(.A1(new_n918), .A2(new_n751), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT123), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT123), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n918), .A2(new_n926), .A3(new_n751), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n925), .A2(G183gat), .A3(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n326), .A2(new_n460), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n930));
  AOI22_X1  g729(.A1(new_n910), .A2(new_n929), .B1(new_n930), .B2(KEYINPUT60), .ZN(new_n931));
  OR2_X1    g730(.A1(new_n930), .A2(KEYINPUT60), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n928), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n932), .B1(new_n928), .B2(new_n931), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n933), .A2(new_n934), .ZN(G1350gat));
  AOI21_X1  g734(.A(new_n463), .B1(new_n918), .B2(new_n370), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n937));
  OR3_X1    g736(.A1(new_n936), .A2(new_n937), .A3(KEYINPUT61), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n910), .A2(new_n463), .A3(new_n370), .ZN(new_n939));
  OAI21_X1  g738(.A(KEYINPUT61), .B1(new_n936), .B2(new_n937), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n936), .A2(new_n937), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n938), .B(new_n939), .C1(new_n940), .C2(new_n941), .ZN(G1351gat));
  NOR4_X1   g741(.A1(new_n889), .A2(new_n521), .A3(new_n586), .A4(new_n849), .ZN(new_n943));
  AOI21_X1  g742(.A(G197gat), .B1(new_n943), .B2(new_n636), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT126), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n890), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n914), .A2(new_n673), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n890), .A2(new_n945), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n636), .A2(G197gat), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n944), .B1(new_n950), .B2(new_n951), .ZN(G1352gat));
  OAI21_X1  g751(.A(G204gat), .B1(new_n949), .B2(new_n392), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT127), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n392), .A2(G204gat), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n943), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n955), .B1(new_n943), .B2(new_n956), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n954), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(new_n959), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n961), .A2(new_n957), .A3(KEYINPUT62), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n953), .A2(new_n960), .A3(new_n962), .ZN(G1353gat));
  NAND3_X1  g762(.A1(new_n890), .A2(new_n751), .A3(new_n947), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(G211gat), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT63), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n965), .B(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(G211gat), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n943), .A2(new_n968), .A3(new_n751), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(new_n969), .ZN(G1354gat));
  AOI21_X1  g769(.A(G218gat), .B1(new_n943), .B2(new_n370), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n370), .A2(G218gat), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n971), .B1(new_n950), .B2(new_n972), .ZN(G1355gat));
endmodule


