

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760;

  INV_X1 U378 ( .A(KEYINPUT64), .ZN(n459) );
  XNOR2_X1 U379 ( .A(n459), .B(G953), .ZN(n748) );
  INV_X1 U380 ( .A(n614), .ZN(n700) );
  BUF_X2 U381 ( .A(n724), .Z(n728) );
  AND2_X2 U382 ( .A1(n629), .A2(n630), .ZN(n472) );
  NAND2_X2 U383 ( .A1(n755), .A2(KEYINPUT44), .ZN(n629) );
  XNOR2_X1 U384 ( .A(n400), .B(n494), .ZN(n744) );
  XNOR2_X2 U385 ( .A(n567), .B(n493), .ZN(n400) );
  NAND2_X1 U386 ( .A1(n601), .A2(n580), .ZN(n683) );
  NOR2_X1 U387 ( .A1(n579), .A2(n584), .ZN(n669) );
  NOR2_X2 U388 ( .A1(n619), .A2(n569), .ZN(n690) );
  NOR2_X1 U389 ( .A1(n578), .A2(n634), .ZN(n675) );
  XNOR2_X1 U390 ( .A(n387), .B(n365), .ZN(n758) );
  NOR2_X1 U391 ( .A1(n602), .A2(n580), .ZN(n387) );
  NOR2_X1 U392 ( .A1(n613), .A2(n464), .ZN(n611) );
  AND2_X1 U393 ( .A1(n398), .A2(n397), .ZN(n396) );
  XNOR2_X1 U394 ( .A(n377), .B(G478), .ZN(n584) );
  NAND2_X1 U395 ( .A1(n483), .A2(n488), .ZN(n382) );
  XNOR2_X1 U396 ( .A(n457), .B(n456), .ZN(n498) );
  XNOR2_X1 U397 ( .A(n458), .B(n495), .ZN(n457) );
  XOR2_X1 U398 ( .A(G131), .B(G134), .Z(n494) );
  XNOR2_X1 U399 ( .A(G113), .B(KEYINPUT3), .ZN(n506) );
  NOR2_X1 U400 ( .A1(n716), .A2(n615), .ZN(n433) );
  XNOR2_X1 U401 ( .A(n379), .B(KEYINPUT72), .ZN(n420) );
  NAND2_X1 U402 ( .A1(n380), .A2(n360), .ZN(n379) );
  XNOR2_X1 U403 ( .A(n593), .B(n381), .ZN(n380) );
  INV_X1 U404 ( .A(KEYINPUT73), .ZN(n381) );
  NOR2_X1 U405 ( .A1(n758), .A2(n759), .ZN(n411) );
  OR2_X1 U406 ( .A1(G237), .A2(G902), .ZN(n518) );
  NAND2_X1 U407 ( .A1(n690), .A2(n576), .ZN(n393) );
  XOR2_X1 U408 ( .A(KEYINPUT41), .B(n572), .Z(n715) );
  XNOR2_X1 U409 ( .A(G140), .B(KEYINPUT101), .ZN(n549) );
  XNOR2_X1 U410 ( .A(G113), .B(G122), .ZN(n552) );
  XOR2_X1 U411 ( .A(G146), .B(G125), .Z(n520) );
  NOR2_X1 U412 ( .A1(n384), .A2(KEYINPUT88), .ZN(n383) );
  INV_X1 U413 ( .A(n485), .ZN(n385) );
  NOR2_X1 U414 ( .A1(n490), .A2(n675), .ZN(n409) );
  NOR2_X1 U415 ( .A1(G953), .A2(G237), .ZN(n544) );
  INV_X1 U416 ( .A(KEYINPUT4), .ZN(n493) );
  XOR2_X1 U417 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n513) );
  XNOR2_X1 U418 ( .A(n520), .B(n512), .ZN(n489) );
  XOR2_X1 U419 ( .A(KEYINPUT77), .B(KEYINPUT89), .Z(n512) );
  NAND2_X1 U420 ( .A1(n649), .A2(n519), .ZN(n488) );
  OR2_X1 U421 ( .A1(n720), .A2(n485), .ZN(n416) );
  XNOR2_X1 U422 ( .A(n448), .B(n447), .ZN(n577) );
  INV_X1 U423 ( .A(KEYINPUT69), .ZN(n447) );
  AND2_X1 U424 ( .A1(n694), .A2(n450), .ZN(n449) );
  INV_X1 U425 ( .A(n569), .ZN(n693) );
  INV_X1 U426 ( .A(KEYINPUT99), .ZN(n478) );
  XOR2_X1 U427 ( .A(KEYINPUT25), .B(KEYINPUT97), .Z(n530) );
  XNOR2_X1 U428 ( .A(KEYINPUT96), .B(KEYINPUT95), .ZN(n529) );
  INV_X1 U429 ( .A(G469), .ZN(n460) );
  XOR2_X1 U430 ( .A(KEYINPUT5), .B(KEYINPUT74), .Z(n503) );
  XNOR2_X1 U431 ( .A(n413), .B(n412), .ZN(n515) );
  XNOR2_X1 U432 ( .A(n505), .B(KEYINPUT70), .ZN(n412) );
  XNOR2_X1 U433 ( .A(n507), .B(n506), .ZN(n413) );
  INV_X1 U434 ( .A(G101), .ZN(n505) );
  NAND2_X1 U435 ( .A1(n462), .A2(n669), .ZN(n594) );
  NOR2_X1 U436 ( .A1(n577), .A2(n464), .ZN(n462) );
  XNOR2_X1 U437 ( .A(n389), .B(n388), .ZN(n602) );
  INV_X1 U438 ( .A(KEYINPUT39), .ZN(n388) );
  XNOR2_X1 U439 ( .A(n594), .B(n415), .ZN(n414) );
  INV_X1 U440 ( .A(KEYINPUT110), .ZN(n415) );
  XNOR2_X1 U441 ( .A(KEYINPUT68), .B(KEYINPUT0), .ZN(n609) );
  XNOR2_X1 U442 ( .A(n570), .B(KEYINPUT28), .ZN(n453) );
  NOR2_X1 U443 ( .A1(n614), .A2(n577), .ZN(n570) );
  XNOR2_X1 U444 ( .A(n378), .B(n566), .ZN(n726) );
  XNOR2_X1 U445 ( .A(n722), .B(n721), .ZN(n723) );
  NAND2_X1 U446 ( .A1(n364), .A2(n718), .ZN(n480) );
  XNOR2_X1 U447 ( .A(n714), .B(n482), .ZN(n481) );
  INV_X1 U448 ( .A(KEYINPUT81), .ZN(n482) );
  NAND2_X1 U449 ( .A1(n527), .A2(n486), .ZN(n485) );
  INV_X1 U450 ( .A(n519), .ZN(n486) );
  XNOR2_X1 U451 ( .A(G116), .B(G119), .ZN(n507) );
  XNOR2_X1 U452 ( .A(n551), .B(n431), .ZN(n553) );
  XNOR2_X1 U453 ( .A(n552), .B(n432), .ZN(n431) );
  INV_X1 U454 ( .A(KEYINPUT102), .ZN(n432) );
  XNOR2_X1 U455 ( .A(G143), .B(G131), .ZN(n547) );
  XOR2_X1 U456 ( .A(KEYINPUT11), .B(G104), .Z(n548) );
  XNOR2_X1 U457 ( .A(n520), .B(KEYINPUT10), .ZN(n545) );
  XOR2_X1 U458 ( .A(KEYINPUT92), .B(G101), .Z(n495) );
  INV_X1 U459 ( .A(n521), .ZN(n456) );
  AND2_X1 U460 ( .A1(n589), .A2(n450), .ZN(n491) );
  XNOR2_X1 U461 ( .A(n611), .B(KEYINPUT33), .ZN(n716) );
  NAND2_X1 U462 ( .A1(G214), .A2(n518), .ZN(n502) );
  INV_X1 U463 ( .A(KEYINPUT48), .ZN(n410) );
  XNOR2_X1 U464 ( .A(n496), .B(G107), .ZN(n514) );
  XNOR2_X1 U465 ( .A(G104), .B(G110), .ZN(n496) );
  INV_X1 U466 ( .A(KEYINPUT45), .ZN(n645) );
  XNOR2_X1 U467 ( .A(n525), .B(n443), .ZN(n564) );
  INV_X1 U468 ( .A(KEYINPUT8), .ZN(n443) );
  XNOR2_X1 U469 ( .A(n526), .B(n359), .ZN(n392) );
  XNOR2_X1 U470 ( .A(KEYINPUT24), .B(KEYINPUT93), .ZN(n522) );
  XNOR2_X1 U471 ( .A(n545), .B(n521), .ZN(n746) );
  XNOR2_X1 U472 ( .A(G116), .B(G134), .ZN(n559) );
  XNOR2_X1 U473 ( .A(G107), .B(KEYINPUT7), .ZN(n560) );
  XNOR2_X1 U474 ( .A(n376), .B(KEYINPUT9), .ZN(n561) );
  INV_X1 U475 ( .A(KEYINPUT104), .ZN(n376) );
  XNOR2_X1 U476 ( .A(n403), .B(n400), .ZN(n517) );
  XNOR2_X1 U477 ( .A(n489), .B(n404), .ZN(n403) );
  XNOR2_X1 U478 ( .A(n405), .B(n513), .ZN(n404) );
  BUF_X1 U479 ( .A(n716), .Z(n419) );
  NOR2_X1 U480 ( .A1(n710), .A2(KEYINPUT2), .ZN(n711) );
  INV_X1 U481 ( .A(KEYINPUT78), .ZN(n463) );
  XNOR2_X1 U482 ( .A(n393), .B(KEYINPUT107), .ZN(n589) );
  OR2_X1 U483 ( .A1(n726), .A2(G902), .ZN(n377) );
  AND2_X1 U484 ( .A1(n615), .A2(n478), .ZN(n473) );
  NAND2_X1 U485 ( .A1(n475), .A2(n476), .ZN(n474) );
  AND2_X1 U486 ( .A1(n477), .A2(n614), .ZN(n476) );
  XNOR2_X1 U487 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U488 ( .A(n509), .B(n504), .ZN(n468) );
  XNOR2_X1 U489 ( .A(n515), .B(n508), .ZN(n509) );
  XNOR2_X1 U490 ( .A(n516), .B(n515), .ZN(n741) );
  XNOR2_X1 U491 ( .A(n514), .B(n434), .ZN(n516) );
  XNOR2_X1 U492 ( .A(n435), .B(KEYINPUT16), .ZN(n434) );
  INV_X1 U493 ( .A(G122), .ZN(n435) );
  XNOR2_X1 U494 ( .A(n372), .B(n442), .ZN(n727) );
  AND2_X1 U495 ( .A1(n564), .A2(G221), .ZN(n442) );
  XNOR2_X1 U496 ( .A(n746), .B(n391), .ZN(n372) );
  XNOR2_X1 U497 ( .A(n524), .B(n392), .ZN(n391) );
  NOR2_X1 U498 ( .A1(n582), .A2(n715), .ZN(n573) );
  INV_X1 U499 ( .A(KEYINPUT109), .ZN(n461) );
  XNOR2_X1 U500 ( .A(n470), .B(n469), .ZN(n578) );
  XNOR2_X1 U501 ( .A(KEYINPUT36), .B(KEYINPUT87), .ZN(n469) );
  AND2_X1 U502 ( .A1(n414), .A2(n581), .ZN(n470) );
  AND2_X1 U503 ( .A1(n579), .A2(n584), .ZN(n671) );
  NOR2_X1 U504 ( .A1(n421), .A2(n452), .ZN(n451) );
  INV_X1 U505 ( .A(n571), .ZN(n452) );
  XNOR2_X1 U506 ( .A(n639), .B(KEYINPUT106), .ZN(n756) );
  BUF_X1 U507 ( .A(n659), .Z(n422) );
  XNOR2_X1 U508 ( .A(n725), .B(n726), .ZN(n417) );
  INV_X1 U509 ( .A(KEYINPUT56), .ZN(n439) );
  NAND2_X1 U510 ( .A1(n481), .A2(n479), .ZN(n418) );
  NOR2_X1 U511 ( .A1(n719), .A2(n480), .ZN(n479) );
  AND2_X1 U512 ( .A1(n416), .A2(n484), .ZN(n357) );
  AND2_X1 U513 ( .A1(n608), .A2(n607), .ZN(n358) );
  XOR2_X1 U514 ( .A(G119), .B(G128), .Z(n359) );
  INV_X1 U515 ( .A(n587), .ZN(n450) );
  AND2_X1 U516 ( .A1(n453), .A2(n451), .ZN(n360) );
  XOR2_X1 U517 ( .A(KEYINPUT38), .B(n597), .Z(n679) );
  INV_X1 U518 ( .A(KEYINPUT88), .ZN(n399) );
  AND2_X1 U519 ( .A1(n585), .A2(n584), .ZN(n361) );
  OR2_X1 U520 ( .A1(n393), .A2(n478), .ZN(n362) );
  AND2_X1 U521 ( .A1(n592), .A2(n666), .ZN(n363) );
  XNOR2_X1 U522 ( .A(KEYINPUT117), .B(n717), .ZN(n364) );
  XOR2_X1 U523 ( .A(n568), .B(n461), .Z(n365) );
  XNOR2_X1 U524 ( .A(n501), .B(n500), .ZN(n366) );
  INV_X1 U525 ( .A(n732), .ZN(n437) );
  XOR2_X1 U526 ( .A(n656), .B(KEYINPUT62), .Z(n367) );
  XNOR2_X1 U527 ( .A(n654), .B(KEYINPUT59), .ZN(n368) );
  XOR2_X1 U528 ( .A(n612), .B(KEYINPUT35), .Z(n369) );
  XOR2_X1 U529 ( .A(KEYINPUT118), .B(KEYINPUT53), .Z(n370) );
  XOR2_X1 U530 ( .A(KEYINPUT122), .B(KEYINPUT60), .Z(n371) );
  NAND2_X1 U531 ( .A1(n357), .A2(n395), .ZN(n394) );
  XNOR2_X1 U532 ( .A(n373), .B(n410), .ZN(n599) );
  NAND2_X1 U533 ( .A1(n408), .A2(n409), .ZN(n373) );
  NAND2_X1 U534 ( .A1(n569), .A2(n449), .ZN(n448) );
  INV_X1 U535 ( .A(n680), .ZN(n484) );
  NAND2_X1 U536 ( .A1(n386), .A2(n383), .ZN(n398) );
  NOR2_X1 U537 ( .A1(n680), .A2(n385), .ZN(n384) );
  NOR2_X1 U538 ( .A1(n656), .A2(G902), .ZN(n510) );
  XNOR2_X1 U539 ( .A(n433), .B(KEYINPUT34), .ZN(n402) );
  NAND2_X1 U540 ( .A1(n402), .A2(n361), .ZN(n401) );
  NAND2_X1 U541 ( .A1(n374), .A2(n375), .ZN(n646) );
  NAND2_X1 U542 ( .A1(n644), .A2(n643), .ZN(n374) );
  NAND2_X1 U543 ( .A1(n631), .A2(n471), .ZN(n375) );
  OR2_X2 U544 ( .A1(n710), .A2(KEYINPUT80), .ZN(n653) );
  NAND2_X1 U545 ( .A1(n618), .A2(n702), .ZN(n425) );
  XNOR2_X1 U546 ( .A(n567), .B(n565), .ZN(n378) );
  INV_X1 U547 ( .A(n382), .ZN(n487) );
  NOR2_X1 U548 ( .A1(n382), .A2(n399), .ZN(n395) );
  NAND2_X1 U549 ( .A1(n382), .A2(n399), .ZN(n397) );
  NAND2_X1 U550 ( .A1(n720), .A2(n484), .ZN(n386) );
  XNOR2_X2 U551 ( .A(n517), .B(n741), .ZN(n720) );
  NAND2_X1 U552 ( .A1(n491), .A2(n428), .ZN(n389) );
  XNOR2_X1 U553 ( .A(n390), .B(n468), .ZN(n656) );
  XNOR2_X2 U554 ( .A(n390), .B(n499), .ZN(n536) );
  XNOR2_X2 U555 ( .A(n744), .B(G146), .ZN(n390) );
  NAND2_X1 U556 ( .A1(n393), .A2(n478), .ZN(n477) );
  NAND2_X1 U557 ( .A1(n396), .A2(n394), .ZN(n581) );
  OR2_X2 U558 ( .A1(n604), .A2(n358), .ZN(n610) );
  XNOR2_X1 U559 ( .A(n581), .B(KEYINPUT19), .ZN(n604) );
  XNOR2_X2 U560 ( .A(n401), .B(n369), .ZN(n755) );
  NAND2_X1 U561 ( .A1(n748), .A2(G224), .ZN(n405) );
  NAND2_X1 U562 ( .A1(n406), .A2(n712), .ZN(n455) );
  NAND2_X1 U563 ( .A1(n710), .A2(KEYINPUT2), .ZN(n712) );
  NAND2_X1 U564 ( .A1(n407), .A2(n652), .ZN(n406) );
  NAND2_X1 U565 ( .A1(n710), .A2(n647), .ZN(n407) );
  AND2_X2 U566 ( .A1(n444), .A2(n603), .ZN(n710) );
  XNOR2_X1 U567 ( .A(n411), .B(n575), .ZN(n408) );
  NAND2_X1 U568 ( .A1(n487), .A2(n416), .ZN(n597) );
  XNOR2_X2 U569 ( .A(n492), .B(G143), .ZN(n567) );
  NOR2_X1 U570 ( .A1(n417), .A2(n732), .ZN(G63) );
  XNOR2_X1 U571 ( .A(n418), .B(n370), .ZN(G75) );
  NAND2_X1 U572 ( .A1(n724), .A2(G475), .ZN(n655) );
  NAND2_X1 U573 ( .A1(n724), .A2(G469), .ZN(n454) );
  NAND2_X2 U574 ( .A1(n455), .A2(n653), .ZN(n724) );
  XNOR2_X2 U575 ( .A(n576), .B(KEYINPUT1), .ZN(n689) );
  XNOR2_X2 U576 ( .A(n537), .B(n460), .ZN(n576) );
  NAND2_X1 U577 ( .A1(n363), .A2(n420), .ZN(n490) );
  NAND2_X1 U578 ( .A1(n724), .A2(G210), .ZN(n441) );
  NOR2_X1 U579 ( .A1(n617), .A2(KEYINPUT47), .ZN(n593) );
  XNOR2_X1 U580 ( .A(n454), .B(n366), .ZN(n436) );
  BUF_X1 U581 ( .A(n604), .Z(n421) );
  XNOR2_X1 U582 ( .A(n441), .B(n723), .ZN(n423) );
  NAND2_X1 U583 ( .A1(n436), .A2(n437), .ZN(n429) );
  NAND2_X1 U584 ( .A1(n757), .A2(n756), .ZN(n641) );
  XNOR2_X2 U585 ( .A(n636), .B(KEYINPUT32), .ZN(n757) );
  NOR2_X2 U586 ( .A1(n672), .A2(n659), .ZN(n616) );
  NAND2_X1 U587 ( .A1(n423), .A2(n437), .ZN(n440) );
  NOR2_X1 U588 ( .A1(n424), .A2(n617), .ZN(n626) );
  XNOR2_X1 U589 ( .A(n616), .B(KEYINPUT100), .ZN(n424) );
  NAND2_X1 U590 ( .A1(n466), .A2(n437), .ZN(n465) );
  XNOR2_X2 U591 ( .A(n425), .B(KEYINPUT31), .ZN(n672) );
  XNOR2_X1 U592 ( .A(n467), .B(n367), .ZN(n466) );
  XNOR2_X2 U593 ( .A(n426), .B(n533), .ZN(n569) );
  NOR2_X1 U594 ( .A1(n727), .A2(G902), .ZN(n426) );
  BUF_X2 U595 ( .A(n748), .Z(n427) );
  NOR2_X1 U596 ( .A1(n586), .A2(n679), .ZN(n428) );
  XNOR2_X1 U597 ( .A(n429), .B(KEYINPUT121), .ZN(G54) );
  XNOR2_X1 U598 ( .A(n430), .B(n371), .ZN(G60) );
  NAND2_X1 U599 ( .A1(n438), .A2(n437), .ZN(n430) );
  NOR2_X2 U600 ( .A1(G902), .A2(n536), .ZN(n537) );
  NOR2_X2 U601 ( .A1(n474), .A2(n473), .ZN(n659) );
  NAND2_X1 U602 ( .A1(n472), .A2(n628), .ZN(n471) );
  XNOR2_X1 U603 ( .A(n655), .B(n368), .ZN(n438) );
  XNOR2_X1 U604 ( .A(n646), .B(n645), .ZN(n736) );
  XNOR2_X1 U605 ( .A(n440), .B(n439), .ZN(G51) );
  NAND2_X1 U606 ( .A1(n603), .A2(n677), .ZN(n446) );
  NOR2_X1 U607 ( .A1(n736), .A2(n445), .ZN(n444) );
  INV_X1 U608 ( .A(n677), .ZN(n445) );
  XNOR2_X1 U609 ( .A(n446), .B(n749), .ZN(n747) );
  NAND2_X1 U610 ( .A1(n453), .A2(n571), .ZN(n582) );
  NAND2_X1 U611 ( .A1(n427), .A2(G227), .ZN(n458) );
  XNOR2_X1 U612 ( .A(n464), .B(n463), .ZN(n633) );
  NAND2_X1 U613 ( .A1(n624), .A2(n464), .ZN(n625) );
  XNOR2_X2 U614 ( .A(n700), .B(KEYINPUT6), .ZN(n464) );
  XNOR2_X1 U615 ( .A(n465), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U616 ( .A1(n724), .A2(G472), .ZN(n467) );
  NOR2_X1 U617 ( .A1(n626), .A2(n657), .ZN(n628) );
  OR2_X2 U618 ( .A1(n615), .A2(n362), .ZN(n475) );
  NAND2_X1 U619 ( .A1(n720), .A2(n519), .ZN(n483) );
  XNOR2_X1 U620 ( .A(n503), .B(G137), .ZN(n504) );
  INV_X1 U621 ( .A(KEYINPUT40), .ZN(n568) );
  NOR2_X1 U622 ( .A1(n427), .A2(G952), .ZN(n732) );
  XNOR2_X1 U623 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n501) );
  XNOR2_X2 U624 ( .A(G128), .B(KEYINPUT66), .ZN(n492) );
  XOR2_X1 U625 ( .A(G137), .B(G140), .Z(n521) );
  XNOR2_X1 U626 ( .A(n514), .B(KEYINPUT76), .ZN(n497) );
  XNOR2_X1 U627 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U628 ( .A(n536), .B(KEYINPUT57), .ZN(n500) );
  XOR2_X1 U629 ( .A(KEYINPUT90), .B(n502), .Z(n680) );
  NAND2_X1 U630 ( .A1(n544), .A2(G210), .ZN(n508) );
  XNOR2_X2 U631 ( .A(n510), .B(G472), .ZN(n614) );
  NOR2_X1 U632 ( .A1(n680), .A2(n614), .ZN(n511) );
  XOR2_X1 U633 ( .A(KEYINPUT30), .B(n511), .Z(n586) );
  XOR2_X1 U634 ( .A(G902), .B(KEYINPUT15), .Z(n649) );
  NAND2_X1 U635 ( .A1(G210), .A2(n518), .ZN(n519) );
  XOR2_X1 U636 ( .A(KEYINPUT94), .B(KEYINPUT75), .Z(n523) );
  XNOR2_X1 U637 ( .A(n523), .B(n522), .ZN(n524) );
  NAND2_X1 U638 ( .A1(n427), .A2(G234), .ZN(n525) );
  XOR2_X1 U639 ( .A(KEYINPUT23), .B(G110), .Z(n526) );
  INV_X1 U640 ( .A(n649), .ZN(n527) );
  NAND2_X1 U641 ( .A1(G234), .A2(n527), .ZN(n528) );
  XNOR2_X1 U642 ( .A(KEYINPUT20), .B(n528), .ZN(n534) );
  NAND2_X1 U643 ( .A1(n534), .A2(G217), .ZN(n532) );
  XNOR2_X1 U644 ( .A(n530), .B(n529), .ZN(n531) );
  NAND2_X1 U645 ( .A1(n534), .A2(G221), .ZN(n535) );
  XOR2_X1 U646 ( .A(n535), .B(KEYINPUT21), .Z(n694) );
  XOR2_X1 U647 ( .A(n694), .B(KEYINPUT98), .Z(n619) );
  NAND2_X1 U648 ( .A1(G234), .A2(G237), .ZN(n538) );
  XNOR2_X1 U649 ( .A(n538), .B(KEYINPUT14), .ZN(n539) );
  NAND2_X1 U650 ( .A1(G952), .A2(n539), .ZN(n709) );
  NOR2_X1 U651 ( .A1(G953), .A2(n709), .ZN(n606) );
  INV_X1 U652 ( .A(n427), .ZN(n541) );
  NAND2_X1 U653 ( .A1(n539), .A2(G902), .ZN(n540) );
  XNOR2_X1 U654 ( .A(n540), .B(KEYINPUT91), .ZN(n605) );
  NAND2_X1 U655 ( .A1(n541), .A2(n605), .ZN(n542) );
  NOR2_X1 U656 ( .A1(G900), .A2(n542), .ZN(n543) );
  NOR2_X1 U657 ( .A1(n606), .A2(n543), .ZN(n587) );
  XNOR2_X1 U658 ( .A(KEYINPUT13), .B(G475), .ZN(n558) );
  NAND2_X1 U659 ( .A1(G214), .A2(n544), .ZN(n546) );
  XNOR2_X1 U660 ( .A(n546), .B(n545), .ZN(n556) );
  XNOR2_X1 U661 ( .A(n548), .B(n547), .ZN(n554) );
  XOR2_X1 U662 ( .A(KEYINPUT103), .B(KEYINPUT12), .Z(n550) );
  XNOR2_X1 U663 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U664 ( .A(n554), .B(n553), .Z(n555) );
  XNOR2_X1 U665 ( .A(n556), .B(n555), .ZN(n654) );
  NOR2_X1 U666 ( .A1(G902), .A2(n654), .ZN(n557) );
  XNOR2_X1 U667 ( .A(n558), .B(n557), .ZN(n585) );
  INV_X1 U668 ( .A(n585), .ZN(n579) );
  XNOR2_X1 U669 ( .A(n559), .B(G122), .ZN(n563) );
  XNOR2_X1 U670 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U671 ( .A(n563), .B(n562), .Z(n566) );
  NAND2_X1 U672 ( .A1(G217), .A2(n564), .ZN(n565) );
  INV_X1 U673 ( .A(n669), .ZN(n580) );
  XNOR2_X1 U674 ( .A(n576), .B(KEYINPUT108), .ZN(n571) );
  NOR2_X1 U675 ( .A1(n585), .A2(n584), .ZN(n681) );
  NOR2_X1 U676 ( .A1(n679), .A2(n680), .ZN(n684) );
  NAND2_X1 U677 ( .A1(n681), .A2(n684), .ZN(n572) );
  XNOR2_X1 U678 ( .A(n573), .B(KEYINPUT42), .ZN(n759) );
  XOR2_X1 U679 ( .A(KEYINPUT65), .B(KEYINPUT46), .Z(n574) );
  XNOR2_X1 U680 ( .A(KEYINPUT84), .B(n574), .ZN(n575) );
  INV_X1 U681 ( .A(n689), .ZN(n634) );
  XNOR2_X1 U682 ( .A(KEYINPUT105), .B(n671), .ZN(n601) );
  NAND2_X1 U683 ( .A1(n683), .A2(n360), .ZN(n583) );
  NAND2_X1 U684 ( .A1(n583), .A2(KEYINPUT47), .ZN(n592) );
  NOR2_X1 U685 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U686 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U687 ( .A1(n597), .A2(n590), .ZN(n591) );
  NAND2_X1 U688 ( .A1(n361), .A2(n591), .ZN(n666) );
  INV_X1 U689 ( .A(n683), .ZN(n617) );
  NOR2_X1 U690 ( .A1(n689), .A2(n594), .ZN(n595) );
  NAND2_X1 U691 ( .A1(n484), .A2(n595), .ZN(n596) );
  XNOR2_X1 U692 ( .A(n596), .B(KEYINPUT43), .ZN(n598) );
  NAND2_X1 U693 ( .A1(n598), .A2(n597), .ZN(n678) );
  NAND2_X1 U694 ( .A1(n599), .A2(n678), .ZN(n600) );
  XNOR2_X1 U695 ( .A(n600), .B(KEYINPUT83), .ZN(n603) );
  OR2_X1 U696 ( .A1(n602), .A2(n601), .ZN(n677) );
  INV_X1 U697 ( .A(G953), .ZN(n718) );
  NOR2_X1 U698 ( .A1(G898), .A2(n718), .ZN(n740) );
  NAND2_X1 U699 ( .A1(n605), .A2(n740), .ZN(n608) );
  INV_X1 U700 ( .A(n606), .ZN(n607) );
  XNOR2_X2 U701 ( .A(n610), .B(n609), .ZN(n615) );
  NAND2_X1 U702 ( .A1(n690), .A2(n689), .ZN(n613) );
  INV_X1 U703 ( .A(KEYINPUT82), .ZN(n612) );
  INV_X1 U704 ( .A(n615), .ZN(n618) );
  NOR2_X1 U705 ( .A1(n614), .A2(n613), .ZN(n702) );
  INV_X1 U706 ( .A(n619), .ZN(n620) );
  NAND2_X1 U707 ( .A1(n681), .A2(n620), .ZN(n621) );
  NOR2_X1 U708 ( .A1(n615), .A2(n621), .ZN(n623) );
  XNOR2_X1 U709 ( .A(KEYINPUT22), .B(KEYINPUT71), .ZN(n622) );
  XNOR2_X1 U710 ( .A(n623), .B(n622), .ZN(n632) );
  NOR2_X1 U711 ( .A1(n632), .A2(n689), .ZN(n624) );
  NOR2_X1 U712 ( .A1(n569), .A2(n625), .ZN(n657) );
  NAND2_X1 U713 ( .A1(n629), .A2(n628), .ZN(n627) );
  NAND2_X1 U714 ( .A1(n627), .A2(KEYINPUT85), .ZN(n631) );
  INV_X1 U715 ( .A(KEYINPUT85), .ZN(n630) );
  NOR2_X2 U716 ( .A1(n632), .A2(n693), .ZN(n638) );
  NOR2_X1 U717 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U718 ( .A1(n638), .A2(n635), .ZN(n636) );
  NOR2_X1 U719 ( .A1(n689), .A2(n700), .ZN(n637) );
  NAND2_X1 U720 ( .A1(n638), .A2(n637), .ZN(n639) );
  INV_X1 U721 ( .A(KEYINPUT44), .ZN(n642) );
  NAND2_X1 U722 ( .A1(KEYINPUT86), .A2(n642), .ZN(n640) );
  XNOR2_X1 U723 ( .A(n641), .B(n640), .ZN(n644) );
  NAND2_X1 U724 ( .A1(n755), .A2(n642), .ZN(n643) );
  AND2_X1 U725 ( .A1(n649), .A2(KEYINPUT80), .ZN(n647) );
  NAND2_X1 U726 ( .A1(n649), .A2(KEYINPUT2), .ZN(n648) );
  XNOR2_X1 U727 ( .A(n648), .B(KEYINPUT67), .ZN(n651) );
  NOR2_X1 U728 ( .A1(n649), .A2(KEYINPUT80), .ZN(n650) );
  NOR2_X1 U729 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U730 ( .A(G101), .B(n657), .Z(G3) );
  NAND2_X1 U731 ( .A1(n669), .A2(n422), .ZN(n658) );
  XNOR2_X1 U732 ( .A(G104), .B(n658), .ZN(G6) );
  XOR2_X1 U733 ( .A(KEYINPUT111), .B(KEYINPUT26), .Z(n661) );
  NAND2_X1 U734 ( .A1(n422), .A2(n671), .ZN(n660) );
  XNOR2_X1 U735 ( .A(n661), .B(n660), .ZN(n663) );
  XOR2_X1 U736 ( .A(G107), .B(KEYINPUT27), .Z(n662) );
  XNOR2_X1 U737 ( .A(n663), .B(n662), .ZN(G9) );
  XOR2_X1 U738 ( .A(G128), .B(KEYINPUT29), .Z(n665) );
  NAND2_X1 U739 ( .A1(n360), .A2(n671), .ZN(n664) );
  XNOR2_X1 U740 ( .A(n665), .B(n664), .ZN(G30) );
  XNOR2_X1 U741 ( .A(G143), .B(n666), .ZN(G45) );
  NAND2_X1 U742 ( .A1(n360), .A2(n669), .ZN(n667) );
  XNOR2_X1 U743 ( .A(n667), .B(KEYINPUT112), .ZN(n668) );
  XNOR2_X1 U744 ( .A(G146), .B(n668), .ZN(G48) );
  NAND2_X1 U745 ( .A1(n672), .A2(n669), .ZN(n670) );
  XNOR2_X1 U746 ( .A(n670), .B(G113), .ZN(G15) );
  XOR2_X1 U747 ( .A(G116), .B(KEYINPUT113), .Z(n674) );
  NAND2_X1 U748 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U749 ( .A(n674), .B(n673), .ZN(G18) );
  XNOR2_X1 U750 ( .A(G125), .B(n675), .ZN(n676) );
  XNOR2_X1 U751 ( .A(n676), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U752 ( .A(G134), .B(n677), .ZN(G36) );
  XNOR2_X1 U753 ( .A(G140), .B(n678), .ZN(G42) );
  NAND2_X1 U754 ( .A1(n680), .A2(n679), .ZN(n682) );
  NAND2_X1 U755 ( .A1(n682), .A2(n681), .ZN(n686) );
  NAND2_X1 U756 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U757 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U758 ( .A(KEYINPUT116), .B(n687), .Z(n688) );
  NOR2_X1 U759 ( .A1(n419), .A2(n688), .ZN(n706) );
  NOR2_X1 U760 ( .A1(n690), .A2(n689), .ZN(n692) );
  XNOR2_X1 U761 ( .A(KEYINPUT50), .B(KEYINPUT115), .ZN(n691) );
  XNOR2_X1 U762 ( .A(n692), .B(n691), .ZN(n698) );
  XOR2_X1 U763 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n696) );
  OR2_X1 U764 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U765 ( .A(n696), .B(n695), .ZN(n697) );
  NAND2_X1 U766 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U767 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U768 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U769 ( .A(KEYINPUT51), .B(n703), .Z(n704) );
  NOR2_X1 U770 ( .A1(n715), .A2(n704), .ZN(n705) );
  NOR2_X1 U771 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U772 ( .A(n707), .B(KEYINPUT52), .ZN(n708) );
  NOR2_X1 U773 ( .A1(n709), .A2(n708), .ZN(n719) );
  XNOR2_X1 U774 ( .A(n711), .B(KEYINPUT79), .ZN(n713) );
  NAND2_X1 U775 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U776 ( .A1(n419), .A2(n715), .ZN(n717) );
  XOR2_X1 U777 ( .A(KEYINPUT55), .B(KEYINPUT54), .Z(n722) );
  XNOR2_X1 U778 ( .A(n720), .B(KEYINPUT119), .ZN(n721) );
  NAND2_X1 U779 ( .A1(G478), .A2(n728), .ZN(n725) );
  XOR2_X1 U780 ( .A(n727), .B(KEYINPUT123), .Z(n730) );
  NAND2_X1 U781 ( .A1(G217), .A2(n728), .ZN(n729) );
  XNOR2_X1 U782 ( .A(n730), .B(n729), .ZN(n731) );
  NOR2_X1 U783 ( .A1(n732), .A2(n731), .ZN(G66) );
  NAND2_X1 U784 ( .A1(G224), .A2(G953), .ZN(n733) );
  XNOR2_X1 U785 ( .A(n733), .B(KEYINPUT124), .ZN(n734) );
  XNOR2_X1 U786 ( .A(KEYINPUT61), .B(n734), .ZN(n735) );
  AND2_X1 U787 ( .A1(n735), .A2(G898), .ZN(n738) );
  NOR2_X1 U788 ( .A1(G953), .A2(n736), .ZN(n737) );
  NOR2_X1 U789 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U790 ( .A(n739), .B(KEYINPUT125), .ZN(n743) );
  NOR2_X1 U791 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U792 ( .A(n743), .B(n742), .ZN(G69) );
  BUF_X1 U793 ( .A(n744), .Z(n745) );
  XOR2_X1 U794 ( .A(n746), .B(n745), .Z(n749) );
  NAND2_X1 U795 ( .A1(n427), .A2(n747), .ZN(n753) );
  XNOR2_X1 U796 ( .A(G227), .B(n749), .ZN(n750) );
  NAND2_X1 U797 ( .A1(n750), .A2(G900), .ZN(n751) );
  NAND2_X1 U798 ( .A1(G953), .A2(n751), .ZN(n752) );
  NAND2_X1 U799 ( .A1(n753), .A2(n752), .ZN(G72) );
  XOR2_X1 U800 ( .A(G122), .B(KEYINPUT126), .Z(n754) );
  XNOR2_X1 U801 ( .A(n755), .B(n754), .ZN(G24) );
  XNOR2_X1 U802 ( .A(n756), .B(G110), .ZN(G12) );
  XNOR2_X1 U803 ( .A(G119), .B(n757), .ZN(G21) );
  XOR2_X1 U804 ( .A(n758), .B(G131), .Z(G33) );
  XNOR2_X1 U805 ( .A(G137), .B(KEYINPUT127), .ZN(n760) );
  XNOR2_X1 U806 ( .A(n760), .B(n759), .ZN(G39) );
endmodule

