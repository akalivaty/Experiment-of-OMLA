//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n560, new_n562, new_n563, new_n564, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT66), .B(G2104), .ZN(new_n462));
  OAI211_X1 g037(.A(G137), .B(new_n461), .C1(new_n462), .C2(new_n460), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(G101), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n459), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI211_X1 g042(.A(KEYINPUT67), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n461), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(KEYINPUT65), .A3(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n476), .B1(new_n472), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n474), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n469), .A2(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n470), .A2(KEYINPUT66), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G2104), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n460), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(new_n466), .ZN(new_n488));
  INV_X1    g063(.A(G136), .ZN(new_n489));
  NOR2_X1   g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(new_n466), .B2(G112), .ZN(new_n491));
  OAI22_X1  g066(.A1(new_n488), .A2(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n487), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n492), .B1(G124), .B2(new_n494), .ZN(new_n495));
  XNOR2_X1  g070(.A(new_n495), .B(KEYINPUT68), .ZN(G162));
  XOR2_X1   g071(.A(KEYINPUT70), .B(KEYINPUT4), .Z(new_n497));
  NAND4_X1  g072(.A1(new_n473), .A2(new_n497), .A3(G138), .A4(new_n466), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n500));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  NOR4_X1   g076(.A1(new_n485), .A2(new_n501), .A3(G2105), .A4(new_n486), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n500), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n483), .A2(G2104), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n470), .A2(KEYINPUT66), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT3), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n507), .A2(G138), .A3(new_n466), .A4(new_n461), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT69), .A3(KEYINPUT4), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n499), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n466), .A2(G102), .A3(G2104), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n487), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n512), .B2(new_n466), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n510), .A2(new_n513), .ZN(G164));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G651), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT71), .ZN(new_n517));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n515), .A2(G651), .ZN(new_n519));
  NOR3_X1   g094(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT5), .ZN(new_n522));
  AND3_X1   g097(.A1(new_n522), .A2(KEYINPUT72), .A3(G543), .ZN(new_n523));
  AOI21_X1  g098(.A(KEYINPUT72), .B1(new_n522), .B2(G543), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n523), .A2(new_n524), .B1(new_n522), .B2(G543), .ZN(new_n525));
  NOR3_X1   g100(.A1(new_n517), .A2(new_n525), .A3(new_n519), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G88), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n521), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n525), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n530), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G651), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n529), .A2(new_n533), .ZN(G303));
  INV_X1    g109(.A(G303), .ZN(G166));
  NAND2_X1  g110(.A1(new_n526), .A2(G89), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n520), .A2(G51), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n530), .A2(G63), .A3(G651), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  NAND4_X1  g115(.A1(new_n536), .A2(new_n537), .A3(new_n538), .A4(new_n540), .ZN(G286));
  INV_X1    g116(.A(G286), .ZN(G168));
  NAND2_X1  g117(.A1(G77), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G64), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n525), .B2(new_n544), .ZN(new_n545));
  XOR2_X1   g120(.A(new_n545), .B(KEYINPUT73), .Z(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G651), .ZN(new_n547));
  AOI22_X1  g122(.A1(G90), .A2(new_n526), .B1(new_n520), .B2(G52), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  AOI22_X1  g125(.A1(G81), .A2(new_n526), .B1(new_n520), .B2(G43), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT75), .ZN(new_n552));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G56), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n525), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G651), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT74), .ZN(new_n557));
  AND2_X1   g132(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  AND3_X1   g134(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G36), .ZN(G176));
  XOR2_X1   g136(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n562));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n560), .A2(new_n564), .ZN(G188));
  INV_X1    g140(.A(KEYINPUT77), .ZN(new_n566));
  INV_X1    g141(.A(G91), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n527), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n526), .A2(KEYINPUT77), .A3(G91), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  XOR2_X1   g145(.A(new_n570), .B(KEYINPUT78), .Z(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n525), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n568), .A2(new_n569), .B1(G651), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n520), .A2(G53), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT9), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(G299));
  NAND2_X1  g152(.A1(new_n526), .A2(G87), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n520), .A2(G49), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n530), .B2(G74), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  AOI22_X1  g156(.A1(G86), .A2(new_n526), .B1(new_n520), .B2(G48), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n525), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G651), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n582), .A2(new_n586), .ZN(G305));
  AOI22_X1  g162(.A1(G85), .A2(new_n526), .B1(new_n520), .B2(G47), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n530), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n532), .B2(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n526), .A2(G92), .ZN(new_n592));
  XOR2_X1   g167(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n593));
  XNOR2_X1  g168(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n525), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n520), .A2(G54), .B1(new_n597), .B2(G651), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT80), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n591), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n591), .B1(new_n601), .B2(G868), .ZN(G321));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(G299), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(new_n604), .B2(G168), .ZN(G297));
  OAI21_X1  g181(.A(new_n605), .B1(new_n604), .B2(G168), .ZN(G280));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n601), .B1(new_n608), .B2(G860), .ZN(G148));
  NAND2_X1  g184(.A1(new_n552), .A2(new_n557), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(new_n604), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n600), .A2(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(new_n604), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT81), .Z(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n494), .A2(G123), .ZN(new_n616));
  INV_X1    g191(.A(new_n488), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G135), .ZN(new_n618));
  NOR2_X1   g193(.A1(G99), .A2(G2105), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(new_n466), .B2(G111), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n616), .B(new_n618), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT82), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT83), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2096), .ZN(new_n624));
  NOR4_X1   g199(.A1(new_n472), .A2(new_n505), .A3(new_n506), .A4(G2105), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT12), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2100), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n624), .A2(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2435), .ZN(new_n631));
  XOR2_X1   g206(.A(G2427), .B(G2438), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(KEYINPUT14), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2451), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2454), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n634), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G2443), .B(G2446), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n640), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(G14), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(G401));
  XOR2_X1   g220(.A(G2072), .B(G2078), .Z(new_n646));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT85), .B(KEYINPUT18), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n646), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2096), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2100), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n647), .A2(new_n648), .ZN(new_n654));
  AND2_X1   g229(.A1(new_n654), .A2(KEYINPUT17), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n650), .B1(new_n655), .B2(new_n649), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n653), .B(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n659), .A2(new_n660), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT20), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n665), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n662), .A2(new_n664), .A3(new_n666), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n669), .B(new_n670), .C1(new_n668), .C2(new_n667), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1991), .B(G1996), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G1981), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n673), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT86), .B(G1986), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n676), .B(new_n677), .Z(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(G229));
  INV_X1    g254(.A(G19), .ZN(new_n680));
  OAI21_X1  g255(.A(KEYINPUT91), .B1(new_n680), .B2(G16), .ZN(new_n681));
  OR3_X1    g256(.A1(new_n680), .A2(KEYINPUT91), .A3(G16), .ZN(new_n682));
  INV_X1    g257(.A(G16), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n681), .B(new_n682), .C1(new_n558), .C2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(G1341), .Z(new_n685));
  NAND2_X1  g260(.A1(G299), .A2(G16), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n683), .A2(KEYINPUT23), .A3(G20), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT23), .ZN(new_n688));
  INV_X1    g263(.A(G20), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n688), .B1(new_n689), .B2(G16), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n686), .A2(new_n687), .A3(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(G1956), .Z(new_n692));
  NAND2_X1  g267(.A1(new_n622), .A2(G29), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n685), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT25), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n617), .A2(G139), .ZN(new_n697));
  AOI22_X1  g272(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT93), .ZN(new_n699));
  AOI211_X1 g274(.A(new_n696), .B(new_n697), .C1(G2105), .C2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G29), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G29), .B2(G33), .ZN(new_n702));
  INV_X1    g277(.A(G2072), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n683), .A2(G21), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G168), .B2(new_n683), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT94), .B(G1966), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NOR3_X1   g283(.A1(new_n694), .A2(new_n704), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  INV_X1    g285(.A(G34), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n711), .A2(KEYINPUT24), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n711), .A2(KEYINPUT24), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n710), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G160), .B2(new_n710), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n715), .A2(G2084), .ZN(new_n716));
  NAND2_X1  g291(.A1(G162), .A2(G29), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G29), .B2(G35), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT29), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n716), .B1(new_n720), .B2(G2090), .ZN(new_n721));
  MUX2_X1   g296(.A(G24), .B(G290), .S(G16), .Z(new_n722));
  XOR2_X1   g297(.A(KEYINPUT87), .B(G1986), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n710), .A2(G25), .ZN(new_n725));
  INV_X1    g300(.A(G131), .ZN(new_n726));
  NOR2_X1   g301(.A1(G95), .A2(G2105), .ZN(new_n727));
  OAI21_X1  g302(.A(G2104), .B1(new_n466), .B2(G107), .ZN(new_n728));
  OAI22_X1  g303(.A1(new_n488), .A2(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G119), .B2(new_n494), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n725), .B1(new_n730), .B2(new_n710), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT35), .B(G1991), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n731), .B(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT36), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n724), .B(new_n734), .C1(KEYINPUT90), .C2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n683), .A2(G6), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n582), .A2(new_n586), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(new_n683), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT89), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT32), .B(G1981), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n683), .A2(G22), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G166), .B2(new_n683), .ZN(new_n744));
  INV_X1    g319(.A(G1971), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(G16), .A2(G23), .ZN(new_n747));
  INV_X1    g322(.A(G288), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(G16), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT33), .B(G1976), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n746), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n742), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT88), .B(KEYINPUT34), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n736), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n735), .A2(KEYINPUT90), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n709), .B(new_n721), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(G4), .A2(G16), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n601), .B2(G16), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G1348), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n757), .A2(new_n758), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n683), .A2(G5), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G171), .B2(new_n683), .ZN(new_n766));
  INV_X1    g341(.A(G1961), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(G2090), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n769), .B1(new_n770), .B2(new_n719), .ZN(new_n771));
  INV_X1    g346(.A(G26), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n772), .A2(G29), .ZN(new_n773));
  NOR2_X1   g348(.A1(G104), .A2(G2105), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT92), .Z(new_n775));
  OAI211_X1 g350(.A(new_n775), .B(G2104), .C1(G116), .C2(new_n466), .ZN(new_n776));
  INV_X1    g351(.A(G140), .ZN(new_n777));
  INV_X1    g352(.A(G128), .ZN(new_n778));
  OAI221_X1 g353(.A(new_n776), .B1(new_n488), .B2(new_n777), .C1(new_n493), .C2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n773), .B1(new_n779), .B2(G29), .ZN(new_n780));
  MUX2_X1   g355(.A(new_n773), .B(new_n780), .S(KEYINPUT28), .Z(new_n781));
  INV_X1    g356(.A(G2067), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n710), .A2(G27), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G164), .B2(new_n710), .ZN(new_n785));
  INV_X1    g360(.A(G2078), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT30), .B(G28), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n715), .A2(G2084), .B1(new_n710), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  AOI211_X1 g365(.A(new_n783), .B(new_n790), .C1(new_n703), .C2(new_n702), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n763), .A2(new_n764), .A3(new_n771), .A4(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G29), .A2(G32), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n494), .A2(G129), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n462), .A2(G105), .A3(new_n466), .ZN(new_n795));
  NAND3_X1  g370(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT26), .Z(new_n797));
  INV_X1    g372(.A(G141), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n795), .B(new_n797), .C1(new_n488), .C2(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n794), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n793), .B1(new_n800), .B2(G29), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT27), .ZN(new_n802));
  INV_X1    g377(.A(G1996), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT31), .B(G11), .Z(new_n805));
  NOR3_X1   g380(.A1(new_n792), .A2(new_n804), .A3(new_n805), .ZN(G311));
  AND3_X1   g381(.A1(new_n763), .A2(new_n771), .A3(new_n791), .ZN(new_n807));
  INV_X1    g382(.A(new_n804), .ZN(new_n808));
  INV_X1    g383(.A(new_n805), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n807), .A2(new_n808), .A3(new_n764), .A4(new_n809), .ZN(G150));
  NAND2_X1  g385(.A1(new_n520), .A2(G55), .ZN(new_n811));
  INV_X1    g386(.A(G93), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n527), .B2(new_n812), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n530), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n814), .A2(new_n532), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(G860), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT37), .ZN(new_n819));
  INV_X1    g394(.A(new_n816), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n558), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n610), .A2(new_n816), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT38), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n601), .A2(G559), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(KEYINPUT39), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT95), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n817), .B1(new_n826), .B2(KEYINPUT39), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n819), .B1(new_n828), .B2(new_n829), .ZN(G145));
  INV_X1    g405(.A(new_n513), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT96), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n504), .A2(new_n509), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(new_n498), .ZN(new_n834));
  AOI211_X1 g409(.A(KEYINPUT96), .B(new_n499), .C1(new_n504), .C2(new_n509), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n831), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n779), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n800), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n700), .ZN(new_n839));
  INV_X1    g414(.A(G142), .ZN(new_n840));
  NOR2_X1   g415(.A1(G106), .A2(G2105), .ZN(new_n841));
  OAI21_X1  g416(.A(G2104), .B1(new_n466), .B2(G118), .ZN(new_n842));
  OAI22_X1  g417(.A1(new_n488), .A2(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(G130), .B2(new_n494), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n626), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n730), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT97), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n839), .B(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(G162), .B(G160), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(new_n622), .Z(new_n850));
  AOI21_X1  g425(.A(G37), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n839), .A2(new_n846), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(KEYINPUT98), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n839), .A2(new_n847), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n850), .B(KEYINPUT99), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT98), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n839), .A2(new_n856), .A3(new_n846), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n853), .A2(new_n854), .A3(new_n855), .A4(new_n857), .ZN(new_n858));
  AND3_X1   g433(.A1(new_n851), .A2(new_n858), .A3(KEYINPUT100), .ZN(new_n859));
  AOI21_X1  g434(.A(KEYINPUT100), .B1(new_n851), .B2(new_n858), .ZN(new_n860));
  OAI21_X1  g435(.A(KEYINPUT40), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n851), .A2(new_n858), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT100), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT40), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n851), .A2(new_n858), .A3(KEYINPUT100), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n861), .A2(new_n867), .ZN(G395));
  NAND2_X1  g443(.A1(new_n820), .A2(new_n604), .ZN(new_n869));
  XNOR2_X1  g444(.A(G303), .B(new_n738), .ZN(new_n870));
  XNOR2_X1  g445(.A(G290), .B(new_n748), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n870), .B1(KEYINPUT101), .B2(new_n871), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n871), .A2(KEYINPUT101), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n872), .B(new_n873), .Z(new_n874));
  XOR2_X1   g449(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n612), .B(new_n823), .ZN(new_n877));
  OR2_X1    g452(.A1(G299), .A2(new_n599), .ZN(new_n878));
  NAND2_X1  g453(.A1(G299), .A2(new_n599), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n878), .A2(KEYINPUT41), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(KEYINPUT41), .B1(new_n878), .B2(new_n879), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n877), .A2(new_n883), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n878), .A2(new_n879), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n884), .B1(new_n885), .B2(new_n877), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n876), .B(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n869), .B1(new_n887), .B2(new_n604), .ZN(G295));
  OAI21_X1  g463(.A(new_n869), .B1(new_n887), .B2(new_n604), .ZN(G331));
  XNOR2_X1  g464(.A(G301), .B(G168), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n823), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(G301), .B(G286), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n892), .A2(new_n821), .A3(new_n822), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(KEYINPUT104), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n823), .A2(new_n895), .A3(new_n890), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(new_n882), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(KEYINPUT105), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n891), .A2(new_n893), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n885), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT105), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n894), .A2(new_n901), .A3(new_n882), .A4(new_n896), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n898), .A2(new_n874), .A3(new_n900), .A4(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(G37), .ZN(new_n904));
  INV_X1    g479(.A(new_n874), .ZN(new_n905));
  INV_X1    g480(.A(new_n885), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n906), .B1(new_n894), .B2(new_n896), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n899), .A2(new_n883), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n905), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n903), .A2(new_n904), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(KEYINPUT43), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n898), .A2(new_n900), .A3(new_n902), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n905), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n913), .A2(new_n904), .A3(new_n903), .ZN(new_n914));
  XOR2_X1   g489(.A(KEYINPUT103), .B(KEYINPUT43), .Z(new_n915));
  OAI211_X1 g490(.A(new_n911), .B(KEYINPUT44), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n915), .ZN(new_n918));
  INV_X1    g493(.A(new_n915), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n903), .A2(new_n904), .A3(new_n909), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n917), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AOI211_X1 g498(.A(KEYINPUT106), .B(KEYINPUT44), .C1(new_n918), .C2(new_n920), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n916), .B1(new_n923), .B2(new_n924), .ZN(G397));
  INV_X1    g500(.A(G1384), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT45), .B1(new_n836), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n465), .A2(new_n466), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT67), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n465), .A2(new_n459), .A3(new_n466), .ZN(new_n930));
  XNOR2_X1  g505(.A(KEYINPUT107), .B(G40), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n929), .A2(new_n480), .A3(new_n930), .A4(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT108), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n469), .A2(new_n934), .A3(new_n480), .A4(new_n931), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n927), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT109), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n779), .B(new_n782), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(new_n803), .B2(new_n800), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n937), .A2(G1996), .ZN(new_n941));
  AOI22_X1  g516(.A1(new_n938), .A2(new_n940), .B1(new_n800), .B2(new_n941), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n730), .A2(new_n733), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n730), .A2(new_n733), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n938), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n937), .A2(G1986), .A3(G290), .ZN(new_n947));
  XOR2_X1   g522(.A(new_n947), .B(KEYINPUT48), .Z(new_n948));
  AND2_X1   g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n939), .A2(new_n800), .ZN(new_n950));
  AOI22_X1  g525(.A1(new_n938), .A2(new_n950), .B1(KEYINPUT123), .B2(KEYINPUT46), .ZN(new_n951));
  NOR2_X1   g526(.A1(KEYINPUT123), .A2(KEYINPUT46), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n941), .B(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(KEYINPUT124), .B(KEYINPUT47), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n954), .B(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n942), .A2(new_n943), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(G2067), .B2(new_n779), .ZN(new_n958));
  AOI211_X1 g533(.A(new_n949), .B(new_n956), .C1(new_n938), .C2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(G303), .A2(G8), .ZN(new_n960));
  XOR2_X1   g535(.A(new_n960), .B(KEYINPUT55), .Z(new_n961));
  OAI21_X1  g536(.A(new_n926), .B1(new_n510), .B2(new_n513), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n936), .B1(new_n963), .B2(KEYINPUT45), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n836), .A2(KEYINPUT45), .A3(new_n926), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n508), .A2(KEYINPUT69), .A3(KEYINPUT4), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT69), .B1(new_n508), .B2(KEYINPUT4), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n498), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT96), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n833), .A2(new_n832), .A3(new_n498), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(G1384), .B1(new_n973), .B2(new_n831), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n974), .A2(KEYINPUT110), .A3(KEYINPUT45), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n964), .B1(new_n967), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n976), .A2(G1971), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n962), .A2(KEYINPUT50), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n978), .A2(new_n936), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT50), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n836), .A2(new_n980), .A3(new_n926), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(KEYINPUT111), .B(G2090), .Z(new_n983));
  NOR2_X1   g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI211_X1 g559(.A(G8), .B(new_n961), .C1(new_n977), .C2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n836), .A2(new_n936), .A3(new_n926), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n748), .A2(G1976), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n986), .A2(G8), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n748), .A2(G1976), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n988), .A2(new_n989), .A3(new_n990), .A4(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1981), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n738), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(G305), .A2(G1981), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT49), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT113), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n997), .B(new_n999), .ZN(new_n1000));
  OR2_X1    g575(.A1(new_n998), .A2(KEYINPUT113), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n1000), .A2(G8), .A3(new_n986), .A4(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n986), .A2(G8), .A3(new_n987), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT112), .B1(new_n1003), .B2(KEYINPUT52), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n1003), .A2(KEYINPUT52), .A3(new_n991), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n993), .B(new_n1002), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n985), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G8), .ZN(new_n1008));
  INV_X1    g583(.A(new_n986), .ZN(new_n1009));
  INV_X1    g584(.A(G1976), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1002), .A2(new_n1010), .A3(new_n748), .ZN(new_n1011));
  AOI211_X1 g586(.A(new_n1008), .B(new_n1009), .C1(new_n1011), .C2(new_n995), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT63), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1006), .ZN(new_n1014));
  INV_X1    g589(.A(new_n961), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n980), .B1(new_n836), .B2(new_n926), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n936), .B1(KEYINPUT50), .B2(new_n962), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n1016), .A2(new_n1017), .A3(new_n983), .ZN(new_n1018));
  INV_X1    g593(.A(new_n964), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT110), .B1(new_n974), .B2(KEYINPUT45), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n513), .B1(new_n971), .B2(new_n972), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT45), .ZN(new_n1022));
  NOR4_X1   g597(.A1(new_n1021), .A2(new_n966), .A3(new_n1022), .A4(G1384), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1019), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1018), .B1(new_n1024), .B2(new_n745), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1015), .B1(new_n1025), .B2(new_n1008), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1014), .A2(new_n1026), .A3(new_n985), .ZN(new_n1027));
  XNOR2_X1  g602(.A(KEYINPUT115), .B(G2084), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n979), .A2(new_n981), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n936), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT114), .B1(new_n927), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n963), .A2(KEYINPUT45), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1034), .B(new_n936), .C1(new_n974), .C2(KEYINPUT45), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1032), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G1966), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1030), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  OR3_X1    g613(.A1(new_n1038), .A2(new_n1008), .A3(G286), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1013), .B1(new_n1027), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(G8), .B1(new_n977), .B2(new_n984), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1013), .B1(new_n1041), .B2(new_n1015), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n1038), .A2(new_n1008), .A3(G286), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1042), .A2(new_n985), .A3(new_n1014), .A4(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1012), .B1(new_n1040), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1027), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT51), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1048), .A2(G168), .A3(new_n1029), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1047), .B1(new_n1049), .B2(G8), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1008), .B1(new_n1038), .B2(G168), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT51), .B1(new_n1038), .B2(G168), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1050), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT62), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1046), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1052), .A2(new_n1051), .ZN(new_n1056));
  AOI211_X1 g631(.A(G286), .B(new_n1030), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1057));
  OAI21_X1  g632(.A(KEYINPUT51), .B1(new_n1057), .B2(new_n1008), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1056), .A2(new_n1058), .A3(new_n1054), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1060), .A2(G2078), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1032), .A2(new_n1033), .A3(new_n1035), .A4(new_n1061), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1021), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n978), .A2(new_n936), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n767), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT53), .B1(new_n976), .B2(new_n786), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1059), .A2(G171), .A3(new_n1069), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1007), .B(new_n1045), .C1(new_n1055), .C2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(G171), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1060), .B1(new_n1024), .B2(G2078), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT120), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1065), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n982), .A2(KEYINPUT120), .A3(new_n767), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(G160), .A2(new_n1061), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n836), .A2(new_n926), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1078), .B1(new_n1079), .B2(new_n1022), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1080), .B(G40), .C1(new_n1020), .C2(new_n1023), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1073), .A2(G301), .A3(new_n1077), .A4(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1072), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n1084));
  AOI22_X1  g659(.A1(new_n1056), .A2(new_n1058), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1084), .B1(new_n1068), .B2(G301), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT120), .B1(new_n982), .B2(new_n767), .ZN(new_n1087));
  AOI211_X1 g662(.A(new_n1074), .B(G1961), .C1(new_n979), .C2(new_n981), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1081), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT121), .B1(new_n1089), .B2(new_n1067), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1073), .A2(new_n1091), .A3(new_n1077), .A4(new_n1081), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1090), .A2(G171), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1027), .B1(new_n1086), .B2(new_n1093), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1085), .A2(new_n1094), .A3(KEYINPUT122), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT122), .B1(new_n1085), .B2(new_n1094), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1098), .A2(G1956), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT56), .B(G2072), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1099), .B1(new_n976), .B2(new_n1100), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n574), .B(new_n576), .C1(KEYINPUT116), .C2(KEYINPUT57), .ZN(new_n1102));
  NAND2_X1  g677(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1102), .B(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1105), .B(KEYINPUT117), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT61), .ZN(new_n1107));
  AND2_X1   g682(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  XOR2_X1   g684(.A(KEYINPUT58), .B(G1341), .Z(new_n1110));
  NAND2_X1  g685(.A1(new_n986), .A2(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1111), .B(KEYINPUT119), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT118), .B(G1996), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n976), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n610), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  XOR2_X1   g690(.A(new_n1115), .B(KEYINPUT59), .Z(new_n1116));
  OAI21_X1  g691(.A(new_n1107), .B1(new_n1108), .B2(new_n1105), .ZN(new_n1117));
  INV_X1    g692(.A(G1348), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n982), .A2(new_n1118), .B1(new_n1009), .B2(new_n782), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT60), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1119), .A2(new_n1120), .A3(new_n598), .A4(new_n594), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1119), .A2(new_n599), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1119), .A2(new_n599), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT60), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1116), .A2(new_n1117), .A3(new_n1121), .A4(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1106), .A2(new_n1123), .ZN(new_n1126));
  OAI22_X1  g701(.A1(new_n1109), .A2(new_n1125), .B1(new_n1126), .B2(new_n1108), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1071), .B1(new_n1097), .B2(new_n1127), .ZN(new_n1128));
  XOR2_X1   g703(.A(G290), .B(G1986), .Z(new_n1129));
  OAI21_X1  g704(.A(new_n946), .B1(new_n937), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n959), .B1(new_n1128), .B2(new_n1130), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g706(.A1(new_n657), .A2(G319), .ZN(new_n1133));
  XNOR2_X1  g707(.A(new_n1133), .B(KEYINPUT125), .ZN(new_n1134));
  NAND3_X1  g708(.A1(new_n644), .A2(KEYINPUT126), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g709(.A(new_n1135), .ZN(new_n1136));
  AOI21_X1  g710(.A(KEYINPUT126), .B1(new_n644), .B2(new_n1134), .ZN(new_n1137));
  OAI21_X1  g711(.A(new_n678), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  AOI22_X1  g712(.A1(new_n918), .A2(new_n920), .B1(KEYINPUT127), .B2(new_n1138), .ZN(new_n1139));
  OR2_X1    g713(.A1(new_n1138), .A2(KEYINPUT127), .ZN(new_n1140));
  OAI211_X1 g714(.A(new_n1139), .B(new_n1140), .C1(new_n859), .C2(new_n860), .ZN(G225));
  INV_X1    g715(.A(G225), .ZN(G308));
endmodule


