//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1 0 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 0 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  NAND4_X1  g005(.A1(new_n189), .A2(new_n191), .A3(KEYINPUT0), .A4(G128), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n190), .A2(G146), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n188), .A2(G143), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT0), .B(G128), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n192), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G137), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(KEYINPUT11), .A3(G134), .ZN(new_n199));
  INV_X1    g013(.A(G134), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G137), .ZN(new_n201));
  AND2_X1   g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT64), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n198), .A2(G134), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT11), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  AOI211_X1 g020(.A(KEYINPUT64), .B(KEYINPUT11), .C1(new_n198), .C2(G134), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n202), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G131), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n205), .B1(new_n200), .B2(G137), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT64), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n204), .A2(new_n203), .A3(new_n205), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G131), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(new_n202), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n197), .B1(new_n209), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n199), .A2(new_n201), .ZN(new_n217));
  AOI211_X1 g031(.A(G131), .B(new_n217), .C1(new_n211), .C2(new_n212), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT1), .B1(new_n190), .B2(G146), .ZN(new_n219));
  OAI211_X1 g033(.A(G128), .B(new_n219), .C1(new_n193), .C2(new_n194), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n204), .A2(new_n201), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G131), .ZN(new_n222));
  INV_X1    g036(.A(G128), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n189), .B(new_n191), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n220), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n218), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT2), .ZN(new_n228));
  INV_X1    g042(.A(G113), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(KEYINPUT68), .A2(KEYINPUT2), .A3(G113), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n228), .A2(new_n229), .A3(KEYINPUT67), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n234), .B1(KEYINPUT2), .B2(G113), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n232), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G119), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT69), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G119), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n239), .A2(new_n241), .A3(G116), .ZN(new_n242));
  INV_X1    g056(.A(G116), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G119), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n237), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n232), .A2(new_n236), .A3(new_n242), .A4(new_n244), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NOR3_X1   g062(.A1(new_n216), .A2(new_n226), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT28), .ZN(new_n250));
  INV_X1    g064(.A(new_n197), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n214), .B1(new_n213), .B2(new_n202), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n251), .B1(new_n218), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n248), .ZN(new_n254));
  AND3_X1   g068(.A1(new_n220), .A2(new_n222), .A3(new_n224), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(new_n215), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n253), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT28), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT66), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n260), .B1(new_n218), .B2(new_n225), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n255), .A2(KEYINPUT66), .A3(new_n215), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT65), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n253), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n216), .A2(KEYINPUT65), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n263), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n250), .B(new_n259), .C1(new_n267), .C2(new_n254), .ZN(new_n268));
  INV_X1    g082(.A(G237), .ZN(new_n269));
  INV_X1    g083(.A(G953), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(new_n270), .A3(G210), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n271), .B(KEYINPUT27), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT26), .B(G101), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n272), .B(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n274), .B(KEYINPUT70), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n268), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT30), .ZN(new_n277));
  NOR3_X1   g091(.A1(new_n216), .A2(new_n226), .A3(new_n277), .ZN(new_n278));
  NOR3_X1   g092(.A1(new_n218), .A2(new_n260), .A3(new_n225), .ZN(new_n279));
  AOI21_X1  g093(.A(KEYINPUT66), .B1(new_n255), .B2(new_n215), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n216), .A2(KEYINPUT65), .ZN(new_n282));
  AOI211_X1 g096(.A(new_n264), .B(new_n197), .C1(new_n209), .C2(new_n215), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n278), .B1(new_n284), .B2(new_n277), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n249), .B1(new_n285), .B2(new_n248), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT31), .B1(new_n286), .B2(new_n274), .ZN(new_n287));
  INV_X1    g101(.A(new_n278), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n248), .B(new_n288), .C1(new_n267), .C2(KEYINPUT30), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n289), .A2(KEYINPUT31), .A3(new_n274), .A4(new_n257), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n276), .B1(new_n287), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(G472), .A2(G902), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n293), .B(KEYINPUT71), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n292), .A2(KEYINPUT32), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT32), .ZN(new_n297));
  INV_X1    g111(.A(new_n276), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n289), .A2(new_n274), .A3(new_n257), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT31), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n298), .B1(new_n301), .B2(new_n290), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n297), .B1(new_n302), .B2(new_n294), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n296), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT72), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n254), .B1(new_n253), .B2(new_n256), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n305), .B(KEYINPUT28), .C1(new_n249), .C2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n259), .A2(KEYINPUT72), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n248), .B1(new_n216), .B2(new_n226), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n258), .B1(new_n309), .B2(new_n257), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n307), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n274), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT29), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(G902), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n313), .B1(new_n268), .B2(new_n275), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n274), .B1(new_n289), .B2(new_n257), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT73), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n318), .A2(new_n319), .A3(G472), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n319), .B1(new_n318), .B2(G472), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n187), .B1(new_n304), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n318), .A2(G472), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT73), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n318), .A2(new_n319), .A3(G472), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n327), .A2(KEYINPUT74), .A3(new_n303), .A4(new_n296), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT82), .ZN(new_n330));
  INV_X1    g144(.A(G140), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G125), .ZN(new_n332));
  INV_X1    g146(.A(G125), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G140), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n332), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n331), .A2(KEYINPUT76), .A3(G125), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(KEYINPUT16), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT16), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n332), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n188), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT77), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n338), .A2(new_n340), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G146), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n338), .A2(KEYINPUT77), .A3(new_n188), .A4(new_n340), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n343), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n238), .A2(G128), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT69), .B(G119), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n348), .B1(new_n349), .B2(G128), .ZN(new_n350));
  XOR2_X1   g164(.A(KEYINPUT24), .B(G110), .Z(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT23), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n239), .A2(new_n241), .A3(G128), .ZN(new_n354));
  INV_X1    g168(.A(new_n348), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n239), .A2(new_n241), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT23), .B1(new_n357), .B2(new_n223), .ZN(new_n358));
  OAI21_X1  g172(.A(KEYINPUT75), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT75), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n353), .B1(new_n349), .B2(G128), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n360), .B(new_n361), .C1(new_n350), .C2(new_n353), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n359), .A2(new_n362), .A3(G110), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n347), .A2(new_n352), .A3(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT78), .B(G110), .ZN(new_n365));
  NOR3_X1   g179(.A1(new_n356), .A2(new_n358), .A3(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n350), .A2(new_n351), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT79), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OR2_X1    g182(.A1(new_n350), .A2(new_n351), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT79), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n361), .B1(new_n350), .B2(new_n353), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n369), .B(new_n370), .C1(new_n371), .C2(new_n365), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n332), .A2(new_n334), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n373), .A2(new_n188), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n374), .B1(new_n344), .B2(G146), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n368), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(KEYINPUT22), .B(G137), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n270), .A2(G221), .A3(G234), .ZN(new_n378));
  XOR2_X1   g192(.A(new_n377), .B(new_n378), .Z(new_n379));
  NAND3_X1  g193(.A1(new_n364), .A2(new_n376), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT80), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT80), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n364), .A2(new_n376), .A3(new_n382), .A4(new_n379), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n364), .A2(new_n376), .ZN(new_n385));
  INV_X1    g199(.A(new_n379), .ZN(new_n386));
  AOI21_X1  g200(.A(G902), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n384), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n389), .B1(new_n384), .B2(new_n387), .ZN(new_n391));
  NAND2_X1  g205(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NOR3_X1   g207(.A1(new_n390), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G217), .ZN(new_n395));
  INV_X1    g209(.A(G902), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n395), .B1(G234), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n330), .B1(new_n394), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n391), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n384), .A2(new_n387), .A3(new_n389), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n400), .A2(new_n401), .A3(new_n392), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(KEYINPUT82), .A3(new_n397), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n385), .A2(new_n386), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n384), .A2(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n397), .A2(G902), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n399), .A2(new_n403), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT20), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n269), .A2(new_n270), .A3(G214), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(new_n190), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(KEYINPUT17), .A3(G131), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n343), .A2(new_n345), .A3(new_n346), .A4(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT17), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n411), .B(G143), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(G131), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n414), .A2(KEYINPUT91), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n345), .A2(new_n346), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT91), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n419), .A2(new_n420), .A3(new_n343), .A4(new_n413), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(G113), .B(G122), .ZN(new_n423));
  INV_X1    g237(.A(G104), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n423), .B(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(KEYINPUT18), .A2(G131), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n416), .B(new_n426), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n336), .A2(new_n337), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n374), .B1(new_n428), .B2(G146), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n422), .A2(new_n425), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n417), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT19), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n373), .A2(KEYINPUT90), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT90), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n428), .B1(new_n436), .B2(new_n373), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n435), .B1(new_n437), .B2(new_n434), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n433), .B(new_n345), .C1(new_n438), .C2(G146), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n431), .ZN(new_n440));
  INV_X1    g254(.A(new_n425), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n432), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(G475), .A2(G902), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n410), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n444), .ZN(new_n446));
  AOI211_X1 g260(.A(KEYINPUT20), .B(new_n446), .C1(new_n432), .C2(new_n442), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n422), .A2(new_n431), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n441), .ZN(new_n449));
  AOI21_X1  g263(.A(G902), .B1(new_n449), .B2(new_n432), .ZN(new_n450));
  INV_X1    g264(.A(G475), .ZN(new_n451));
  OAI22_X1  g265(.A1(new_n445), .A2(new_n447), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  XOR2_X1   g266(.A(G128), .B(G143), .Z(new_n453));
  INV_X1    g267(.A(KEYINPUT93), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(G128), .B(G143), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT93), .ZN(new_n457));
  AOI21_X1  g271(.A(G134), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT13), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(new_n190), .A3(G128), .ZN(new_n461));
  OAI211_X1 g275(.A(G134), .B(new_n461), .C1(new_n453), .C2(new_n460), .ZN(new_n462));
  INV_X1    g276(.A(G107), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT92), .ZN(new_n464));
  INV_X1    g278(.A(G122), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n464), .B1(new_n465), .B2(G116), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n243), .A2(KEYINPUT92), .A3(G122), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n465), .A2(G116), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n463), .A3(new_n469), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n459), .B(new_n462), .C1(new_n470), .C2(new_n472), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n468), .A2(KEYINPUT14), .B1(G116), .B2(new_n465), .ZN(new_n474));
  OR2_X1    g288(.A1(new_n474), .A2(KEYINPUT95), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n468), .A2(KEYINPUT14), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n476), .B1(new_n474), .B2(KEYINPUT95), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n463), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  OR2_X1    g292(.A1(new_n471), .A2(KEYINPUT94), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n471), .A2(KEYINPUT94), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n455), .A2(G134), .A3(new_n457), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n479), .B(new_n480), .C1(new_n481), .C2(new_n458), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n473), .B1(new_n478), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT9), .B(G234), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n484), .A2(new_n395), .A3(G953), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n485), .B(KEYINPUT96), .Z(new_n486));
  NAND2_X1  g300(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT97), .ZN(new_n488));
  INV_X1    g302(.A(new_n486), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n489), .B(new_n473), .C1(new_n478), .C2(new_n482), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n487), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  OR3_X1    g305(.A1(new_n483), .A2(new_n488), .A3(new_n486), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(new_n492), .A3(new_n396), .ZN(new_n493));
  INV_X1    g307(.A(G478), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n494), .A2(KEYINPUT15), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n493), .B(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G952), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n497), .A2(G953), .ZN(new_n498));
  INV_X1    g312(.A(G234), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n498), .B1(new_n499), .B2(new_n269), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  AOI211_X1 g315(.A(new_n396), .B(new_n270), .C1(G234), .C2(G237), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT21), .B(G898), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n452), .A2(new_n496), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n424), .A2(G107), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n463), .A2(KEYINPUT3), .A3(G104), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT3), .B1(new_n463), .B2(G104), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT4), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n510), .A3(G101), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n509), .A2(G101), .ZN(new_n512));
  INV_X1    g326(.A(G101), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n513), .B(new_n506), .C1(new_n507), .C2(new_n508), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(KEYINPUT4), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n248), .B(new_n511), .C1(new_n512), .C2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT84), .B1(new_n463), .B2(G104), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT84), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(new_n424), .A3(G107), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n463), .A2(G104), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n517), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(G101), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n522), .A2(new_n514), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n242), .A2(KEYINPUT5), .A3(new_n244), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT5), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n349), .A2(new_n525), .A3(G116), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n524), .A2(G113), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n523), .A2(new_n247), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n516), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(G110), .B(G122), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n516), .A2(new_n528), .A3(new_n530), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n532), .A2(KEYINPUT6), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n220), .A2(new_n224), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n333), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n251), .A2(G125), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(G224), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n540), .A2(G953), .ZN(new_n541));
  XOR2_X1   g355(.A(new_n539), .B(new_n541), .Z(new_n542));
  INV_X1    g356(.A(KEYINPUT6), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n529), .A2(new_n543), .A3(new_n531), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n534), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n545), .A2(new_n396), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT89), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT88), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n537), .B(new_n538), .C1(new_n548), .C2(new_n541), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT7), .B1(new_n540), .B2(G953), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n549), .B(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT87), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT86), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n242), .A2(KEYINPUT5), .A3(new_n244), .ZN(new_n554));
  OAI21_X1  g368(.A(G113), .B1(new_n242), .B2(KEYINPUT5), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n247), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n522), .A2(new_n514), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n553), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n557), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n556), .A2(new_n553), .A3(new_n557), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n530), .B(KEYINPUT8), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n552), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n563), .ZN(new_n565));
  AOI211_X1 g379(.A(KEYINPUT87), .B(new_n565), .C1(new_n560), .C2(new_n561), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n547), .B(new_n551), .C1(new_n564), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n533), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n527), .A2(new_n247), .B1(new_n514), .B2(new_n522), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n569), .B1(new_n528), .B2(new_n553), .ZN(new_n570));
  INV_X1    g384(.A(new_n561), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n563), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT87), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n562), .A2(new_n552), .A3(new_n563), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n547), .B1(new_n575), .B2(new_n551), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n546), .B1(new_n568), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(G210), .B1(G237), .B2(G902), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n578), .B(new_n546), .C1(new_n568), .C2(new_n576), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(G214), .B1(G237), .B2(G902), .ZN(new_n583));
  OAI21_X1  g397(.A(G221), .B1(new_n484), .B2(G902), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n522), .A2(new_n514), .A3(new_n224), .A4(new_n220), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(KEYINPUT10), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT85), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n218), .A2(new_n252), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n251), .B(new_n511), .C1(new_n512), .C2(new_n515), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n587), .A2(new_n588), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n523), .A2(KEYINPUT10), .A3(new_n536), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT10), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n586), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n592), .A2(new_n590), .A3(new_n589), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(KEYINPUT85), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n209), .A2(new_n215), .ZN(new_n598));
  INV_X1    g412(.A(new_n586), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n522), .A2(new_n514), .B1(new_n224), .B2(new_n220), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT12), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n597), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(G110), .B(G140), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n270), .A2(G227), .ZN(new_n606));
  XOR2_X1   g420(.A(new_n605), .B(new_n606), .Z(new_n607));
  XOR2_X1   g421(.A(new_n607), .B(KEYINPUT83), .Z(new_n608));
  AOI21_X1  g422(.A(new_n607), .B1(new_n591), .B2(new_n596), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n587), .A2(new_n590), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n598), .ZN(new_n611));
  AOI22_X1  g425(.A1(new_n604), .A2(new_n608), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(G469), .B1(new_n612), .B2(G902), .ZN(new_n613));
  INV_X1    g427(.A(G469), .ZN(new_n614));
  INV_X1    g428(.A(new_n607), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n597), .A2(new_n615), .A3(new_n603), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n615), .B1(new_n597), .B2(new_n611), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n614), .B(new_n396), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n585), .B1(new_n613), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n582), .A2(new_n583), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n329), .A2(new_n409), .A3(new_n505), .A4(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT98), .B(G101), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G3));
  INV_X1    g438(.A(KEYINPUT99), .ZN(new_n625));
  INV_X1    g439(.A(new_n581), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n551), .B1(new_n564), .B2(new_n566), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(KEYINPUT89), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n628), .A2(new_n533), .A3(new_n567), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n578), .B1(new_n629), .B2(new_n546), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n583), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n625), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n582), .A2(KEYINPUT99), .A3(new_n583), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n504), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n425), .B1(new_n439), .B2(new_n431), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n430), .B1(new_n418), .B2(new_n421), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n636), .B1(new_n425), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(KEYINPUT20), .B1(new_n638), .B2(new_n446), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n443), .A2(new_n410), .A3(new_n444), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n432), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n637), .A2(new_n425), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n396), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(G475), .ZN(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT100), .B(G478), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n493), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT33), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n491), .A2(new_n492), .A3(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n487), .A2(KEYINPUT33), .A3(new_n490), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n649), .A2(G478), .A3(new_n396), .A4(new_n650), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n641), .A2(new_n645), .B1(new_n647), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g466(.A(G472), .B1(new_n302), .B2(G902), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n292), .A2(new_n295), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n653), .A2(new_n654), .A3(new_n619), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n408), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n635), .A2(new_n652), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n657), .B(KEYINPUT101), .Z(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT34), .B(G104), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G6));
  INV_X1    g474(.A(new_n495), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n493), .B(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n452), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n635), .A2(new_n656), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT35), .B(G107), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  XNOR2_X1  g480(.A(new_n385), .B(KEYINPUT102), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n386), .A2(KEYINPUT36), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n667), .B(new_n668), .Z(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n406), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n399), .A2(new_n403), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n505), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n653), .A2(new_n654), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n620), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT103), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT37), .B(G110), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G12));
  NAND2_X1  g493(.A1(new_n633), .A2(new_n634), .ZN(new_n680));
  AOI22_X1  g494(.A1(new_n640), .A2(new_n639), .B1(new_n644), .B2(G475), .ZN(new_n681));
  INV_X1    g495(.A(G900), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n502), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n500), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n681), .A2(new_n496), .A3(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n671), .A2(new_n619), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n329), .A2(new_n680), .A3(new_n686), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G128), .ZN(G30));
  NOR2_X1   g504(.A1(new_n681), .A2(new_n662), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n684), .B(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n619), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n691), .B1(new_n695), .B2(KEYINPUT40), .ZN(new_n696));
  AOI211_X1 g510(.A(new_n632), .B(new_n696), .C1(KEYINPUT40), .C2(new_n695), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n582), .B(KEYINPUT38), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n309), .A2(new_n257), .ZN(new_n699));
  AOI22_X1  g513(.A1(new_n286), .A2(new_n274), .B1(new_n275), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g514(.A(G472), .B1(new_n700), .B2(G902), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n296), .A2(new_n701), .A3(new_n303), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n671), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n697), .A2(new_n698), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G143), .ZN(G45));
  NAND2_X1  g520(.A1(new_n651), .A2(new_n647), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n452), .A2(new_n707), .A3(new_n684), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n329), .A2(new_n680), .A3(new_n688), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G146), .ZN(G48));
  AOI21_X1  g525(.A(new_n408), .B1(new_n323), .B2(new_n328), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n616), .A2(new_n617), .ZN(new_n713));
  OAI21_X1  g527(.A(G469), .B1(new_n713), .B2(G902), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n714), .A2(new_n584), .A3(new_n618), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n712), .A2(new_n635), .A3(new_n652), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT41), .B(G113), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  NAND4_X1  g532(.A1(new_n712), .A2(new_n635), .A3(new_n663), .A4(new_n715), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G116), .ZN(G18));
  AOI21_X1  g534(.A(new_n672), .B1(new_n323), .B2(new_n328), .ZN(new_n721));
  INV_X1    g535(.A(new_n715), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n633), .B2(new_n634), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G119), .ZN(G21));
  NAND2_X1  g539(.A1(new_n691), .A2(new_n715), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n301), .A2(new_n290), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n307), .B(new_n275), .C1(new_n308), .C2(new_n310), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n295), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n653), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n408), .A2(new_n726), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n635), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G122), .ZN(G24));
  AND2_X1   g548(.A1(new_n730), .A2(new_n653), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n671), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(new_n708), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n723), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  NAND3_X1  g553(.A1(new_n654), .A2(KEYINPUT108), .A3(new_n297), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT108), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n303), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT107), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n296), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n740), .A2(new_n742), .A3(new_n744), .A4(new_n296), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n327), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n580), .A2(new_n583), .A3(new_n581), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n609), .A2(new_n611), .ZN(new_n750));
  INV_X1    g564(.A(new_n604), .ZN(new_n751));
  INV_X1    g565(.A(new_n608), .ZN(new_n752));
  OAI211_X1 g566(.A(G469), .B(new_n750), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(G469), .A2(G902), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n618), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n755), .A2(KEYINPUT105), .A3(new_n584), .ZN(new_n756));
  AOI21_X1  g570(.A(KEYINPUT105), .B1(new_n755), .B2(new_n584), .ZN(new_n757));
  NOR4_X1   g571(.A1(new_n749), .A2(new_n756), .A3(new_n757), .A4(new_n708), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n748), .A2(KEYINPUT42), .A3(new_n409), .A4(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n329), .A2(KEYINPUT106), .A3(new_n758), .A4(new_n409), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT42), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(KEYINPUT106), .B1(new_n712), .B2(new_n758), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n759), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G131), .ZN(G33));
  NOR4_X1   g579(.A1(new_n749), .A2(new_n756), .A3(new_n685), .A4(new_n757), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n329), .A2(new_n409), .A3(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G134), .ZN(G36));
  INV_X1    g582(.A(KEYINPUT43), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n769), .A2(KEYINPUT109), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n771), .B1(new_n681), .B2(new_n707), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n681), .A2(new_n707), .ZN(new_n773));
  XNOR2_X1  g587(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(new_n674), .A3(new_n671), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT44), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT112), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n775), .A2(KEYINPUT44), .A3(new_n674), .A4(new_n671), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT110), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n749), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n783), .B1(new_n780), .B2(KEYINPUT110), .ZN(new_n784));
  OAI21_X1  g598(.A(KEYINPUT111), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n780), .A2(KEYINPUT110), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT111), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n786), .A2(new_n787), .A3(new_n783), .A4(new_n781), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n779), .A2(new_n785), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT45), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n612), .A2(KEYINPUT45), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(G469), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT46), .B1(new_n796), .B2(new_n754), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n713), .A2(G469), .A3(G902), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n796), .A2(KEYINPUT46), .A3(new_n754), .ZN(new_n800));
  AOI211_X1 g614(.A(new_n585), .B(new_n693), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n779), .A2(new_n785), .A3(new_n788), .A4(KEYINPUT113), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n791), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G137), .ZN(G39));
  INV_X1    g618(.A(new_n329), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n805), .A2(new_n408), .A3(new_n709), .A4(new_n783), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n799), .A2(new_n800), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT47), .B1(new_n807), .B2(new_n584), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT47), .ZN(new_n809));
  AOI211_X1 g623(.A(new_n809), .B(new_n585), .C1(new_n799), .C2(new_n800), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n806), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(new_n331), .ZN(G42));
  NOR2_X1   g627(.A1(new_n698), .A2(new_n702), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n714), .A2(new_n618), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT49), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n583), .B(new_n584), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n817), .B1(new_n816), .B2(new_n815), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n814), .A2(new_n409), .A3(new_n773), .A4(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n394), .A2(new_n330), .A3(new_n398), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT82), .B1(new_n402), .B2(new_n397), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n822), .A2(KEYINPUT116), .A3(new_n670), .A4(new_n684), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n824));
  INV_X1    g638(.A(new_n684), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n824), .B1(new_n671), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n691), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n828), .B1(new_n633), .B2(new_n634), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n702), .A2(new_n619), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n827), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n689), .A3(new_n710), .A4(new_n738), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT52), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n832), .B(new_n833), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n721), .A2(new_n723), .B1(new_n635), .B2(new_n732), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n835), .A2(new_n716), .A3(new_n719), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n836), .A2(new_n764), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT114), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n452), .A2(new_n496), .A3(new_n825), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n631), .A2(new_n838), .A3(new_n839), .A4(new_n583), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n681), .A2(new_n662), .A3(new_n684), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT114), .B1(new_n749), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n329), .A2(new_n688), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT115), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n687), .B1(new_n323), .B2(new_n328), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT115), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(new_n847), .A3(new_n843), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n504), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n582), .A2(new_n850), .A3(new_n583), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n663), .A2(new_n652), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n673), .A2(new_n675), .B1(new_n853), .B2(new_n656), .ZN(new_n854));
  INV_X1    g668(.A(new_n736), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n758), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n622), .A2(new_n854), .A3(new_n767), .A4(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n849), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n689), .A2(new_n738), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n859), .B1(new_n860), .B2(new_n833), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n834), .A2(new_n837), .A3(new_n858), .A4(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n858), .A2(new_n764), .A3(new_n836), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n860), .A2(new_n833), .A3(new_n710), .A4(new_n831), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n832), .A2(KEYINPUT52), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n859), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT54), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n689), .A2(new_n738), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n859), .B1(new_n870), .B2(KEYINPUT52), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n836), .A2(new_n764), .A3(new_n871), .ZN(new_n872));
  AND4_X1   g686(.A1(new_n622), .A2(new_n854), .A3(new_n767), .A4(new_n856), .ZN(new_n873));
  AND4_X1   g687(.A1(new_n847), .A2(new_n329), .A3(new_n688), .A4(new_n843), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n847), .B1(new_n846), .B2(new_n843), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n873), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT117), .B1(new_n849), .B2(new_n857), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n872), .A2(new_n880), .A3(new_n834), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT54), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n881), .A2(new_n867), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n869), .A2(new_n883), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n775), .A2(new_n501), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(new_n409), .A3(new_n735), .ZN(new_n886));
  NOR4_X1   g700(.A1(new_n886), .A2(new_n583), .A3(new_n698), .A4(new_n722), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT50), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n886), .A2(new_n749), .ZN(new_n889));
  INV_X1    g703(.A(new_n811), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n815), .A2(new_n585), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n722), .A2(new_n749), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n409), .A2(new_n893), .A3(new_n703), .A4(new_n501), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n894), .A2(new_n452), .A3(new_n707), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n885), .A2(new_n893), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n895), .B1(new_n855), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n888), .A2(new_n892), .A3(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT51), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n898), .A2(new_n899), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n748), .A2(new_n409), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n896), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT48), .ZN(new_n904));
  INV_X1    g718(.A(new_n652), .ZN(new_n905));
  INV_X1    g719(.A(new_n723), .ZN(new_n906));
  OAI221_X1 g720(.A(new_n498), .B1(new_n905), .B2(new_n894), .C1(new_n886), .C2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n901), .A2(new_n904), .A3(new_n908), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n884), .A2(new_n900), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n497), .A2(new_n270), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT118), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n819), .B1(new_n910), .B2(new_n912), .ZN(G75));
  NOR2_X1   g727(.A1(new_n270), .A2(G952), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n396), .B1(new_n881), .B2(new_n867), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT56), .B1(new_n916), .B2(G210), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n534), .A2(new_n544), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(new_n542), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT55), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n915), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n917), .B2(new_n920), .ZN(G51));
  INV_X1    g736(.A(KEYINPUT119), .ZN(new_n923));
  AOI211_X1 g737(.A(new_n396), .B(new_n796), .C1(new_n881), .C2(new_n867), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n754), .B(KEYINPUT57), .Z(new_n925));
  AND3_X1   g739(.A1(new_n881), .A2(new_n867), .A3(new_n882), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n882), .B1(new_n881), .B2(new_n867), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n713), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n924), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n923), .B1(new_n930), .B2(new_n914), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n881), .A2(new_n867), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(KEYINPUT54), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n883), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n713), .B1(new_n934), .B2(new_n925), .ZN(new_n935));
  OAI211_X1 g749(.A(KEYINPUT119), .B(new_n915), .C1(new_n935), .C2(new_n924), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n931), .A2(new_n936), .ZN(G54));
  AND2_X1   g751(.A1(KEYINPUT58), .A2(G475), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n916), .A2(new_n443), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n443), .B1(new_n916), .B2(new_n938), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n939), .A2(new_n940), .A3(new_n914), .ZN(G60));
  INV_X1    g755(.A(KEYINPUT120), .ZN(new_n942));
  NAND2_X1  g756(.A1(G478), .A2(G902), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT59), .Z(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n869), .B2(new_n883), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n649), .A2(new_n650), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n946), .A2(new_n944), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(new_n926), .B2(new_n927), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n915), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n942), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n914), .B1(new_n934), .B2(new_n949), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n953), .B(KEYINPUT120), .C1(new_n947), .C2(new_n945), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n952), .A2(new_n954), .ZN(G63));
  NAND2_X1  g769(.A1(G217), .A2(G902), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT60), .Z(new_n957));
  NAND2_X1  g771(.A1(new_n932), .A2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n405), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n914), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT61), .B1(new_n960), .B2(KEYINPUT121), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n932), .A2(new_n669), .A3(new_n957), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n960), .B(new_n962), .C1(KEYINPUT121), .C2(KEYINPUT61), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(G66));
  OAI21_X1  g780(.A(G953), .B1(new_n503), .B2(new_n540), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n836), .A2(new_n622), .A3(new_n854), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n967), .B1(new_n968), .B2(G953), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n918), .B1(G898), .B2(new_n270), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(G69));
  INV_X1    g785(.A(KEYINPUT125), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n860), .A2(new_n710), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n767), .B1(new_n806), .B2(new_n811), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n801), .A2(new_n748), .A3(new_n409), .A4(new_n829), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT124), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n976), .B(new_n977), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n975), .A2(new_n978), .A3(new_n764), .ZN(new_n979));
  AOI21_X1  g793(.A(G953), .B1(new_n979), .B2(new_n803), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n270), .A2(G900), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n972), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n981), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n975), .A2(new_n978), .A3(new_n764), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n802), .A2(new_n801), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n984), .B1(new_n985), .B2(new_n791), .ZN(new_n986));
  OAI211_X1 g800(.A(KEYINPUT125), .B(new_n983), .C1(new_n986), .C2(G953), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n285), .B(new_n438), .Z(new_n988));
  NAND3_X1  g802(.A1(new_n982), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n852), .A2(new_n695), .A3(new_n749), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n712), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n991), .B1(new_n806), .B2(new_n811), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n860), .A2(new_n705), .A3(new_n710), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n992), .B1(new_n993), .B2(KEYINPUT62), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT62), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n860), .A2(new_n705), .A3(new_n995), .A4(new_n710), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(G953), .B1(new_n997), .B2(new_n803), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n988), .B(KEYINPUT122), .ZN(new_n999));
  INV_X1    g813(.A(new_n999), .ZN(new_n1000));
  OAI21_X1  g814(.A(KEYINPUT123), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT123), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n994), .A2(new_n996), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1003), .B1(new_n985), .B2(new_n791), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n1002), .B(new_n999), .C1(new_n1004), .C2(G953), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n270), .B1(G227), .B2(G900), .ZN(new_n1007));
  AND3_X1   g821(.A1(new_n989), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1007), .B1(new_n989), .B2(new_n1006), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1008), .A2(new_n1009), .ZN(G72));
  NAND2_X1  g824(.A1(G472), .A2(G902), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1011), .B(KEYINPUT127), .ZN(new_n1012));
  XNOR2_X1  g826(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1014), .B1(new_n1004), .B2(new_n968), .ZN(new_n1015));
  OR3_X1    g829(.A1(new_n1015), .A2(new_n312), .A3(new_n286), .ZN(new_n1016));
  AND2_X1   g830(.A1(new_n986), .A2(new_n968), .ZN(new_n1017));
  OAI211_X1 g831(.A(new_n312), .B(new_n286), .C1(new_n1017), .C2(new_n1014), .ZN(new_n1018));
  INV_X1    g832(.A(new_n317), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1014), .B1(new_n1019), .B2(new_n299), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n914), .B1(new_n868), .B2(new_n1020), .ZN(new_n1021));
  AND3_X1   g835(.A1(new_n1016), .A2(new_n1018), .A3(new_n1021), .ZN(G57));
endmodule


