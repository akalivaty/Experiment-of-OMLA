

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U325 ( .A(n420), .B(n419), .ZN(n545) );
  XNOR2_X1 U326 ( .A(n471), .B(KEYINPUT105), .ZN(n472) );
  INV_X1 U327 ( .A(KEYINPUT37), .ZN(n471) );
  XNOR2_X1 U328 ( .A(n348), .B(n293), .ZN(n349) );
  XNOR2_X1 U329 ( .A(n317), .B(n316), .ZN(n527) );
  XNOR2_X1 U330 ( .A(n429), .B(n428), .ZN(n517) );
  AND2_X1 U331 ( .A1(G232GAT), .A2(G233GAT), .ZN(n293) );
  XOR2_X1 U332 ( .A(G85GAT), .B(KEYINPUT76), .Z(n294) );
  AND2_X1 U333 ( .A1(G226GAT), .A2(G233GAT), .ZN(n295) );
  NOR2_X1 U334 ( .A1(n545), .A2(n517), .ZN(n430) );
  NOR2_X1 U335 ( .A1(n544), .A2(n490), .ZN(n529) );
  XNOR2_X1 U336 ( .A(n421), .B(n295), .ZN(n422) );
  NOR2_X1 U337 ( .A1(n461), .A2(n567), .ZN(n450) );
  XNOR2_X1 U338 ( .A(n423), .B(n422), .ZN(n425) );
  XNOR2_X1 U339 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U340 ( .A(n473), .B(n472), .ZN(n514) );
  NOR2_X1 U341 ( .A1(n527), .A2(n451), .ZN(n563) );
  INV_X1 U342 ( .A(G43GAT), .ZN(n475) );
  XNOR2_X1 U343 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U344 ( .A(n475), .B(KEYINPUT40), .ZN(n476) );
  XNOR2_X1 U345 ( .A(n455), .B(n454), .ZN(G1349GAT) );
  XNOR2_X1 U346 ( .A(n477), .B(n476), .ZN(G1330GAT) );
  XOR2_X1 U347 ( .A(KEYINPUT20), .B(KEYINPUT88), .Z(n297) );
  XNOR2_X1 U348 ( .A(G190GAT), .B(G99GAT), .ZN(n296) );
  XNOR2_X1 U349 ( .A(n297), .B(n296), .ZN(n299) );
  XOR2_X1 U350 ( .A(G43GAT), .B(G134GAT), .Z(n298) );
  XNOR2_X1 U351 ( .A(n299), .B(n298), .ZN(n315) );
  XOR2_X1 U352 ( .A(G127GAT), .B(KEYINPUT90), .Z(n301) );
  XNOR2_X1 U353 ( .A(G176GAT), .B(KEYINPUT86), .ZN(n300) );
  XNOR2_X1 U354 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U355 ( .A(KEYINPUT85), .B(KEYINPUT89), .Z(n303) );
  XNOR2_X1 U356 ( .A(G169GAT), .B(G15GAT), .ZN(n302) );
  XNOR2_X1 U357 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n305), .B(n304), .ZN(n313) );
  XNOR2_X1 U359 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n306) );
  XNOR2_X1 U360 ( .A(n306), .B(KEYINPUT84), .ZN(n444) );
  XOR2_X1 U361 ( .A(G71GAT), .B(n444), .Z(n311) );
  XOR2_X1 U362 ( .A(KEYINPUT87), .B(KEYINPUT19), .Z(n308) );
  XNOR2_X1 U363 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n307) );
  XNOR2_X1 U364 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U365 ( .A(KEYINPUT18), .B(n309), .Z(n426) );
  XNOR2_X1 U366 ( .A(n426), .B(G120GAT), .ZN(n310) );
  XNOR2_X1 U367 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U368 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U369 ( .A(n315), .B(n314), .ZN(n317) );
  NAND2_X1 U370 ( .A1(G227GAT), .A2(G233GAT), .ZN(n316) );
  XOR2_X1 U371 ( .A(KEYINPUT2), .B(KEYINPUT91), .Z(n319) );
  XNOR2_X1 U372 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n318) );
  XNOR2_X1 U373 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U374 ( .A(G141GAT), .B(n320), .Z(n436) );
  XOR2_X1 U375 ( .A(KEYINPUT24), .B(KEYINPUT92), .Z(n322) );
  XNOR2_X1 U376 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n321) );
  XNOR2_X1 U377 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U378 ( .A(G106GAT), .B(G218GAT), .Z(n324) );
  XOR2_X1 U379 ( .A(G50GAT), .B(G162GAT), .Z(n345) );
  XOR2_X1 U380 ( .A(KEYINPUT72), .B(G78GAT), .Z(n381) );
  XNOR2_X1 U381 ( .A(n345), .B(n381), .ZN(n323) );
  XNOR2_X1 U382 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U383 ( .A(n326), .B(n325), .Z(n328) );
  NAND2_X1 U384 ( .A1(G228GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U385 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U386 ( .A(n329), .B(G148GAT), .Z(n333) );
  XOR2_X1 U387 ( .A(G204GAT), .B(G211GAT), .Z(n331) );
  XNOR2_X1 U388 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n424) );
  XNOR2_X1 U390 ( .A(G22GAT), .B(n424), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U392 ( .A(n436), .B(n334), .ZN(n461) );
  XOR2_X1 U393 ( .A(G92GAT), .B(KEYINPUT77), .Z(n336) );
  XNOR2_X1 U394 ( .A(G190GAT), .B(G218GAT), .ZN(n335) );
  XNOR2_X1 U395 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U396 ( .A(G36GAT), .B(n337), .Z(n423) );
  XOR2_X1 U397 ( .A(G43GAT), .B(KEYINPUT8), .Z(n339) );
  XNOR2_X1 U398 ( .A(KEYINPUT67), .B(KEYINPUT7), .ZN(n338) );
  XNOR2_X1 U399 ( .A(n339), .B(n338), .ZN(n364) );
  XNOR2_X1 U400 ( .A(G29GAT), .B(G134GAT), .ZN(n340) );
  XNOR2_X1 U401 ( .A(n294), .B(n340), .ZN(n443) );
  XNOR2_X1 U402 ( .A(n364), .B(n443), .ZN(n344) );
  XOR2_X1 U403 ( .A(KEYINPUT75), .B(KEYINPUT74), .Z(n342) );
  XNOR2_X1 U404 ( .A(KEYINPUT9), .B(KEYINPUT11), .ZN(n341) );
  XNOR2_X1 U405 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U406 ( .A(n344), .B(n343), .ZN(n350) );
  XOR2_X1 U407 ( .A(KEYINPUT78), .B(KEYINPUT10), .Z(n347) );
  XOR2_X1 U408 ( .A(G99GAT), .B(G106GAT), .Z(n371) );
  XNOR2_X1 U409 ( .A(n345), .B(n371), .ZN(n346) );
  XNOR2_X1 U410 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U411 ( .A(n423), .B(n351), .Z(n559) );
  INV_X1 U412 ( .A(n559), .ZN(n412) );
  XOR2_X1 U413 ( .A(G169GAT), .B(G8GAT), .Z(n427) );
  XOR2_X1 U414 ( .A(G197GAT), .B(G50GAT), .Z(n353) );
  XNOR2_X1 U415 ( .A(G29GAT), .B(G36GAT), .ZN(n352) );
  XNOR2_X1 U416 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U417 ( .A(n427), .B(n354), .Z(n356) );
  NAND2_X1 U418 ( .A1(G229GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U419 ( .A(n356), .B(n355), .ZN(n368) );
  XOR2_X1 U420 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n358) );
  XNOR2_X1 U421 ( .A(KEYINPUT69), .B(KEYINPUT29), .ZN(n357) );
  XNOR2_X1 U422 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U423 ( .A(KEYINPUT65), .B(G1GAT), .Z(n360) );
  XNOR2_X1 U424 ( .A(G141GAT), .B(G113GAT), .ZN(n359) );
  XNOR2_X1 U425 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U426 ( .A(n362), .B(n361), .Z(n366) );
  XNOR2_X1 U427 ( .A(G22GAT), .B(G15GAT), .ZN(n363) );
  XNOR2_X1 U428 ( .A(n363), .B(KEYINPUT68), .ZN(n397) );
  XNOR2_X1 U429 ( .A(n364), .B(n397), .ZN(n365) );
  XNOR2_X1 U430 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U431 ( .A(n368), .B(n367), .ZN(n548) );
  INV_X1 U432 ( .A(n548), .ZN(n569) );
  XNOR2_X1 U433 ( .A(G120GAT), .B(G148GAT), .ZN(n369) );
  XNOR2_X1 U434 ( .A(n369), .B(G57GAT), .ZN(n432) );
  XNOR2_X1 U435 ( .A(G71GAT), .B(KEYINPUT70), .ZN(n370) );
  XNOR2_X1 U436 ( .A(n370), .B(KEYINPUT13), .ZN(n401) );
  XNOR2_X1 U437 ( .A(n432), .B(n401), .ZN(n385) );
  XOR2_X1 U438 ( .A(G176GAT), .B(G64GAT), .Z(n421) );
  XOR2_X1 U439 ( .A(n371), .B(n421), .Z(n373) );
  NAND2_X1 U440 ( .A1(G230GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U441 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U442 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n375) );
  XNOR2_X1 U443 ( .A(KEYINPUT71), .B(KEYINPUT31), .ZN(n374) );
  XNOR2_X1 U444 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U445 ( .A(n377), .B(n376), .Z(n383) );
  XOR2_X1 U446 ( .A(KEYINPUT32), .B(G92GAT), .Z(n379) );
  XNOR2_X1 U447 ( .A(G204GAT), .B(G85GAT), .ZN(n378) );
  XNOR2_X1 U448 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U449 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U450 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U451 ( .A(n385), .B(n384), .Z(n573) );
  XOR2_X1 U452 ( .A(n573), .B(KEYINPUT41), .Z(n532) );
  NAND2_X1 U453 ( .A1(n569), .A2(n532), .ZN(n388) );
  XOR2_X1 U454 ( .A(KEYINPUT46), .B(KEYINPUT115), .Z(n386) );
  XNOR2_X1 U455 ( .A(KEYINPUT114), .B(n386), .ZN(n387) );
  XNOR2_X1 U456 ( .A(n388), .B(n387), .ZN(n408) );
  XOR2_X1 U457 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n390) );
  XNOR2_X1 U458 ( .A(KEYINPUT14), .B(KEYINPUT15), .ZN(n389) );
  XNOR2_X1 U459 ( .A(n390), .B(n389), .ZN(n407) );
  XOR2_X1 U460 ( .A(KEYINPUT83), .B(G64GAT), .Z(n392) );
  XNOR2_X1 U461 ( .A(G8GAT), .B(G57GAT), .ZN(n391) );
  XNOR2_X1 U462 ( .A(n392), .B(n391), .ZN(n396) );
  XOR2_X1 U463 ( .A(G78GAT), .B(G211GAT), .Z(n394) );
  XNOR2_X1 U464 ( .A(G183GAT), .B(G155GAT), .ZN(n393) );
  XNOR2_X1 U465 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U466 ( .A(n396), .B(n395), .ZN(n405) );
  XOR2_X1 U467 ( .A(G1GAT), .B(G127GAT), .Z(n431) );
  XOR2_X1 U468 ( .A(n431), .B(n397), .Z(n399) );
  NAND2_X1 U469 ( .A1(G231GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U470 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U471 ( .A(n400), .B(KEYINPUT80), .Z(n403) );
  XNOR2_X1 U472 ( .A(n401), .B(KEYINPUT12), .ZN(n402) );
  XNOR2_X1 U473 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U474 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U475 ( .A(n407), .B(n406), .Z(n578) );
  INV_X1 U476 ( .A(n578), .ZN(n555) );
  NAND2_X1 U477 ( .A1(n408), .A2(n555), .ZN(n409) );
  NOR2_X1 U478 ( .A1(n412), .A2(n409), .ZN(n411) );
  XNOR2_X1 U479 ( .A(KEYINPUT47), .B(KEYINPUT116), .ZN(n410) );
  XNOR2_X1 U480 ( .A(n411), .B(n410), .ZN(n418) );
  XOR2_X1 U481 ( .A(KEYINPUT79), .B(n412), .Z(n564) );
  XNOR2_X1 U482 ( .A(KEYINPUT36), .B(KEYINPUT104), .ZN(n413) );
  XNOR2_X1 U483 ( .A(n564), .B(n413), .ZN(n582) );
  NAND2_X1 U484 ( .A1(n582), .A2(n578), .ZN(n414) );
  XOR2_X1 U485 ( .A(KEYINPUT45), .B(n414), .Z(n416) );
  NOR2_X1 U486 ( .A1(n573), .A2(n569), .ZN(n415) );
  NAND2_X1 U487 ( .A1(n416), .A2(n415), .ZN(n417) );
  NAND2_X1 U488 ( .A1(n418), .A2(n417), .ZN(n420) );
  XNOR2_X1 U489 ( .A(KEYINPUT117), .B(KEYINPUT48), .ZN(n419) );
  XOR2_X1 U490 ( .A(n425), .B(n424), .Z(n429) );
  XNOR2_X1 U491 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U492 ( .A(n430), .B(KEYINPUT54), .ZN(n449) );
  XOR2_X1 U493 ( .A(n432), .B(n431), .Z(n434) );
  NAND2_X1 U494 ( .A1(G225GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U495 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U496 ( .A(n436), .B(n435), .ZN(n448) );
  XOR2_X1 U497 ( .A(KEYINPUT1), .B(KEYINPUT94), .Z(n438) );
  XNOR2_X1 U498 ( .A(G162GAT), .B(KEYINPUT4), .ZN(n437) );
  XNOR2_X1 U499 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U500 ( .A(KEYINPUT6), .B(KEYINPUT5), .Z(n440) );
  XNOR2_X1 U501 ( .A(KEYINPUT93), .B(KEYINPUT95), .ZN(n439) );
  XNOR2_X1 U502 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U503 ( .A(n442), .B(n441), .Z(n446) );
  XNOR2_X1 U504 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U505 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U506 ( .A(n448), .B(n447), .ZN(n467) );
  XNOR2_X1 U507 ( .A(KEYINPUT96), .B(n467), .ZN(n515) );
  NAND2_X1 U508 ( .A1(n449), .A2(n515), .ZN(n567) );
  XNOR2_X1 U509 ( .A(n450), .B(KEYINPUT55), .ZN(n451) );
  NAND2_X1 U510 ( .A1(n563), .A2(n532), .ZN(n455) );
  XOR2_X1 U511 ( .A(KEYINPUT124), .B(KEYINPUT56), .Z(n453) );
  XNOR2_X1 U512 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n452) );
  XNOR2_X1 U513 ( .A(n517), .B(KEYINPUT27), .ZN(n463) );
  NOR2_X1 U514 ( .A1(n463), .A2(n515), .ZN(n456) );
  XNOR2_X1 U515 ( .A(n456), .B(KEYINPUT97), .ZN(n544) );
  XOR2_X1 U516 ( .A(KEYINPUT28), .B(KEYINPUT64), .Z(n457) );
  XOR2_X1 U517 ( .A(n457), .B(n461), .Z(n490) );
  XNOR2_X1 U518 ( .A(n529), .B(KEYINPUT98), .ZN(n458) );
  NAND2_X1 U519 ( .A1(n527), .A2(n458), .ZN(n469) );
  NOR2_X1 U520 ( .A1(n527), .A2(n517), .ZN(n459) );
  NOR2_X1 U521 ( .A1(n461), .A2(n459), .ZN(n460) );
  XNOR2_X1 U522 ( .A(n460), .B(KEYINPUT25), .ZN(n465) );
  NAND2_X1 U523 ( .A1(n461), .A2(n527), .ZN(n462) );
  XOR2_X1 U524 ( .A(n462), .B(KEYINPUT26), .Z(n546) );
  INV_X1 U525 ( .A(n546), .ZN(n568) );
  OR2_X1 U526 ( .A1(n463), .A2(n568), .ZN(n464) );
  NAND2_X1 U527 ( .A1(n465), .A2(n464), .ZN(n466) );
  NAND2_X1 U528 ( .A1(n467), .A2(n466), .ZN(n468) );
  NAND2_X1 U529 ( .A1(n469), .A2(n468), .ZN(n479) );
  NAND2_X1 U530 ( .A1(n582), .A2(n479), .ZN(n470) );
  NOR2_X1 U531 ( .A1(n578), .A2(n470), .ZN(n473) );
  OR2_X1 U532 ( .A1(n548), .A2(n573), .ZN(n481) );
  NOR2_X1 U533 ( .A1(n514), .A2(n481), .ZN(n474) );
  XOR2_X1 U534 ( .A(KEYINPUT38), .B(n474), .Z(n499) );
  NOR2_X1 U535 ( .A1(n527), .A2(n499), .ZN(n477) );
  NOR2_X1 U536 ( .A1(n564), .A2(n555), .ZN(n478) );
  XNOR2_X1 U537 ( .A(n478), .B(KEYINPUT16), .ZN(n480) );
  NAND2_X1 U538 ( .A1(n480), .A2(n479), .ZN(n501) );
  OR2_X1 U539 ( .A1(n481), .A2(n501), .ZN(n491) );
  NOR2_X1 U540 ( .A1(n515), .A2(n491), .ZN(n483) );
  XNOR2_X1 U541 ( .A(KEYINPUT34), .B(KEYINPUT99), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U543 ( .A(G1GAT), .B(n484), .ZN(G1324GAT) );
  NOR2_X1 U544 ( .A1(n517), .A2(n491), .ZN(n485) );
  XOR2_X1 U545 ( .A(KEYINPUT100), .B(n485), .Z(n486) );
  XNOR2_X1 U546 ( .A(G8GAT), .B(n486), .ZN(G1325GAT) );
  NOR2_X1 U547 ( .A1(n527), .A2(n491), .ZN(n488) );
  XNOR2_X1 U548 ( .A(KEYINPUT101), .B(KEYINPUT35), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U550 ( .A(G15GAT), .B(n489), .Z(G1326GAT) );
  INV_X1 U551 ( .A(n490), .ZN(n523) );
  NOR2_X1 U552 ( .A1(n523), .A2(n491), .ZN(n493) );
  XNOR2_X1 U553 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U555 ( .A(G22GAT), .B(n494), .ZN(G1327GAT) );
  NOR2_X1 U556 ( .A1(n499), .A2(n515), .ZN(n496) );
  XNOR2_X1 U557 ( .A(KEYINPUT106), .B(KEYINPUT39), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U559 ( .A(G29GAT), .B(n497), .ZN(G1328GAT) );
  NOR2_X1 U560 ( .A1(n517), .A2(n499), .ZN(n498) );
  XOR2_X1 U561 ( .A(G36GAT), .B(n498), .Z(G1329GAT) );
  NOR2_X1 U562 ( .A1(n523), .A2(n499), .ZN(n500) );
  XOR2_X1 U563 ( .A(G50GAT), .B(n500), .Z(G1331GAT) );
  NAND2_X1 U564 ( .A1(n548), .A2(n532), .ZN(n513) );
  NOR2_X1 U565 ( .A1(n513), .A2(n501), .ZN(n502) );
  XNOR2_X1 U566 ( .A(KEYINPUT107), .B(n502), .ZN(n510) );
  NOR2_X1 U567 ( .A1(n515), .A2(n510), .ZN(n504) );
  XNOR2_X1 U568 ( .A(KEYINPUT42), .B(KEYINPUT108), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U570 ( .A(G57GAT), .B(n505), .Z(G1332GAT) );
  NOR2_X1 U571 ( .A1(n517), .A2(n510), .ZN(n507) );
  XNOR2_X1 U572 ( .A(G64GAT), .B(KEYINPUT109), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n507), .B(n506), .ZN(G1333GAT) );
  NOR2_X1 U574 ( .A1(n527), .A2(n510), .ZN(n508) );
  XOR2_X1 U575 ( .A(KEYINPUT110), .B(n508), .Z(n509) );
  XNOR2_X1 U576 ( .A(G71GAT), .B(n509), .ZN(G1334GAT) );
  NOR2_X1 U577 ( .A1(n523), .A2(n510), .ZN(n512) );
  XNOR2_X1 U578 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n511) );
  XNOR2_X1 U579 ( .A(n512), .B(n511), .ZN(G1335GAT) );
  OR2_X1 U580 ( .A1(n514), .A2(n513), .ZN(n522) );
  NOR2_X1 U581 ( .A1(n515), .A2(n522), .ZN(n516) );
  XOR2_X1 U582 ( .A(G85GAT), .B(n516), .Z(G1336GAT) );
  NOR2_X1 U583 ( .A1(n517), .A2(n522), .ZN(n519) );
  XNOR2_X1 U584 ( .A(G92GAT), .B(KEYINPUT111), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(G1337GAT) );
  NOR2_X1 U586 ( .A1(n527), .A2(n522), .ZN(n520) );
  XOR2_X1 U587 ( .A(KEYINPUT112), .B(n520), .Z(n521) );
  XNOR2_X1 U588 ( .A(G99GAT), .B(n521), .ZN(G1338GAT) );
  NOR2_X1 U589 ( .A1(n523), .A2(n522), .ZN(n525) );
  XNOR2_X1 U590 ( .A(KEYINPUT44), .B(KEYINPUT113), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  NOR2_X1 U593 ( .A1(n545), .A2(n527), .ZN(n528) );
  NAND2_X1 U594 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U595 ( .A(KEYINPUT118), .B(n530), .Z(n540) );
  INV_X1 U596 ( .A(n540), .ZN(n536) );
  NOR2_X1 U597 ( .A1(n536), .A2(n548), .ZN(n531) );
  XOR2_X1 U598 ( .A(G113GAT), .B(n531), .Z(G1340GAT) );
  XNOR2_X1 U599 ( .A(KEYINPUT119), .B(KEYINPUT49), .ZN(n534) );
  INV_X1 U600 ( .A(n532), .ZN(n552) );
  NOR2_X1 U601 ( .A1(n552), .A2(n536), .ZN(n533) );
  XNOR2_X1 U602 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U603 ( .A(G120GAT), .B(n535), .Z(G1341GAT) );
  NOR2_X1 U604 ( .A1(n536), .A2(n555), .ZN(n538) );
  XNOR2_X1 U605 ( .A(KEYINPUT50), .B(KEYINPUT120), .ZN(n537) );
  XNOR2_X1 U606 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U607 ( .A(G127GAT), .B(n539), .Z(G1342GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT121), .B(KEYINPUT51), .Z(n542) );
  NAND2_X1 U609 ( .A1(n540), .A2(n564), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U611 ( .A(G134GAT), .B(n543), .Z(G1343GAT) );
  NOR2_X1 U612 ( .A1(n545), .A2(n544), .ZN(n547) );
  NAND2_X1 U613 ( .A1(n547), .A2(n546), .ZN(n558) );
  NOR2_X1 U614 ( .A1(n548), .A2(n558), .ZN(n549) );
  XOR2_X1 U615 ( .A(G141GAT), .B(n549), .Z(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT52), .B(KEYINPUT122), .Z(n551) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(n554) );
  NOR2_X1 U619 ( .A1(n552), .A2(n558), .ZN(n553) );
  XOR2_X1 U620 ( .A(n554), .B(n553), .Z(G1345GAT) );
  NOR2_X1 U621 ( .A1(n555), .A2(n558), .ZN(n557) );
  XNOR2_X1 U622 ( .A(G155GAT), .B(KEYINPUT123), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1346GAT) );
  NOR2_X1 U624 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U625 ( .A(G162GAT), .B(n560), .Z(G1347GAT) );
  NAND2_X1 U626 ( .A1(n563), .A2(n569), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U628 ( .A1(n563), .A2(n578), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(KEYINPUT58), .ZN(n566) );
  XNOR2_X1 U632 ( .A(G190GAT), .B(n566), .ZN(G1351GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n571) );
  NOR2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n581) );
  NAND2_X1 U635 ( .A1(n581), .A2(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n575) );
  NAND2_X1 U639 ( .A1(n581), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n577) );
  XOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT125), .Z(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  XOR2_X1 U643 ( .A(G211GAT), .B(KEYINPUT127), .Z(n580) );
  NAND2_X1 U644 ( .A1(n581), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1354GAT) );
  NAND2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(n583), .B(KEYINPUT62), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

