//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n786,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n866, new_n867, new_n869, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n992, new_n993, new_n994;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT13), .Z(new_n203));
  AND2_X1   g002(.A1(G43gat), .A2(G50gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(G43gat), .A2(G50gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT91), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G43gat), .ZN(new_n207));
  INV_X1    g006(.A(G50gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT91), .ZN(new_n210));
  NAND2_X1  g009(.A1(G43gat), .A2(G50gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n206), .A2(new_n212), .A3(KEYINPUT15), .ZN(new_n213));
  INV_X1    g012(.A(G29gat), .ZN(new_n214));
  INV_X1    g013(.A(G36gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n215), .A3(KEYINPUT14), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT14), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(G29gat), .B2(G36gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT92), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n216), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n220), .A2(KEYINPUT92), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n213), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G15gat), .B(G22gat), .ZN(new_n226));
  INV_X1    g025(.A(G1gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT16), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  OAI221_X1 g028(.A(new_n229), .B1(KEYINPUT97), .B2(G8gat), .C1(G1gat), .C2(new_n226), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n229), .B1(G1gat), .B2(new_n226), .ZN(new_n231));
  INV_X1    g030(.A(G8gat), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT97), .B1(new_n226), .B2(G1gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT93), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n204), .A2(new_n205), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT15), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NOR4_X1   g037(.A1(new_n204), .A2(new_n205), .A3(KEYINPUT93), .A4(KEYINPUT15), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n213), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AND3_X1   g039(.A1(new_n217), .A2(new_n219), .A3(KEYINPUT94), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT94), .B1(new_n217), .B2(new_n219), .ZN(new_n242));
  OAI22_X1  g041(.A1(new_n241), .A2(new_n242), .B1(new_n214), .B2(new_n215), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT95), .B1(new_n240), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT94), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n220), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n217), .A2(new_n219), .A3(KEYINPUT94), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n216), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT95), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n209), .A2(new_n211), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT93), .B1(new_n250), .B2(KEYINPUT15), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n236), .A2(new_n235), .A3(new_n237), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n248), .A2(new_n249), .A3(new_n253), .A4(new_n213), .ZN(new_n254));
  AOI221_X4 g053(.A(new_n225), .B1(new_n230), .B2(new_n234), .C1(new_n244), .C2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n234), .A2(new_n230), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n244), .A2(new_n254), .ZN(new_n257));
  INV_X1    g056(.A(new_n225), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n203), .B1(new_n255), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT99), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT99), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n262), .B(new_n203), .C1(new_n255), .C2(new_n259), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n257), .A2(new_n258), .ZN(new_n264));
  INV_X1    g063(.A(new_n256), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n225), .B1(new_n244), .B2(new_n254), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT96), .B(KEYINPUT17), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n256), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT17), .ZN(new_n270));
  AOI211_X1 g069(.A(new_n270), .B(new_n225), .C1(new_n244), .C2(new_n254), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n266), .B(new_n202), .C1(new_n269), .C2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT18), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n261), .A2(new_n263), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n273), .B1(G229gat), .B2(G233gat), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n266), .B(new_n275), .C1(new_n269), .C2(new_n271), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT98), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n267), .A2(KEYINPUT17), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n278), .B(new_n256), .C1(new_n267), .C2(new_n268), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT98), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n279), .A2(new_n280), .A3(new_n266), .A4(new_n275), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G113gat), .B(G141gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(G197gat), .ZN(new_n284));
  XOR2_X1   g083(.A(KEYINPUT11), .B(G169gat), .Z(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT90), .B(KEYINPUT12), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  AND3_X1   g087(.A1(new_n274), .A2(new_n282), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n288), .B1(new_n274), .B2(new_n282), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G78gat), .B(G106gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n292), .B(G22gat), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  XOR2_X1   g093(.A(G141gat), .B(G148gat), .Z(new_n295));
  INV_X1    g094(.A(G155gat), .ZN(new_n296));
  INV_X1    g095(.A(G162gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(KEYINPUT2), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n295), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G141gat), .B(G148gat), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n299), .B(new_n298), .C1(new_n303), .C2(KEYINPUT2), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G197gat), .B(G204gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT22), .ZN(new_n307));
  INV_X1    g106(.A(G211gat), .ZN(new_n308));
  INV_X1    g107(.A(G218gat), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G211gat), .B(G218gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(KEYINPUT29), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n305), .B1(new_n314), .B2(KEYINPUT3), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(KEYINPUT74), .ZN(new_n316));
  INV_X1    g115(.A(new_n312), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n311), .B(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT74), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  XOR2_X1   g119(.A(KEYINPUT80), .B(KEYINPUT3), .Z(new_n321));
  NAND3_X1  g120(.A1(new_n302), .A2(new_n304), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n316), .A2(new_n320), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n315), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n326), .A2(G228gat), .A3(G233gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(KEYINPUT88), .ZN(new_n328));
  NAND2_X1  g127(.A1(G228gat), .A2(G233gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT88), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n316), .A2(new_n320), .A3(new_n330), .A4(new_n324), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n321), .B1(new_n313), .B2(KEYINPUT29), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(new_n305), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n328), .A2(new_n329), .A3(new_n331), .A4(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT31), .B(G50gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  AND3_X1   g135(.A1(new_n327), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n336), .B1(new_n327), .B2(new_n334), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n294), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n327), .A2(new_n334), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(new_n335), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n327), .A2(new_n334), .A3(new_n336), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n341), .A2(new_n293), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n316), .A2(new_n320), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G226gat), .A2(G233gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n347), .B(KEYINPUT75), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n350));
  AND3_X1   g149(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n352));
  OAI22_X1  g151(.A1(new_n351), .A2(KEYINPUT65), .B1(new_n352), .B2(KEYINPUT66), .ZN(new_n353));
  NAND3_X1  g152(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT65), .ZN(new_n355));
  OAI22_X1  g154(.A1(new_n354), .A2(new_n355), .B1(G183gat), .B2(G190gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(G183gat), .A2(G190gat), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT24), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n357), .A2(KEYINPUT66), .A3(new_n358), .ZN(new_n359));
  NOR3_X1   g158(.A1(new_n353), .A2(new_n356), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(G169gat), .ZN(new_n361));
  INV_X1    g160(.A(G176gat), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT23), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(G169gat), .A2(G176gat), .ZN(new_n364));
  MUX2_X1   g163(.A(new_n363), .B(KEYINPUT23), .S(new_n364), .Z(new_n365));
  OAI21_X1  g164(.A(new_n350), .B1(new_n360), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n357), .A2(KEYINPUT68), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT68), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n368), .A2(G183gat), .A3(G190gat), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n367), .A2(new_n369), .A3(new_n358), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT69), .ZN(new_n371));
  INV_X1    g170(.A(G183gat), .ZN(new_n372));
  INV_X1    g171(.A(G190gat), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT69), .B1(G183gat), .B2(G190gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n370), .A2(new_n354), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT25), .ZN(new_n378));
  INV_X1    g177(.A(new_n364), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n378), .B1(new_n363), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT67), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(KEYINPUT23), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT70), .B1(new_n377), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n376), .A3(new_n354), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT70), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n387), .A2(new_n388), .A3(new_n384), .A4(new_n380), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n366), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n361), .A2(new_n362), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n391), .B1(KEYINPUT26), .B2(new_n379), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT26), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n382), .A2(new_n393), .A3(new_n383), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n392), .A2(new_n394), .B1(G183gat), .B2(G190gat), .ZN(new_n395));
  OAI211_X1 g194(.A(KEYINPUT71), .B(new_n373), .C1(new_n372), .C2(KEYINPUT27), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT28), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT72), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n372), .A2(KEYINPUT27), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n373), .B1(new_n372), .B2(KEYINPUT27), .ZN(new_n402));
  OR2_X1    g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n396), .A2(KEYINPUT72), .A3(new_n397), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n400), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n403), .B1(new_n400), .B2(new_n404), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n395), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n349), .B1(new_n390), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT76), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n390), .A2(new_n410), .A3(new_n407), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n410), .B1(new_n390), .B2(new_n407), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n411), .A2(new_n412), .A3(KEYINPUT29), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n346), .B(new_n409), .C1(new_n413), .C2(new_n348), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n348), .B1(new_n411), .B2(new_n412), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n390), .A2(new_n407), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n348), .A2(KEYINPUT29), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n415), .A2(new_n345), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT77), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT77), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n414), .A2(new_n422), .A3(new_n419), .ZN(new_n423));
  XNOR2_X1  g222(.A(G8gat), .B(G36gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n424), .B(KEYINPUT78), .ZN(new_n425));
  XNOR2_X1  g224(.A(G64gat), .B(G92gat), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n425), .B(new_n426), .Z(new_n427));
  NAND3_X1  g226(.A1(new_n421), .A2(new_n423), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n427), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n416), .A2(KEYINPUT76), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n390), .A2(new_n410), .A3(new_n407), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(new_n323), .A3(new_n431), .ZN(new_n432));
  AOI211_X1 g231(.A(new_n345), .B(new_n408), .C1(new_n432), .C2(new_n349), .ZN(new_n433));
  INV_X1    g232(.A(new_n419), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n429), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT79), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT30), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n427), .B1(new_n414), .B2(new_n419), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT79), .B1(new_n439), .B2(KEYINPUT30), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(KEYINPUT30), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n428), .A2(new_n438), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(G57gat), .B(G85gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n443), .B(KEYINPUT84), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n444), .B(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(G1gat), .B(G29gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n446), .B(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT5), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n305), .A2(KEYINPUT3), .ZN(new_n450));
  AND2_X1   g249(.A1(KEYINPUT73), .A2(G127gat), .ZN(new_n451));
  NOR2_X1   g250(.A1(KEYINPUT73), .A2(G127gat), .ZN(new_n452));
  OAI21_X1  g251(.A(G134gat), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  OR2_X1    g252(.A1(G127gat), .A2(G134gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(G113gat), .B(G120gat), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n453), .B(new_n454), .C1(KEYINPUT1), .C2(new_n455), .ZN(new_n456));
  XOR2_X1   g255(.A(G113gat), .B(G120gat), .Z(new_n457));
  INV_X1    g256(.A(KEYINPUT1), .ZN(new_n458));
  XNOR2_X1  g257(.A(G127gat), .B(G134gat), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n450), .A2(new_n461), .A3(new_n322), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT81), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n450), .A2(KEYINPUT81), .A3(new_n461), .A4(new_n322), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(G225gat), .A2(G233gat), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n456), .A2(new_n302), .A3(new_n460), .A4(new_n304), .ZN(new_n469));
  OR2_X1    g268(.A1(new_n469), .A2(KEYINPUT4), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(KEYINPUT4), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n449), .B1(new_n466), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n461), .A2(new_n305), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(new_n469), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n468), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n476), .B(KEYINPUT82), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n448), .B1(new_n473), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT85), .B1(new_n469), .B2(KEYINPUT4), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n469), .A2(KEYINPUT86), .A3(KEYINPUT4), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT86), .B1(new_n469), .B2(KEYINPUT4), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n479), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT86), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n471), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n485), .A2(new_n470), .A3(KEYINPUT85), .A4(new_n480), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n468), .A2(KEYINPUT5), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n483), .A2(new_n466), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n478), .A2(KEYINPUT87), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT6), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n448), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n473), .A2(new_n477), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n492), .B1(new_n493), .B2(new_n488), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT87), .B1(new_n478), .B2(new_n488), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n490), .B1(new_n497), .B2(new_n494), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n344), .B1(new_n442), .B2(new_n499), .ZN(new_n500));
  XOR2_X1   g299(.A(G15gat), .B(G43gat), .Z(new_n501));
  XNOR2_X1  g300(.A(G71gat), .B(G99gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n390), .A2(new_n461), .A3(new_n407), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n461), .B1(new_n390), .B2(new_n407), .ZN(new_n505));
  NAND2_X1  g304(.A1(G227gat), .A2(G233gat), .ZN(new_n506));
  NOR3_X1   g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n503), .B1(new_n507), .B2(KEYINPUT33), .ZN(new_n508));
  INV_X1    g307(.A(new_n461), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n416), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n390), .A2(new_n461), .A3(new_n407), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(new_n506), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT34), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT34), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n515), .B(new_n506), .C1(new_n504), .C2(new_n505), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n508), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n503), .ZN(new_n518));
  INV_X1    g317(.A(new_n506), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n510), .A2(new_n519), .A3(new_n511), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT33), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n515), .B1(new_n512), .B2(new_n506), .ZN(new_n523));
  INV_X1    g322(.A(new_n516), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n520), .A2(KEYINPUT32), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n517), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n527), .B1(new_n517), .B2(new_n525), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT36), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n339), .A2(new_n343), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT38), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT37), .ZN(new_n534));
  AOI211_X1 g333(.A(new_n533), .B(new_n429), .C1(new_n420), .C2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n421), .A2(new_n423), .A3(KEYINPUT37), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n420), .A2(new_n534), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n415), .A2(new_n418), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n346), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n408), .B1(new_n432), .B2(new_n349), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n539), .B(KEYINPUT37), .C1(new_n540), .C2(new_n346), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n537), .A2(new_n427), .A3(new_n541), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n535), .A2(new_n536), .B1(new_n542), .B2(new_n533), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n499), .A2(new_n435), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n532), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AND4_X1   g344(.A1(new_n428), .A2(new_n438), .A3(new_n440), .A4(new_n441), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT39), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n483), .A2(new_n466), .A3(new_n486), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT89), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n548), .A2(new_n549), .A3(new_n468), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n549), .B1(new_n548), .B2(new_n468), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n547), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n552), .ZN(new_n554));
  INV_X1    g353(.A(new_n475), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n547), .B1(new_n555), .B2(new_n467), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n554), .A2(new_n550), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n553), .A2(new_n557), .A3(new_n492), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT40), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n553), .A2(new_n557), .A3(KEYINPUT40), .A4(new_n492), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(new_n495), .A3(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n546), .A2(new_n562), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n500), .B(new_n531), .C1(new_n545), .C2(new_n563), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n428), .A2(new_n441), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n438), .A2(new_n440), .ZN(new_n566));
  NOR3_X1   g365(.A1(new_n528), .A2(new_n529), .A3(new_n344), .ZN(new_n567));
  INV_X1    g366(.A(new_n499), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n565), .A2(new_n566), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT35), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n442), .A2(new_n499), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT35), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n571), .A2(new_n572), .A3(new_n567), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n291), .B1(new_n564), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT103), .ZN(new_n576));
  XNOR2_X1  g375(.A(G134gat), .B(G162gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT41), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n577), .B(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(G92gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT101), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT101), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(G92gat), .ZN(new_n585));
  INV_X1    g384(.A(G85gat), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n583), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G85gat), .A2(G92gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT7), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT7), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n590), .A2(G85gat), .A3(G92gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G99gat), .A2(G106gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(KEYINPUT8), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n587), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  OR2_X1    g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT102), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n596), .A2(new_n597), .A3(new_n593), .ZN(new_n598));
  AND2_X1   g397(.A1(G99gat), .A2(G106gat), .ZN(new_n599));
  NOR2_X1   g398(.A1(G99gat), .A2(G106gat), .ZN(new_n600));
  OAI21_X1  g399(.A(KEYINPUT102), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n595), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n595), .A2(new_n602), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI22_X1  g404(.A1(new_n267), .A2(new_n605), .B1(new_n579), .B2(new_n578), .ZN(new_n606));
  INV_X1    g405(.A(new_n605), .ZN(new_n607));
  INV_X1    g406(.A(new_n268), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n607), .B1(new_n264), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n606), .B1(new_n609), .B2(new_n278), .ZN(new_n610));
  XNOR2_X1  g409(.A(G190gat), .B(G218gat), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT100), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n278), .B(new_n605), .C1(new_n267), .C2(new_n268), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n578), .A2(new_n579), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n614), .B1(new_n264), .B2(new_n607), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n611), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n581), .B1(new_n612), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n605), .B1(new_n267), .B2(new_n268), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n615), .B(new_n611), .C1(new_n271), .C2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT100), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n581), .ZN(new_n623));
  NOR3_X1   g422(.A1(new_n622), .A2(new_n616), .A3(new_n623), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n618), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(G57gat), .B(G64gat), .Z(new_n626));
  OR2_X1    g425(.A1(G71gat), .A2(G78gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(G71gat), .A2(G78gat), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT9), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n626), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G57gat), .B(G64gat), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n628), .B(new_n627), .C1(new_n633), .C2(new_n630), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT21), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(G231gat), .A2(G233gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(G127gat), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n256), .B1(new_n636), .B2(new_n635), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(new_n296), .ZN(new_n644));
  XNOR2_X1  g443(.A(G183gat), .B(G211gat), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n644), .B(new_n645), .Z(new_n646));
  XNOR2_X1  g445(.A(new_n642), .B(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n576), .B1(new_n625), .B2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n646), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n642), .B(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n618), .A2(new_n624), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n650), .A2(KEYINPUT103), .A3(new_n651), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n632), .A2(new_n634), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n653), .B1(new_n603), .B2(new_n604), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT10), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT101), .B(G92gat), .ZN(new_n656));
  AOI22_X1  g455(.A1(new_n656), .A2(new_n586), .B1(KEYINPUT8), .B2(new_n593), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n657), .A2(new_n601), .A3(new_n598), .A4(new_n592), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n595), .A2(new_n602), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(new_n635), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n654), .A2(new_n655), .A3(new_n660), .ZN(new_n661));
  OAI211_X1 g460(.A(new_n653), .B(KEYINPUT10), .C1(new_n603), .C2(new_n604), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(G230gat), .A2(G233gat), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n664), .B(KEYINPUT104), .Z(new_n665));
  OAI21_X1  g464(.A(KEYINPUT105), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n665), .B1(new_n661), .B2(new_n662), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT105), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n665), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n670), .B1(new_n654), .B2(new_n660), .ZN(new_n671));
  XNOR2_X1  g470(.A(G120gat), .B(G148gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(G176gat), .B(G204gat), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n672), .B(new_n673), .Z(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n666), .A2(new_n669), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n675), .B1(new_n667), .B2(new_n671), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(KEYINPUT106), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT106), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n677), .A2(new_n681), .A3(new_n678), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  AND3_X1   g483(.A1(new_n648), .A2(new_n652), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n575), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n686), .A2(new_n568), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(new_n227), .ZN(G1324gat));
  AND2_X1   g487(.A1(new_n575), .A2(new_n442), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT16), .B(G8gat), .Z(new_n690));
  AND3_X1   g489(.A1(new_n689), .A2(new_n685), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n232), .B1(new_n689), .B2(new_n685), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT42), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n693), .B1(KEYINPUT42), .B2(new_n691), .ZN(G1325gat));
  OAI21_X1  g493(.A(G15gat), .B1(new_n686), .B2(new_n531), .ZN(new_n695));
  INV_X1    g494(.A(new_n530), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n696), .A2(G15gat), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n695), .B1(new_n686), .B2(new_n697), .ZN(G1326gat));
  NOR2_X1   g497(.A1(new_n686), .A2(new_n532), .ZN(new_n699));
  XOR2_X1   g498(.A(KEYINPUT43), .B(G22gat), .Z(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1327gat));
  AOI21_X1  g500(.A(new_n572), .B1(new_n571), .B2(new_n567), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n517), .A2(new_n525), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(new_n526), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n517), .A2(new_n525), .A3(new_n527), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n704), .A2(new_n532), .A3(new_n705), .ZN(new_n706));
  NOR4_X1   g505(.A1(new_n442), .A2(new_n706), .A3(new_n499), .A4(KEYINPUT35), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT109), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n702), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(KEYINPUT109), .B1(new_n570), .B2(new_n573), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n564), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n711), .A2(new_n712), .A3(new_n625), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n564), .A2(new_n574), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n712), .B1(new_n714), .B2(new_n625), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n650), .A2(new_n683), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n719), .A2(new_n291), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT108), .Z(new_n721));
  NAND2_X1  g520(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(G29gat), .B1(new_n722), .B2(new_n568), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n714), .A2(new_n625), .A3(new_n720), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT107), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n568), .A2(G29gat), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n725), .B1(new_n724), .B2(new_n726), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT45), .ZN(new_n729));
  OR3_X1    g528(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n729), .B1(new_n727), .B2(new_n728), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n723), .A2(new_n730), .A3(new_n731), .ZN(G1328gat));
  OAI21_X1  g531(.A(G36gat), .B1(new_n722), .B2(new_n546), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n719), .A2(G36gat), .A3(new_n651), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n689), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT46), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n735), .B1(KEYINPUT110), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(KEYINPUT110), .B(KEYINPUT46), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n733), .B(new_n737), .C1(new_n735), .C2(new_n738), .ZN(G1329gat));
  INV_X1    g538(.A(new_n531), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n625), .A2(new_n712), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n708), .B1(new_n702), .B2(new_n707), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n570), .A2(new_n573), .A3(KEYINPUT109), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n741), .B1(new_n744), .B2(new_n564), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n740), .B(new_n721), .C1(new_n745), .C2(new_n715), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(G43gat), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n724), .A2(new_n207), .A3(new_n530), .ZN(new_n748));
  XNOR2_X1  g547(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n749), .B1(new_n747), .B2(new_n748), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n750), .A2(new_n751), .ZN(G1330gat));
  OAI211_X1 g551(.A(new_n344), .B(new_n721), .C1(new_n745), .C2(new_n715), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G50gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(KEYINPUT112), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n724), .A2(new_n208), .A3(new_n344), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT48), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n755), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n754), .B(new_n756), .C1(KEYINPUT112), .C2(KEYINPUT48), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(G1331gat));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n762));
  OR2_X1    g561(.A1(new_n545), .A2(new_n563), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n531), .A2(new_n500), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n742), .A2(new_n743), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n648), .A2(new_n652), .A3(new_n291), .A4(new_n683), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n762), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n766), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n711), .A2(KEYINPUT113), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n499), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g572(.A(KEYINPUT49), .B(G64gat), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n771), .A2(new_n442), .A3(new_n774), .ZN(new_n775));
  OAI22_X1  g574(.A1(new_n770), .A2(new_n546), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(G1333gat));
  OAI21_X1  g576(.A(G71gat), .B1(new_n770), .B2(new_n531), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n696), .A2(G71gat), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n767), .A2(new_n769), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n778), .A2(KEYINPUT50), .A3(new_n780), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(G1334gat));
  NAND2_X1  g584(.A1(new_n771), .A2(new_n344), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(G78gat), .ZN(G1335gat));
  INV_X1    g586(.A(new_n291), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n650), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n683), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n717), .A2(new_n499), .A3(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n790), .B1(new_n713), .B2(new_n716), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n795), .A2(KEYINPUT114), .A3(new_n499), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n794), .A2(G85gat), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n789), .A2(new_n625), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n765), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n799), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n711), .A2(KEYINPUT51), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n803), .A2(new_n586), .A3(new_n499), .A4(new_n683), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n797), .A2(new_n804), .ZN(G1336gat));
  OAI211_X1 g604(.A(new_n442), .B(new_n791), .C1(new_n745), .C2(new_n715), .ZN(new_n806));
  INV_X1    g605(.A(new_n656), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n803), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n546), .A2(G92gat), .A3(new_n684), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n808), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(KEYINPUT52), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n808), .B(new_n814), .C1(new_n809), .C2(new_n811), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n815), .ZN(G1337gat));
  NAND2_X1  g615(.A1(new_n795), .A2(new_n740), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(G99gat), .ZN(new_n818));
  OR3_X1    g617(.A1(new_n696), .A2(G99gat), .A3(new_n684), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n818), .B1(new_n809), .B2(new_n819), .ZN(G1338gat));
  OAI211_X1 g619(.A(new_n344), .B(new_n791), .C1(new_n745), .C2(new_n715), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(G106gat), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n684), .A2(new_n532), .A3(G106gat), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n803), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(KEYINPUT115), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(KEYINPUT115), .ZN(new_n828));
  AND4_X1   g627(.A1(new_n822), .A2(new_n824), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n826), .B1(new_n803), .B2(new_n823), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n828), .B1(new_n830), .B2(new_n822), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n829), .A2(new_n831), .ZN(G1339gat));
  NAND4_X1  g631(.A1(new_n648), .A2(new_n652), .A3(new_n291), .A4(new_n684), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n274), .A2(new_n282), .A3(new_n288), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n202), .B1(new_n279), .B2(new_n266), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n255), .A2(new_n259), .A3(new_n203), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n286), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n834), .B(new_n837), .C1(new_n618), .C2(new_n624), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n661), .A2(new_n662), .A3(new_n665), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT116), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n661), .A2(KEYINPUT116), .A3(new_n662), .A4(new_n665), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n843), .A2(new_n666), .A3(KEYINPUT54), .A4(new_n669), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n674), .B1(new_n667), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT55), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n844), .A2(KEYINPUT55), .A3(new_n846), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n849), .A2(new_n677), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n838), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n683), .A2(new_n834), .A3(new_n837), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n853), .B1(new_n291), .B2(new_n851), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n852), .B1(new_n854), .B2(new_n651), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n833), .B1(new_n855), .B2(new_n650), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n856), .A2(new_n532), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n857), .A2(new_n499), .A3(new_n530), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n546), .ZN(new_n859));
  OAI21_X1  g658(.A(G113gat), .B1(new_n859), .B2(new_n291), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n291), .A2(G113gat), .ZN(new_n861));
  XOR2_X1   g660(.A(new_n861), .B(KEYINPUT117), .Z(new_n862));
  OAI21_X1  g661(.A(new_n860), .B1(new_n859), .B2(new_n862), .ZN(G1340gat));
  NOR2_X1   g662(.A1(new_n859), .A2(new_n684), .ZN(new_n864));
  XOR2_X1   g663(.A(new_n864), .B(G120gat), .Z(G1341gat));
  NOR2_X1   g664(.A1(new_n859), .A2(new_n647), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n451), .A2(new_n452), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n866), .B(new_n867), .ZN(G1342gat));
  NOR3_X1   g667(.A1(new_n442), .A2(G134gat), .A3(new_n651), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n858), .A2(new_n869), .ZN(new_n870));
  XOR2_X1   g669(.A(new_n870), .B(KEYINPUT56), .Z(new_n871));
  OAI21_X1  g670(.A(G134gat), .B1(new_n859), .B2(new_n651), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(G1343gat));
  NOR2_X1   g672(.A1(new_n442), .A2(new_n568), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n740), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT57), .B1(new_n856), .B2(new_n344), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n532), .A2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n847), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n844), .A2(KEYINPUT118), .A3(new_n846), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n882), .A2(new_n848), .A3(new_n883), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n850), .A2(new_n677), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n884), .B(new_n885), .C1(new_n290), .C2(new_n289), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n625), .B1(new_n886), .B2(new_n853), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n647), .B1(new_n887), .B2(new_n852), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n880), .B1(new_n888), .B2(new_n833), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n876), .B1(new_n877), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(G141gat), .B1(new_n890), .B2(new_n291), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n531), .A2(new_n344), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n875), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n531), .A2(KEYINPUT119), .A3(new_n344), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n894), .A2(new_n856), .A3(new_n895), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n291), .A2(G141gat), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n891), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n740), .A2(new_n684), .A3(new_n875), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n885), .B1(new_n289), .B2(new_n290), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n882), .A2(new_n848), .A3(new_n883), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n853), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n852), .B1(new_n904), .B2(new_n651), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n833), .B1(new_n905), .B2(new_n650), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT57), .B1(new_n906), .B2(new_n344), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n856), .A2(new_n879), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n901), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n900), .B1(new_n910), .B2(G148gat), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n683), .B(new_n876), .C1(new_n877), .C2(new_n889), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n900), .A2(G148gat), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT120), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT120), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n912), .A2(new_n916), .A3(new_n913), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n911), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n896), .A2(G148gat), .A3(new_n684), .ZN(new_n919));
  OAI21_X1  g718(.A(KEYINPUT121), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT121), .ZN(new_n921));
  INV_X1    g720(.A(new_n919), .ZN(new_n922));
  AND3_X1   g721(.A1(new_n912), .A2(new_n916), .A3(new_n913), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n916), .B1(new_n912), .B2(new_n913), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n921), .B(new_n922), .C1(new_n925), .C2(new_n911), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n920), .A2(new_n926), .ZN(G1345gat));
  OAI21_X1  g726(.A(G155gat), .B1(new_n890), .B2(new_n647), .ZN(new_n928));
  INV_X1    g727(.A(new_n896), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n929), .A2(new_n296), .A3(new_n650), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1346gat));
  OAI21_X1  g730(.A(G162gat), .B1(new_n890), .B2(new_n651), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n929), .A2(new_n297), .A3(new_n625), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1347gat));
  NOR3_X1   g733(.A1(new_n546), .A2(new_n696), .A3(new_n499), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n857), .A2(new_n935), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n936), .A2(new_n361), .A3(new_n291), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n856), .A2(new_n568), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n938), .A2(new_n442), .A3(new_n567), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(new_n788), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n937), .B1(new_n940), .B2(new_n361), .ZN(G1348gat));
  NAND3_X1  g740(.A1(new_n939), .A2(new_n362), .A3(new_n683), .ZN(new_n942));
  OAI21_X1  g741(.A(G176gat), .B1(new_n936), .B2(new_n684), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1349gat));
  NOR2_X1   g743(.A1(new_n372), .A2(KEYINPUT27), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n647), .A2(new_n401), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n857), .A2(new_n650), .A3(new_n935), .ZN(new_n947));
  AOI22_X1  g746(.A1(new_n939), .A2(new_n946), .B1(new_n947), .B2(G183gat), .ZN(new_n948));
  XOR2_X1   g747(.A(new_n948), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g748(.A1(new_n939), .A2(new_n373), .A3(new_n625), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n856), .A2(new_n532), .A3(new_n625), .A4(new_n935), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(G190gat), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(KEYINPUT61), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT122), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n952), .A2(new_n955), .A3(KEYINPUT61), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT123), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n958), .B1(new_n952), .B2(KEYINPUT61), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n951), .A2(KEYINPUT123), .A3(new_n960), .A4(G190gat), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n950), .B1(new_n957), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(KEYINPUT124), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT124), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n965), .B(new_n950), .C1(new_n957), .C2(new_n962), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n964), .A2(new_n966), .ZN(G1351gat));
  NOR2_X1   g766(.A1(new_n892), .A2(new_n546), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n938), .A2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  XNOR2_X1  g769(.A(KEYINPUT125), .B(G197gat), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n970), .A2(new_n788), .A3(new_n971), .ZN(new_n972));
  OR2_X1    g771(.A1(new_n907), .A2(new_n909), .ZN(new_n973));
  NOR3_X1   g772(.A1(new_n740), .A2(new_n499), .A3(new_n546), .ZN(new_n974));
  AND2_X1   g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT126), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n975), .A2(new_n976), .A3(new_n788), .ZN(new_n977));
  INV_X1    g776(.A(new_n971), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n976), .B1(new_n975), .B2(new_n788), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n972), .B1(new_n979), .B2(new_n980), .ZN(G1352gat));
  NAND2_X1  g780(.A1(new_n975), .A2(new_n683), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(G204gat), .ZN(new_n983));
  NOR3_X1   g782(.A1(new_n969), .A2(G204gat), .A3(new_n684), .ZN(new_n984));
  XNOR2_X1  g783(.A(new_n984), .B(KEYINPUT62), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n983), .A2(new_n985), .ZN(G1353gat));
  NAND3_X1  g785(.A1(new_n970), .A2(new_n308), .A3(new_n650), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n973), .A2(new_n650), .A3(new_n974), .ZN(new_n988));
  AND3_X1   g787(.A1(new_n988), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n989));
  AOI21_X1  g788(.A(KEYINPUT63), .B1(new_n988), .B2(G211gat), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n987), .B1(new_n989), .B2(new_n990), .ZN(G1354gat));
  NAND3_X1  g790(.A1(new_n970), .A2(new_n309), .A3(new_n625), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n975), .A2(new_n625), .ZN(new_n993));
  INV_X1    g792(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n992), .B1(new_n994), .B2(new_n309), .ZN(G1355gat));
endmodule


