//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 1 0 0 1 1 0 0 0 1 1 1 0 1 1 0 0 1 0 1 0 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 1 1 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  INV_X1    g0016(.A(new_n201), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  OR3_X1    g0019(.A1(new_n218), .A2(new_n211), .A3(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G87), .ZN(new_n224));
  INV_X1    g0024(.A(G250), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n227));
  INV_X1    g0027(.A(G58), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  INV_X1    g0029(.A(G257), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n227), .B1(new_n228), .B2(new_n229), .C1(new_n206), .C2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n213), .B1(new_n226), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n216), .B(new_n220), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n229), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT65), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(G13), .ZN(new_n251));
  NOR3_X1   g0051(.A1(new_n251), .A2(new_n211), .A3(G1), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n202), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n219), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n255), .B1(new_n210), .B2(G20), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n253), .B1(new_n257), .B2(new_n202), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT8), .B(G58), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT66), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n259), .B(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n211), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n258), .B1(new_n267), .B2(new_n255), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT9), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n268), .B(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT10), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(KEYINPUT70), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G1), .A3(G13), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  OR2_X1    g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AND2_X1   g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NOR2_X1   g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI22_X1  g0081(.A1(new_n278), .A2(G223), .B1(new_n281), .B2(G77), .ZN(new_n282));
  AOI21_X1  g0082(.A(G1698), .B1(new_n276), .B2(new_n277), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G222), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n274), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G41), .ZN(new_n286));
  INV_X1    g0086(.A(G45), .ZN(new_n287));
  AOI21_X1  g0087(.A(G1), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n288), .A2(new_n274), .A3(G274), .ZN(new_n289));
  INV_X1    g0089(.A(G226), .ZN(new_n290));
  AND2_X1   g0090(.A1(G33), .A2(G41), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G41), .A2(G45), .ZN(new_n292));
  OAI22_X1  g0092(.A1(new_n291), .A2(new_n219), .B1(new_n292), .B2(G1), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n289), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n285), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n272), .B1(new_n295), .B2(G190), .ZN(new_n296));
  INV_X1    g0096(.A(G200), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT69), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NOR3_X1   g0098(.A1(new_n295), .A2(KEYINPUT69), .A3(new_n297), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n270), .A2(new_n296), .A3(new_n298), .A4(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n271), .A2(KEYINPUT70), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n301), .B(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  INV_X1    g0104(.A(new_n295), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n268), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(G179), .B2(new_n305), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n290), .A2(G1698), .ZN(new_n309));
  OAI221_X1 g0109(.A(new_n309), .B1(G223), .B2(G1698), .C1(new_n279), .C2(new_n280), .ZN(new_n310));
  NAND2_X1  g0110(.A1(G33), .A2(G87), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n274), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n289), .B1(new_n229), .B2(new_n293), .ZN(new_n313));
  INV_X1    g0113(.A(G190), .ZN(new_n314));
  NOR3_X1   g0114(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n312), .A2(new_n313), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n315), .B1(new_n317), .B2(G200), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n259), .B(KEYINPUT66), .ZN(new_n319));
  INV_X1    g0119(.A(new_n252), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n261), .A2(new_n257), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n228), .A2(new_n222), .ZN(new_n324));
  OAI21_X1  g0124(.A(G20), .B1(new_n324), .B2(new_n201), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n265), .A2(G159), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(KEYINPUT7), .B1(new_n281), .B2(new_n211), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n276), .A2(KEYINPUT7), .A3(new_n211), .A4(new_n277), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(G68), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT75), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n327), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n276), .A2(new_n211), .A3(new_n277), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT7), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n222), .B1(new_n336), .B2(new_n329), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT75), .ZN(new_n338));
  AOI21_X1  g0138(.A(KEYINPUT16), .B1(new_n333), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n327), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n331), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT16), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n255), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n318), .B(new_n323), .C1(new_n339), .C2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT17), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n344), .B(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n323), .B1(new_n339), .B2(new_n343), .ZN(new_n347));
  INV_X1    g0147(.A(G179), .ZN(new_n348));
  NOR3_X1   g0148(.A1(new_n312), .A2(new_n313), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n349), .B1(new_n317), .B2(G169), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(KEYINPUT18), .B1(new_n347), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n347), .A2(KEYINPUT18), .A3(new_n351), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n352), .B1(KEYINPUT76), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n340), .B1(new_n337), .B2(KEYINPUT75), .ZN(new_n355));
  AOI211_X1 g0155(.A(new_n332), .B(new_n222), .C1(new_n336), .C2(new_n329), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n342), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n255), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n337), .A2(new_n327), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n358), .B1(new_n359), .B2(KEYINPUT16), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n350), .B1(new_n361), .B2(new_n323), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT76), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(new_n363), .A3(KEYINPUT18), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n346), .B1(new_n354), .B2(new_n364), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n320), .A2(KEYINPUT12), .A3(G68), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT12), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n252), .B2(new_n222), .ZN(new_n368));
  OAI22_X1  g0168(.A1(new_n366), .A2(new_n368), .B1(new_n257), .B2(new_n222), .ZN(new_n369));
  INV_X1    g0169(.A(new_n265), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n370), .A2(new_n202), .B1(new_n211), .B2(G68), .ZN(new_n371));
  INV_X1    g0171(.A(G77), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n262), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n255), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT11), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n369), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n375), .B2(new_n374), .ZN(new_n378));
  NOR2_X1   g0178(.A1(G226), .A2(G1698), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(new_n229), .B2(G1698), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n276), .A2(new_n277), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n380), .A2(new_n381), .B1(G33), .B2(G97), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n289), .B1(new_n382), .B2(new_n274), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT71), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n293), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n274), .B(KEYINPUT71), .C1(G1), .C2(new_n292), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n385), .A2(G238), .A3(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT13), .B1(new_n383), .B2(new_n387), .ZN(new_n388));
  AND3_X1   g0188(.A1(new_n288), .A2(new_n274), .A3(G274), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n290), .A2(new_n275), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n229), .A2(G1698), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n390), .B(new_n391), .C1(new_n279), .C2(new_n280), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G97), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n291), .A2(new_n219), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n389), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT13), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n385), .A2(G238), .A3(new_n386), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n297), .B1(new_n388), .B2(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n397), .A2(KEYINPUT72), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n383), .B2(new_n387), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n396), .A2(new_n398), .A3(new_n401), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n314), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NOR3_X1   g0205(.A1(new_n378), .A2(new_n400), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n304), .B1(new_n388), .B2(new_n399), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT14), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n407), .A2(KEYINPUT74), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n348), .B1(new_n403), .B2(new_n404), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n394), .A2(new_n395), .ZN(new_n411));
  AND4_X1   g0211(.A1(new_n397), .A2(new_n398), .A3(new_n411), .A4(new_n289), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n397), .B1(new_n396), .B2(new_n398), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n408), .B(G169), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT74), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n410), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NOR3_X1   g0216(.A1(new_n407), .A2(KEYINPUT73), .A3(new_n408), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT73), .ZN(new_n418));
  OAI21_X1  g0218(.A(G169), .B1(new_n412), .B2(new_n413), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n418), .B1(new_n419), .B2(KEYINPUT14), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n409), .B(new_n416), .C1(new_n417), .C2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n406), .B1(new_n421), .B2(new_n378), .ZN(new_n422));
  OAI22_X1  g0222(.A1(new_n259), .A2(new_n370), .B1(new_n211), .B2(new_n372), .ZN(new_n423));
  XNOR2_X1  g0223(.A(KEYINPUT15), .B(G87), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n424), .A2(new_n262), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n255), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT67), .ZN(new_n427));
  XNOR2_X1  g0227(.A(new_n426), .B(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n320), .A2(G77), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(new_n256), .B2(G77), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT68), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n428), .A2(KEYINPUT68), .A3(new_n430), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(G244), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n289), .B1(new_n436), .B2(new_n293), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n283), .A2(G232), .B1(new_n281), .B2(G107), .ZN(new_n438));
  INV_X1    g0238(.A(new_n278), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n438), .B1(new_n223), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n437), .B1(new_n440), .B2(new_n395), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(G190), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n442), .B1(new_n297), .B2(new_n441), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n435), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n441), .A2(new_n348), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n445), .B1(G169), .B2(new_n441), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n446), .B1(new_n433), .B2(new_n434), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n308), .A2(new_n365), .A3(new_n422), .A4(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n287), .A2(G1), .ZN(new_n450));
  AND2_X1   g0250(.A1(KEYINPUT5), .A2(G41), .ZN(new_n451));
  NOR2_X1   g0251(.A1(KEYINPUT5), .A2(G41), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n453), .A2(G264), .A3(new_n274), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT5), .B(G41), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n455), .A2(G274), .A3(new_n274), .A4(new_n450), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n225), .A2(G1698), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(new_n279), .B2(new_n280), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT87), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT87), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n381), .A2(new_n461), .A3(new_n458), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  OAI211_X1 g0263(.A(G257), .B(G1698), .C1(new_n279), .C2(new_n280), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT86), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT86), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n464), .A2(new_n467), .B1(G33), .B2(G294), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n463), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n457), .B1(new_n469), .B2(new_n395), .ZN(new_n470));
  OAI21_X1  g0270(.A(KEYINPUT88), .B1(new_n470), .B2(new_n304), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT88), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n460), .A2(new_n462), .B1(new_n465), .B2(KEYINPUT86), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n274), .B1(new_n473), .B2(new_n468), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n472), .B(G169), .C1(new_n474), .C2(new_n457), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n470), .A2(G179), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n471), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT89), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT23), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n479), .B1(new_n211), .B2(G107), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n207), .A2(KEYINPUT23), .A3(G20), .ZN(new_n481));
  NAND2_X1  g0281(.A1(G33), .A2(G116), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n480), .A2(new_n481), .B1(new_n483), .B2(new_n211), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n381), .A2(new_n211), .A3(G87), .ZN(new_n485));
  AND2_X1   g0285(.A1(new_n485), .A2(KEYINPUT22), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n485), .A2(KEYINPUT22), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT24), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT24), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n490), .B(new_n484), .C1(new_n486), .C2(new_n487), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n358), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n252), .A2(new_n207), .ZN(new_n493));
  OR2_X1    g0293(.A1(new_n493), .A2(KEYINPUT85), .ZN(new_n494));
  XNOR2_X1  g0294(.A(KEYINPUT84), .B(KEYINPUT25), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n495), .B1(new_n493), .B2(KEYINPUT85), .ZN(new_n496));
  OR2_X1    g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n494), .A2(new_n496), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n210), .A2(G33), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n320), .A2(new_n358), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G107), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n497), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n492), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT89), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n471), .A2(new_n475), .A3(new_n505), .A4(new_n476), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n478), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT90), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT82), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n453), .A2(new_n509), .A3(G270), .A4(new_n274), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n510), .A2(new_n456), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n453), .A2(G270), .A3(new_n274), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT82), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT83), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n278), .A2(new_n515), .A3(G264), .ZN(new_n516));
  OAI211_X1 g0316(.A(G264), .B(G1698), .C1(new_n279), .C2(new_n280), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(KEYINPUT83), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(G257), .B(new_n275), .C1(new_n279), .C2(new_n280), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n276), .A2(G303), .A3(new_n277), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n274), .B1(new_n519), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n514), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(G116), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n254), .A2(new_n219), .B1(G20), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(G20), .B1(G33), .B2(G283), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(G33), .B2(new_n206), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT20), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n527), .A2(new_n529), .A3(KEYINPUT20), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n252), .A2(new_n526), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n320), .A2(new_n358), .A3(new_n499), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n536), .B1(new_n537), .B2(new_n526), .ZN(new_n538));
  OAI21_X1  g0338(.A(G169), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(KEYINPUT21), .B1(new_n525), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n522), .B1(new_n516), .B2(new_n518), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n511), .B(new_n513), .C1(new_n541), .C2(new_n274), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n534), .B(new_n536), .C1(new_n526), .C2(new_n537), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT21), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n542), .A2(new_n543), .A3(new_n544), .A4(G169), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(G244), .B(G1698), .C1(new_n279), .C2(new_n280), .ZN(new_n547));
  OAI211_X1 g0347(.A(G238), .B(new_n275), .C1(new_n279), .C2(new_n280), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n547), .A2(new_n548), .A3(new_n482), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n395), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n210), .A2(G45), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n274), .A2(G250), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n274), .A2(G274), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n552), .B1(new_n553), .B2(new_n551), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n556), .A2(new_n314), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n500), .A2(G87), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n424), .A2(new_n252), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n211), .B(G68), .C1(new_n279), .C2(new_n280), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT19), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(new_n262), .B2(new_n206), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n211), .B1(new_n393), .B2(new_n561), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n224), .A2(new_n206), .A3(new_n207), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT80), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n564), .A2(KEYINPUT80), .A3(new_n565), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n563), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n558), .B(new_n559), .C1(new_n570), .C2(new_n358), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n557), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n556), .A2(G200), .ZN(new_n573));
  AOI21_X1  g0373(.A(G169), .B1(new_n550), .B2(new_n555), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n554), .B1(new_n395), .B2(new_n549), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n574), .B1(new_n348), .B2(new_n575), .ZN(new_n576));
  XOR2_X1   g0376(.A(new_n424), .B(KEYINPUT81), .Z(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n500), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n578), .B(new_n559), .C1(new_n570), .C2(new_n358), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n572), .A2(new_n573), .B1(new_n576), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n524), .A2(new_n348), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n513), .A2(new_n456), .A3(new_n510), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(new_n582), .A3(new_n543), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n543), .B1(new_n542), .B2(G200), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n314), .B2(new_n542), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n546), .A2(new_n580), .A3(new_n583), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n453), .A2(new_n274), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n456), .B1(new_n587), .B2(new_n230), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n278), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n589));
  OAI211_X1 g0389(.A(G244), .B(new_n275), .C1(new_n279), .C2(new_n280), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT4), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n591), .A2(G1698), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n593), .B(G244), .C1(new_n280), .C2(new_n279), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT78), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT78), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n381), .A2(new_n596), .A3(G244), .A4(new_n593), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n589), .A2(new_n592), .A3(new_n595), .A4(new_n597), .ZN(new_n598));
  AOI211_X1 g0398(.A(new_n314), .B(new_n588), .C1(new_n598), .C2(new_n395), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n265), .A2(G77), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT6), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT77), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT77), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(KEYINPUT6), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n207), .A2(G97), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(G97), .A2(G107), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n208), .A2(new_n602), .A3(new_n604), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n600), .B1(new_n610), .B2(new_n211), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n207), .B1(new_n336), .B2(new_n329), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n255), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n320), .A2(G97), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n500), .B2(G97), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n599), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n598), .A2(new_n395), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT79), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n598), .A2(KEYINPUT79), .A3(new_n395), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n588), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n617), .B1(new_n622), .B2(new_n297), .ZN(new_n623));
  INV_X1    g0423(.A(new_n588), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n598), .A2(KEYINPUT79), .A3(new_n395), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT79), .B1(new_n598), .B2(new_n395), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n348), .B(new_n624), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n588), .B1(new_n598), .B2(new_n395), .ZN(new_n628));
  OR2_X1    g0428(.A1(new_n628), .A2(G169), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n627), .A2(new_n629), .A3(new_n616), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n623), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n586), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT90), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n478), .A2(new_n504), .A3(new_n633), .A4(new_n506), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n470), .A2(G190), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n503), .B(new_n635), .C1(new_n297), .C2(new_n470), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n508), .A2(new_n632), .A3(new_n634), .A4(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n449), .A2(new_n637), .ZN(G372));
  NAND2_X1  g0438(.A1(new_n421), .A2(new_n378), .ZN(new_n639));
  INV_X1    g0439(.A(new_n447), .ZN(new_n640));
  AOI211_X1 g0440(.A(new_n406), .B(new_n346), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT18), .ZN(new_n642));
  INV_X1    g0442(.A(new_n323), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n643), .B1(new_n357), .B2(new_n360), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n642), .B1(new_n644), .B2(new_n350), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n645), .A2(new_n353), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n303), .B1(new_n641), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n307), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n631), .ZN(new_n650));
  INV_X1    g0450(.A(new_n574), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n575), .A2(new_n348), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n579), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT91), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n575), .B2(new_n297), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n556), .A2(KEYINPUT91), .A3(G200), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n570), .A2(new_n358), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n575), .A2(G190), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n658), .A2(new_n659), .A3(new_n559), .A4(new_n558), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n653), .B1(new_n657), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT92), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n653), .B(KEYINPUT92), .C1(new_n660), .C2(new_n657), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n650), .A2(new_n636), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n546), .A2(new_n583), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT93), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n504), .A2(new_n477), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n666), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n627), .A2(new_n629), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT94), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n672), .A2(new_n673), .B1(new_n613), .B2(new_n615), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n627), .A2(KEYINPUT94), .A3(new_n629), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n665), .A2(new_n674), .A3(new_n675), .A4(new_n676), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n580), .A2(new_n629), .A3(new_n627), .A4(new_n616), .ZN(new_n678));
  AOI22_X1  g0478(.A1(new_n678), .A2(KEYINPUT26), .B1(new_n579), .B2(new_n576), .ZN(new_n679));
  AND3_X1   g0479(.A1(new_n677), .A2(new_n679), .A3(KEYINPUT95), .ZN(new_n680));
  AOI21_X1  g0480(.A(KEYINPUT95), .B1(new_n677), .B2(new_n679), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n671), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n649), .B1(new_n683), .B2(new_n449), .ZN(G369));
  NAND3_X1  g0484(.A1(new_n210), .A2(new_n211), .A3(G13), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(G213), .A3(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(G343), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n668), .A2(new_n543), .A3(new_n690), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n546), .A2(new_n583), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n543), .A2(new_n690), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(new_n585), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G330), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n508), .A2(new_n634), .ZN(new_n698));
  INV_X1    g0498(.A(new_n690), .ZN(new_n699));
  OAI211_X1 g0499(.A(new_n698), .B(new_n636), .C1(new_n503), .C2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n507), .B2(new_n699), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n670), .A2(new_n699), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n692), .A2(new_n690), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n698), .A2(new_n636), .A3(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(G399));
  INV_X1    g0506(.A(new_n214), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G41), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n565), .A2(G116), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(G1), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n218), .B2(new_n709), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT28), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT29), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n682), .A2(new_n714), .A3(new_n699), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n508), .A2(new_n634), .A3(new_n692), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(KEYINPUT97), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT97), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n508), .A2(new_n718), .A3(new_n634), .A4(new_n692), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n717), .A2(new_n666), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n653), .B1(new_n678), .B2(KEYINPUT26), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n665), .A2(new_n676), .A3(new_n674), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n721), .B1(new_n722), .B2(KEYINPUT26), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n690), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n715), .B1(new_n724), .B2(new_n714), .ZN(new_n725));
  INV_X1    g0525(.A(G330), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n698), .A2(new_n636), .A3(new_n632), .A4(new_n699), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT96), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n575), .A2(G179), .ZN(new_n729));
  OAI211_X1 g0529(.A(new_n542), .B(new_n729), .C1(new_n474), .C2(new_n457), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n728), .B1(new_n622), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n556), .A2(new_n348), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n470), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n732), .A2(KEYINPUT96), .A3(new_n542), .A4(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n469), .A2(new_n395), .ZN(new_n736));
  AND4_X1   g0536(.A1(new_n736), .A2(new_n582), .A3(new_n454), .A4(new_n575), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n737), .A2(KEYINPUT30), .A3(new_n628), .A4(new_n581), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT30), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n581), .A2(new_n628), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n736), .A2(new_n582), .A3(new_n454), .A4(new_n575), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n731), .A2(new_n735), .A3(new_n738), .A4(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(KEYINPUT31), .B1(new_n743), .B2(new_n690), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n738), .B(new_n742), .C1(new_n622), .C2(new_n730), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n690), .A2(KEYINPUT31), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n726), .B1(new_n727), .B2(new_n748), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n725), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n713), .B1(new_n751), .B2(G1), .ZN(G364));
  NOR2_X1   g0552(.A1(new_n695), .A2(G330), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT98), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n251), .A2(G20), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n210), .B1(new_n755), .B2(G45), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n754), .B1(new_n708), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n709), .A2(KEYINPUT98), .A3(new_n756), .ZN(new_n759));
  AOI211_X1 g0559(.A(new_n753), .B(new_n697), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G13), .A2(G33), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n219), .B1(G20), .B2(new_n304), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n246), .A2(G45), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n707), .A2(new_n381), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n767), .B(new_n768), .C1(G45), .C2(new_n218), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n707), .A2(new_n281), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n770), .A2(G355), .B1(new_n526), .B2(new_n707), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n766), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n764), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n211), .A2(new_n348), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G200), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n314), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT32), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n211), .A2(G179), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G190), .A2(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G159), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n777), .A2(new_n202), .B1(new_n778), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n775), .A2(G190), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n784), .B1(G68), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n774), .A2(new_n780), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n381), .B1(new_n787), .B2(new_n372), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n774), .A2(G190), .A3(new_n297), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n788), .B1(G58), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n779), .A2(G190), .A3(G200), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n224), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n314), .A2(G179), .A3(G200), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n211), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n793), .B1(G97), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n779), .A2(new_n314), .A3(G200), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n778), .A2(new_n783), .B1(new_n799), .B2(G107), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n786), .A2(new_n791), .A3(new_n797), .A4(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G322), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n789), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G311), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n281), .B1(new_n787), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n781), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n803), .B(new_n805), .C1(G329), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n776), .A2(G326), .ZN(new_n808));
  XNOR2_X1  g0608(.A(KEYINPUT33), .B(G317), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G294), .A2(new_n796), .B1(new_n785), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n792), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n811), .A2(G303), .B1(new_n799), .B2(G283), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n807), .A2(new_n808), .A3(new_n810), .A4(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n773), .B1(new_n801), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n759), .A2(new_n758), .ZN(new_n815));
  NOR3_X1   g0615(.A1(new_n772), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n763), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n816), .B1(new_n695), .B2(new_n817), .ZN(new_n818));
  XOR2_X1   g0618(.A(new_n818), .B(KEYINPUT99), .Z(new_n819));
  NOR2_X1   g0619(.A1(new_n760), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(G396));
  NAND2_X1  g0621(.A1(new_n435), .A2(new_n690), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n441), .A2(G169), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(new_n348), .B2(new_n441), .ZN(new_n824));
  AOI21_X1  g0624(.A(KEYINPUT68), .B1(new_n428), .B2(new_n430), .ZN(new_n825));
  INV_X1    g0625(.A(new_n434), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n824), .B(new_n690), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(KEYINPUT101), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT101), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n447), .A2(new_n829), .A3(new_n690), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n448), .A2(new_n822), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n683), .B2(new_n690), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n828), .A2(new_n830), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n640), .B(new_n822), .C1(new_n435), .C2(new_n443), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n682), .A2(new_n699), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n832), .A2(new_n749), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n815), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT102), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n832), .A2(new_n836), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n841), .A2(new_n749), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n837), .A2(KEYINPUT102), .A3(new_n815), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n840), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n764), .A2(new_n761), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n846), .A2(G77), .ZN(new_n847));
  INV_X1    g0647(.A(G303), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n777), .A2(new_n848), .B1(new_n798), .B2(new_n224), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(G107), .B2(new_n811), .ZN(new_n850));
  INV_X1    g0650(.A(G294), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n789), .A2(new_n851), .B1(new_n781), .B2(new_n804), .ZN(new_n852));
  INV_X1    g0652(.A(new_n787), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n381), .B(new_n852), .C1(G116), .C2(new_n853), .ZN(new_n854));
  AOI22_X1  g0654(.A1(G97), .A2(new_n796), .B1(new_n785), .B2(G283), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n850), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(G132), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n381), .B1(new_n781), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(G68), .B2(new_n799), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n796), .A2(G58), .B1(new_n811), .B2(G50), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n790), .A2(G143), .B1(new_n853), .B2(G159), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n776), .A2(G137), .ZN(new_n862));
  INV_X1    g0662(.A(G150), .ZN(new_n863));
  INV_X1    g0663(.A(new_n785), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n861), .B(new_n862), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  XNOR2_X1  g0665(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n859), .B(new_n860), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n865), .A2(new_n866), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n856), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n815), .B(new_n847), .C1(new_n869), .C2(new_n764), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n835), .B2(new_n762), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n844), .A2(new_n871), .ZN(G384));
  NOR2_X1   g0672(.A1(new_n755), .A2(new_n210), .ZN(new_n873));
  INV_X1    g0673(.A(new_n449), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n725), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n649), .ZN(new_n876));
  XOR2_X1   g0676(.A(new_n876), .B(KEYINPUT105), .Z(new_n877));
  OAI211_X1 g0677(.A(new_n378), .B(new_n690), .C1(new_n421), .C2(new_n406), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n378), .A2(new_n690), .ZN(new_n880));
  AOI211_X1 g0680(.A(new_n406), .B(new_n880), .C1(new_n421), .C2(new_n378), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n640), .A2(new_n690), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n882), .B1(new_n836), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n359), .A2(KEYINPUT16), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n323), .B1(new_n343), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n688), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n353), .A2(KEYINPUT76), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n891), .A2(new_n364), .A3(new_n645), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n344), .B(KEYINPUT17), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n890), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT103), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT37), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n344), .A2(new_n896), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n361), .A2(new_n323), .B1(new_n350), .B2(new_n688), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n895), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n350), .A2(new_n688), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n347), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n901), .A2(KEYINPUT103), .A3(new_n896), .A4(new_n344), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n900), .A2(new_n888), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n344), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n899), .A2(new_n902), .B1(KEYINPUT37), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n886), .B1(new_n894), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n899), .A2(new_n902), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n904), .A2(KEYINPUT37), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n909), .B(KEYINPUT38), .C1(new_n365), .C2(new_n890), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n885), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n646), .A2(new_n688), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n639), .A2(new_n690), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT104), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n344), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n901), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n344), .A2(new_n916), .ZN(new_n919));
  OAI21_X1  g0719(.A(KEYINPUT37), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n907), .A2(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n347), .B(new_n889), .C1(new_n646), .C2(new_n346), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT38), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n910), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT39), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n911), .B2(new_n926), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n912), .B(new_n913), .C1(new_n915), .C2(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n877), .B(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n743), .A2(KEYINPUT31), .A3(new_n690), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n932), .A2(new_n744), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n637), .B2(new_n690), .ZN(new_n934));
  INV_X1    g0734(.A(new_n880), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n422), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n831), .B1(new_n936), .B2(new_n878), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n894), .A2(new_n886), .A3(new_n905), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n934), .B(new_n937), .C1(new_n938), .C2(new_n923), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n835), .B1(new_n879), .B2(new_n881), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(new_n727), .B2(new_n933), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT40), .B1(new_n906), .B2(new_n910), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n939), .A2(KEYINPUT40), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n449), .B1(new_n727), .B2(new_n933), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n726), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n945), .B2(new_n944), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n873), .B1(new_n931), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n931), .B2(new_n947), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n219), .A2(new_n211), .A3(new_n526), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT35), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n950), .B1(new_n610), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(new_n951), .B2(new_n610), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT36), .Z(new_n954));
  NOR3_X1   g0754(.A1(new_n218), .A2(new_n372), .A3(new_n324), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n222), .A2(G50), .ZN(new_n956));
  OAI211_X1 g0756(.A(G1), .B(new_n251), .C1(new_n955), .C2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n949), .A2(new_n954), .A3(new_n957), .ZN(G367));
  INV_X1    g0758(.A(new_n815), .ZN(new_n959));
  AND2_X1   g0759(.A1(new_n768), .A2(new_n241), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n765), .B1(new_n214), .B2(new_n424), .ZN(new_n961));
  INV_X1    g0761(.A(G143), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n962), .A2(new_n777), .B1(new_n864), .B2(new_n782), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n381), .B1(new_n789), .B2(new_n863), .ZN(new_n964));
  XNOR2_X1  g0764(.A(KEYINPUT108), .B(G137), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n787), .A2(new_n202), .B1(new_n781), .B2(new_n965), .ZN(new_n966));
  NOR3_X1   g0766(.A1(new_n963), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n798), .A2(new_n372), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(G58), .B2(new_n811), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n967), .B(new_n969), .C1(new_n222), .C2(new_n795), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n798), .A2(new_n206), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(G294), .B2(new_n785), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n972), .B1(new_n207), .B2(new_n795), .C1(new_n804), .C2(new_n777), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n790), .A2(G303), .B1(new_n806), .B2(G317), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT46), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n792), .B2(new_n526), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n811), .A2(KEYINPUT46), .A3(G116), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n381), .B1(new_n853), .B2(G283), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n974), .A2(new_n976), .A3(new_n977), .A4(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n970), .B1(new_n973), .B2(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT47), .Z(new_n981));
  OAI221_X1 g0781(.A(new_n959), .B1(new_n960), .B2(new_n961), .C1(new_n981), .C2(new_n773), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT109), .Z(new_n983));
  NAND2_X1  g0783(.A1(new_n571), .A2(new_n690), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n665), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n653), .B2(new_n984), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n983), .B1(new_n817), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n631), .B1(new_n616), .B2(new_n690), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n674), .A2(new_n676), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n988), .B1(new_n989), .B2(new_n690), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n705), .A2(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT42), .Z(new_n992));
  OAI21_X1  g0792(.A(new_n630), .B1(new_n990), .B2(new_n698), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n992), .B1(new_n699), .B2(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n986), .B(KEYINPUT43), .ZN(new_n995));
  OR3_X1    g0795(.A1(new_n994), .A2(KEYINPUT106), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(KEYINPUT106), .B1(new_n994), .B2(new_n995), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n994), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n996), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n702), .A2(new_n990), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1000), .B(new_n1001), .Z(new_n1002));
  NAND2_X1  g0802(.A1(new_n705), .A2(new_n703), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n990), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT44), .Z(new_n1005));
  NOR2_X1   g0805(.A1(new_n1003), .A2(new_n990), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT45), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(new_n702), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n705), .B1(new_n701), .B2(new_n704), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(new_n696), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n751), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT107), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1012), .A2(KEYINPUT107), .A3(new_n751), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1009), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n751), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n708), .B(KEYINPUT41), .Z(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n757), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n987), .B1(new_n1002), .B2(new_n1021), .ZN(G387));
  NAND2_X1  g0822(.A1(new_n1011), .A2(new_n750), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1013), .A2(new_n1023), .A3(new_n708), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n701), .A2(new_n817), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n710), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n770), .A2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(G107), .B2(new_n214), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n238), .A2(new_n287), .ZN(new_n1029));
  AOI211_X1 g0829(.A(G45), .B(new_n1026), .C1(G68), .C2(G77), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n259), .A2(G50), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT50), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n707), .B(new_n381), .C1(new_n1030), .C2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1028), .B1(new_n1029), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n959), .B1(new_n1034), .B2(new_n766), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n789), .A2(new_n202), .B1(new_n781), .B2(new_n863), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n281), .B(new_n1036), .C1(G68), .C2(new_n853), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n792), .A2(new_n372), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n971), .B(new_n1038), .C1(G159), .C2(new_n776), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n261), .A2(new_n785), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n577), .A2(new_n796), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1037), .A2(new_n1039), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT110), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n796), .A2(G283), .B1(new_n811), .B2(G294), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n790), .A2(G317), .B1(new_n853), .B2(G303), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n777), .B2(new_n802), .C1(new_n804), .C2(new_n864), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT48), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1044), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT111), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1049), .A2(KEYINPUT49), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n381), .B1(new_n806), .B2(G326), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1051), .B(new_n1052), .C1(new_n526), .C2(new_n798), .ZN(new_n1053));
  AOI21_X1  g0853(.A(KEYINPUT49), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1043), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1035), .B1(new_n1055), .B2(new_n764), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT112), .Z(new_n1057));
  AOI22_X1  g0857(.A1(new_n1012), .A2(new_n757), .B1(new_n1025), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1024), .A2(new_n1058), .ZN(G393));
  AOI22_X1  g0859(.A1(G317), .A2(new_n776), .B1(new_n790), .B2(G311), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT52), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n281), .B1(new_n781), .B2(new_n802), .C1(new_n851), .C2(new_n787), .ZN(new_n1062));
  INV_X1    g0862(.A(G283), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n207), .A2(new_n798), .B1(new_n792), .B2(new_n1063), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n864), .A2(new_n848), .B1(new_n526), .B2(new_n795), .ZN(new_n1065));
  OR4_X1    g0865(.A1(new_n1061), .A2(new_n1062), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n777), .A2(new_n863), .B1(new_n782), .B2(new_n789), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT51), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n381), .B1(new_n781), .B2(new_n962), .C1(new_n259), .C2(new_n787), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n785), .A2(G50), .B1(new_n799), .B2(G87), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n795), .A2(new_n372), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(G68), .B2(new_n811), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1068), .A2(new_n1070), .A3(new_n1071), .A4(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n773), .B1(new_n1066), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n765), .B1(new_n206), .B2(new_n214), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n768), .B2(new_n249), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n1075), .A2(new_n815), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n990), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1078), .B1(new_n1079), .B2(new_n817), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n702), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1008), .B(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1080), .B1(new_n1082), .B2(new_n756), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n709), .B1(new_n1082), .B2(new_n1013), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1083), .B1(new_n1017), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(G390));
  INV_X1    g0886(.A(KEYINPUT114), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n726), .B1(new_n727), .B2(new_n933), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n937), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n748), .B1(new_n637), .B2(new_n690), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1090), .A2(G330), .A3(new_n835), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n882), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1089), .A2(new_n1092), .B1(new_n836), .B2(new_n884), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n690), .B(new_n831), .C1(new_n720), .C2(new_n723), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1091), .A2(new_n882), .ZN(new_n1095));
  NOR3_X1   g0895(.A1(new_n1094), .A2(new_n1095), .A3(new_n883), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n835), .B1(new_n1088), .B2(KEYINPUT113), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n934), .A2(G330), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT113), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n882), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1093), .B1(new_n1096), .B2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n449), .A2(new_n1098), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n875), .A2(new_n649), .A3(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1087), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1093), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n883), .B1(new_n724), .B2(new_n835), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1095), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n882), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n831), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1088), .A2(KEYINPUT113), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1107), .B1(new_n1110), .B2(new_n1114), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n648), .B(new_n1103), .C1(new_n725), .C2(new_n874), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1115), .A2(new_n1116), .A3(KEYINPUT114), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1106), .A2(new_n1117), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n915), .B(new_n925), .C1(new_n1108), .C2(new_n882), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n928), .B1(new_n885), .B2(new_n914), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1119), .A2(new_n1120), .A3(new_n1109), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1089), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n708), .B1(new_n1118), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1118), .A2(new_n1123), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT115), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1118), .A2(KEYINPUT115), .A3(new_n1123), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1124), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1123), .A2(new_n757), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n928), .A2(new_n761), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n792), .A2(new_n863), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT53), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n864), .A2(new_n965), .B1(new_n782), .B2(new_n795), .ZN(new_n1134));
  INV_X1    g0934(.A(G128), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n777), .A2(new_n1135), .B1(new_n798), .B2(new_n202), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(KEYINPUT54), .B(G143), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n381), .B1(new_n787), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(G125), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n789), .A2(new_n857), .B1(new_n781), .B2(new_n1139), .ZN(new_n1140));
  NOR4_X1   g0940(.A1(new_n1134), .A2(new_n1136), .A3(new_n1138), .A4(new_n1140), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n207), .A2(new_n864), .B1(new_n777), .B2(new_n1063), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n281), .B1(new_n787), .B2(new_n206), .C1(new_n526), .C2(new_n789), .ZN(new_n1143));
  NOR4_X1   g0943(.A1(new_n1142), .A2(new_n793), .A3(new_n1072), .A4(new_n1143), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n798), .A2(new_n222), .B1(new_n781), .B2(new_n851), .ZN(new_n1145));
  XOR2_X1   g0945(.A(new_n1145), .B(KEYINPUT116), .Z(new_n1146));
  AOI22_X1  g0946(.A1(new_n1133), .A2(new_n1141), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n959), .B1(new_n261), .B2(new_n846), .C1(new_n1147), .C2(new_n773), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT117), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1130), .B1(new_n1131), .B2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1129), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(G378));
  NAND2_X1  g0952(.A1(new_n303), .A2(new_n307), .ZN(new_n1153));
  XOR2_X1   g0953(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1154));
  XNOR2_X1  g0954(.A(new_n1153), .B(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n268), .A2(new_n688), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT119), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1155), .B(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n761), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n959), .B1(G50), .B2(new_n846), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n1139), .A2(new_n777), .B1(new_n864), .B2(new_n857), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n790), .A2(G128), .B1(new_n853), .B2(G137), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n792), .B2(new_n1137), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1162), .B(new_n1164), .C1(G150), .C2(new_n796), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  OR2_X1    g0966(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n799), .A2(G159), .ZN(new_n1169));
  AOI211_X1 g0969(.A(G33), .B(G41), .C1(new_n806), .C2(G124), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n381), .A2(G41), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1172), .B1(new_n1063), .B2(new_n781), .C1(new_n207), .C2(new_n789), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1038), .B(new_n1173), .C1(G68), .C2(new_n796), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n777), .A2(new_n526), .B1(new_n798), .B2(new_n228), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(G97), .B2(new_n785), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n577), .A2(new_n853), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1174), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  XOR2_X1   g0978(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1172), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1181), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1171), .A2(new_n1180), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1161), .B1(new_n1184), .B2(new_n764), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1160), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT120), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n943), .B2(new_n726), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT40), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n941), .B2(new_n925), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n890), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n363), .B1(new_n362), .B2(KEYINPUT18), .ZN(new_n1192));
  NOR4_X1   g0992(.A1(new_n644), .A2(KEYINPUT76), .A3(new_n642), .A4(new_n350), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1192), .A2(new_n1193), .A3(new_n352), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1191), .B1(new_n1194), .B2(new_n346), .ZN(new_n1195));
  AOI21_X1  g0995(.A(KEYINPUT38), .B1(new_n1195), .B2(new_n909), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1189), .B1(new_n1196), .B2(new_n938), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n934), .A2(new_n937), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  OAI211_X1 g0999(.A(KEYINPUT120), .B(G330), .C1(new_n1190), .C2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1188), .A2(new_n1200), .A3(new_n1159), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1155), .B(new_n1157), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1202), .B(new_n1187), .C1(new_n726), .C2(new_n943), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1201), .A2(new_n929), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(KEYINPUT121), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n929), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  XOR2_X1   g1008(.A(new_n1205), .B(new_n1208), .Z(new_n1209));
  OAI21_X1  g1009(.A(new_n1186), .B1(new_n1209), .B2(new_n756), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n1118), .A2(KEYINPUT115), .A3(new_n1123), .ZN(new_n1212));
  AOI21_X1  g1012(.A(KEYINPUT115), .B1(new_n1118), .B2(new_n1123), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1116), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT122), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1208), .A2(new_n1215), .A3(new_n1204), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1206), .A2(KEYINPUT122), .A3(new_n1207), .ZN(new_n1217));
  AND3_X1   g1017(.A1(new_n1216), .A2(KEYINPUT57), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1214), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n708), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1205), .B(new_n1208), .ZN(new_n1221));
  AOI21_X1  g1021(.A(KEYINPUT57), .B1(new_n1214), .B2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1211), .B1(new_n1220), .B2(new_n1222), .ZN(G375));
  NAND2_X1  g1023(.A1(new_n882), .A2(new_n761), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n864), .A2(new_n1137), .B1(new_n228), .B2(new_n798), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n381), .B1(new_n789), .B2(new_n965), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n787), .A2(new_n863), .B1(new_n781), .B2(new_n1135), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(G50), .A2(new_n796), .B1(new_n776), .B2(G132), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1228), .B(new_n1229), .C1(new_n782), .C2(new_n792), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n789), .A2(new_n1063), .B1(new_n787), .B2(new_n207), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n381), .B(new_n1231), .C1(G303), .C2(new_n806), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n968), .B1(G97), .B2(new_n811), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(G116), .A2(new_n785), .B1(new_n776), .B2(G294), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1232), .A2(new_n1041), .A3(new_n1233), .A4(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n773), .B1(new_n1230), .B2(new_n1235), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n815), .B(new_n1236), .C1(new_n222), .C2(new_n845), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1115), .A2(new_n757), .B1(new_n1224), .B2(new_n1237), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT123), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1239), .B(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1106), .A2(new_n1117), .A3(new_n1020), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1238), .B1(new_n1241), .B2(new_n1242), .ZN(G381));
  NAND3_X1  g1043(.A1(new_n1024), .A2(new_n820), .A3(new_n1058), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1244), .A2(G384), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT124), .ZN(new_n1246));
  NOR4_X1   g1046(.A1(G387), .A2(new_n1246), .A3(G390), .A4(G381), .ZN(new_n1247));
  XOR2_X1   g1047(.A(new_n1247), .B(KEYINPUT125), .Z(new_n1248));
  INV_X1    g1048(.A(KEYINPUT57), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1105), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1249), .B1(new_n1250), .B2(new_n1209), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n709), .B1(new_n1214), .B2(new_n1218), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1210), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1151), .ZN(new_n1254));
  OR2_X1    g1054(.A1(new_n1248), .A2(new_n1254), .ZN(G407));
  INV_X1    g1055(.A(new_n1254), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n689), .A2(G213), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1257), .B(KEYINPUT126), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1256), .A2(new_n1258), .ZN(new_n1259));
  OAI211_X1 g1059(.A(G213), .B(new_n1259), .C1(new_n1248), .C2(new_n1254), .ZN(G409));
  NAND3_X1  g1060(.A1(new_n1216), .A2(new_n757), .A3(new_n1217), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1186), .ZN(new_n1262));
  NOR3_X1   g1062(.A1(new_n1129), .A2(new_n1262), .A3(new_n1150), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1214), .A2(new_n1020), .A3(new_n1221), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1258), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n1253), .B2(new_n1151), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1239), .A2(KEYINPUT60), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n708), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(new_n1239), .B(KEYINPUT123), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1106), .A2(new_n1117), .A3(KEYINPUT60), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1268), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1238), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n844), .B(new_n871), .C1(new_n1271), .C2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1270), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1241), .A2(new_n1274), .ZN(new_n1275));
  OAI211_X1 g1075(.A(G384), .B(new_n1238), .C1(new_n1275), .C2(new_n1268), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1258), .A2(G2897), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1273), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1277), .B1(new_n1273), .B2(new_n1276), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(KEYINPUT61), .B1(new_n1266), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1273), .A2(new_n1276), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1265), .B(new_n1283), .C1(new_n1253), .C2(new_n1151), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(KEYINPUT62), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(G375), .A2(G378), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT62), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1286), .A2(new_n1287), .A3(new_n1283), .A4(new_n1265), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1281), .A2(new_n1285), .A3(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1244), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n820), .B1(new_n1024), .B2(new_n1058), .ZN(new_n1291));
  OR3_X1    g1091(.A1(new_n1085), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1085), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(G387), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT127), .ZN(new_n1296));
  OR2_X1    g1096(.A1(new_n1002), .A2(new_n1021), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1297), .A2(new_n987), .A3(new_n1292), .A4(new_n1293), .ZN(new_n1298));
  AND3_X1   g1098(.A1(new_n1295), .A2(new_n1296), .A3(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1296), .B1(new_n1295), .B2(new_n1298), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1289), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT63), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1284), .A2(new_n1303), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1286), .A2(KEYINPUT63), .A3(new_n1283), .A4(new_n1265), .ZN(new_n1305));
  AND2_X1   g1105(.A1(new_n1295), .A2(new_n1298), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1281), .A2(new_n1304), .A3(new_n1305), .A4(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1302), .A2(new_n1307), .ZN(G405));
  NOR2_X1   g1108(.A1(new_n1253), .A2(new_n1151), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1283), .B1(new_n1256), .B2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1286), .A2(new_n1254), .A3(new_n1282), .ZN(new_n1311));
  AND3_X1   g1111(.A1(new_n1310), .A2(new_n1306), .A3(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1306), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1312), .A2(new_n1313), .ZN(G402));
endmodule


