//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 0 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 1 1 0 1 1 0 1 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT65), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT65), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G134), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G137), .ZN(new_n194));
  AOI21_X1  g008(.A(KEYINPUT11), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n190), .A2(new_n192), .A3(G137), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT66), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(new_n194), .ZN(new_n198));
  NAND2_X1  g012(.A1(KEYINPUT66), .A2(G137), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT11), .A2(G134), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n198), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n196), .A2(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(G131), .B1(new_n195), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT11), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT65), .B(G134), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G137), .ZN(new_n206));
  INV_X1    g020(.A(G131), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n206), .A2(new_n207), .A3(new_n196), .A4(new_n201), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n203), .A2(new_n208), .ZN(new_n209));
  XOR2_X1   g023(.A(KEYINPUT83), .B(KEYINPUT12), .Z(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT78), .B(G104), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT3), .B1(new_n212), .B2(G107), .ZN(new_n213));
  INV_X1    g027(.A(G101), .ZN(new_n214));
  INV_X1    g028(.A(G104), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT78), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT78), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G104), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(new_n218), .A3(G107), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n220));
  INV_X1    g034(.A(G107), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(G104), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n213), .A2(new_n214), .A3(new_n219), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT81), .B1(new_n221), .B2(G104), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n224), .B1(new_n212), .B2(G107), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n216), .A2(new_n218), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(KEYINPUT81), .A3(new_n221), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n214), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT82), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AOI211_X1 g044(.A(KEYINPUT82), .B(new_n214), .C1(new_n225), .C2(new_n227), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n223), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G146), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G143), .ZN(new_n234));
  INV_X1    g048(.A(G143), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G146), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n234), .A2(KEYINPUT1), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(new_n238), .A3(G128), .ZN(new_n239));
  INV_X1    g053(.A(G128), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n234), .B(new_n236), .C1(KEYINPUT1), .C2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n232), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n242), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n244), .B(new_n223), .C1(new_n230), .C2(new_n231), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n211), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n245), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n209), .A2(KEYINPUT70), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n203), .A2(new_n249), .A3(new_n208), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT12), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n246), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n225), .A2(new_n227), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G101), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT82), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n228), .A2(new_n229), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n260), .A2(KEYINPUT10), .A3(new_n244), .A4(new_n223), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT10), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n245), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT79), .B(KEYINPUT4), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n220), .B1(new_n226), .B2(new_n221), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n219), .A2(new_n222), .ZN(new_n266));
  OAI211_X1 g080(.A(G101), .B(new_n264), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT80), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n213), .A2(new_n219), .A3(new_n222), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT80), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n269), .A2(new_n270), .A3(G101), .A4(new_n264), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT0), .B(G128), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n274), .A2(KEYINPUT64), .A3(new_n237), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT64), .ZN(new_n276));
  XNOR2_X1  g090(.A(G143), .B(G146), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n276), .B1(new_n277), .B2(new_n273), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n277), .A2(KEYINPUT0), .A3(G128), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n275), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT69), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n269), .A2(G101), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(new_n223), .A3(KEYINPUT4), .ZN(new_n284));
  AND3_X1   g098(.A1(new_n275), .A2(new_n278), .A3(new_n279), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(KEYINPUT69), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n272), .A2(new_n282), .A3(new_n284), .A4(new_n286), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n261), .A2(new_n263), .A3(new_n287), .A4(new_n251), .ZN(new_n288));
  XNOR2_X1  g102(.A(G110), .B(G140), .ZN(new_n289));
  INV_X1    g103(.A(G227), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n290), .A2(G953), .ZN(new_n291));
  XOR2_X1   g105(.A(new_n289), .B(new_n291), .Z(new_n292));
  NAND2_X1  g106(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n255), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n261), .A2(new_n263), .A3(new_n287), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n252), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n292), .B1(new_n296), .B2(new_n288), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n187), .B(new_n188), .C1(new_n294), .C2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT85), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT84), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n293), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n288), .A2(KEYINPUT84), .A3(new_n292), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n296), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n292), .ZN(new_n304));
  INV_X1    g118(.A(new_n288), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n304), .B1(new_n255), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n188), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n299), .B1(new_n308), .B2(G469), .ZN(new_n309));
  AOI21_X1  g123(.A(G902), .B1(new_n303), .B2(new_n306), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n310), .A2(KEYINPUT85), .A3(new_n187), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n298), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G475), .ZN(new_n313));
  NOR2_X1   g127(.A1(G237), .A2(G953), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n314), .A2(G143), .A3(G214), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(G143), .B1(new_n314), .B2(G214), .ZN(new_n317));
  OAI21_X1  g131(.A(G131), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n317), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(new_n207), .A3(new_n315), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT17), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n318), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n207), .B1(new_n319), .B2(new_n315), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT17), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT16), .ZN(new_n325));
  INV_X1    g139(.A(G140), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(new_n326), .A3(G125), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(G125), .ZN(new_n328));
  INV_X1    g142(.A(G125), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G140), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n327), .B1(new_n331), .B2(new_n325), .ZN(new_n332));
  OR2_X1    g146(.A1(new_n332), .A2(new_n233), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n233), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n322), .A2(new_n324), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n328), .A2(new_n330), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT75), .B1(new_n336), .B2(new_n233), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n338));
  NOR3_X1   g152(.A1(new_n331), .A2(new_n338), .A3(G146), .ZN(new_n339));
  OAI22_X1  g153(.A1(new_n337), .A2(new_n339), .B1(new_n233), .B2(new_n336), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n323), .A2(KEYINPUT18), .ZN(new_n341));
  NAND2_X1  g155(.A1(KEYINPUT18), .A2(G131), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n319), .A2(new_n315), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n340), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(G113), .B(G122), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n345), .B(new_n215), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n335), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT97), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n346), .B1(new_n335), .B2(new_n344), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(G902), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n349), .A2(new_n351), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n313), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n335), .A2(new_n344), .A3(new_n346), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n318), .A2(new_n320), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n331), .B(KEYINPUT19), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n333), .B(new_n358), .C1(G146), .C2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n346), .B1(new_n360), .B2(new_n344), .ZN(new_n361));
  OAI21_X1  g175(.A(KEYINPUT96), .B1(new_n357), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n344), .ZN(new_n363));
  INV_X1    g177(.A(new_n346), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT96), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n366), .A3(new_n347), .ZN(new_n367));
  NOR2_X1   g181(.A1(G475), .A2(G902), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n362), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT20), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n365), .A2(new_n347), .ZN(new_n371));
  NOR3_X1   g185(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT98), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n356), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  AOI22_X1  g190(.A1(new_n369), .A2(KEYINPUT20), .B1(new_n371), .B2(new_n372), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT98), .B1(new_n377), .B2(new_n355), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G116), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G122), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n380), .A2(G122), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n381), .B1(new_n382), .B2(KEYINPUT14), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n383), .B1(KEYINPUT14), .B2(new_n381), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G107), .ZN(new_n385));
  XNOR2_X1  g199(.A(G116), .B(G122), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n221), .ZN(new_n387));
  XNOR2_X1  g201(.A(G128), .B(G143), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n205), .B(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n385), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n386), .B(new_n221), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n240), .A2(G143), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n240), .A2(G143), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n392), .B1(KEYINPUT13), .B2(new_n393), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n392), .A2(KEYINPUT13), .ZN(new_n395));
  OAI21_X1  g209(.A(G134), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n205), .A2(new_n388), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n391), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(KEYINPUT9), .B(G234), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(G953), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n400), .A2(G217), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n390), .A2(new_n398), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n403), .B1(new_n390), .B2(new_n398), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n407), .A2(G902), .ZN(new_n408));
  INV_X1    g222(.A(G478), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n409), .A2(KEYINPUT15), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(KEYINPUT99), .A3(new_n410), .ZN(new_n411));
  OAI211_X1 g225(.A(KEYINPUT99), .B(new_n188), .C1(new_n405), .C2(new_n406), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n412), .B1(KEYINPUT15), .B2(new_n409), .ZN(new_n413));
  OR2_X1    g227(.A1(new_n405), .A2(new_n406), .ZN(new_n414));
  AOI21_X1  g228(.A(KEYINPUT99), .B1(new_n414), .B2(new_n188), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n411), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT100), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n416), .B(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(G234), .A2(G237), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n419), .A2(G952), .A3(new_n401), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT21), .B(G898), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(KEYINPUT101), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n419), .A2(G902), .A3(G953), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n420), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NOR3_X1   g239(.A1(new_n379), .A2(new_n418), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G221), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n427), .B1(new_n400), .B2(new_n188), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n312), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(G214), .B1(G237), .B2(G902), .ZN(new_n431));
  XOR2_X1   g245(.A(G116), .B(G119), .Z(new_n432));
  XNOR2_X1  g246(.A(KEYINPUT2), .B(G113), .ZN(new_n433));
  OR2_X1    g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n433), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(KEYINPUT68), .A3(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT68), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n432), .A2(new_n433), .A3(new_n437), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n272), .A2(new_n439), .A3(new_n284), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT86), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n272), .A2(new_n439), .A3(new_n284), .A4(KEYINPUT86), .ZN(new_n443));
  INV_X1    g257(.A(new_n223), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n444), .B1(new_n258), .B2(new_n259), .ZN(new_n445));
  INV_X1    g259(.A(new_n434), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n380), .A2(KEYINPUT5), .A3(G119), .ZN(new_n447));
  OR2_X1    g261(.A1(new_n447), .A2(KEYINPUT87), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(KEYINPUT87), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(G113), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G116), .B(G119), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT5), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n446), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n445), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(G110), .B(G122), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n442), .A2(new_n443), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT89), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n440), .A2(new_n441), .B1(new_n445), .B2(new_n454), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n460), .A2(KEYINPUT89), .A3(new_n443), .A4(new_n456), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT6), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n460), .A2(new_n443), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n456), .B(KEYINPUT88), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT90), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n244), .A2(new_n329), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n469), .B1(new_n329), .B2(new_n280), .ZN(new_n470));
  XOR2_X1   g284(.A(new_n470), .B(KEYINPUT91), .Z(new_n471));
  INV_X1    g285(.A(G224), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n472), .A2(G953), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n471), .B(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT90), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n462), .A2(new_n475), .A3(new_n466), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n464), .A2(new_n463), .A3(new_n465), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n468), .A2(new_n474), .A3(new_n476), .A4(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT7), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n470), .B(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n454), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n232), .A2(new_n482), .ZN(new_n483));
  OR2_X1    g297(.A1(new_n483), .A2(KEYINPUT94), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(KEYINPUT94), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n453), .B(KEYINPUT92), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n446), .B1(new_n486), .B2(new_n451), .ZN(new_n487));
  OR2_X1    g301(.A1(new_n487), .A2(KEYINPUT93), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(KEYINPUT93), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n488), .A2(new_n489), .A3(new_n445), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n484), .A2(new_n485), .A3(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n456), .B(KEYINPUT8), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n481), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT95), .ZN(new_n494));
  AOI22_X1  g308(.A1(new_n493), .A2(new_n494), .B1(new_n459), .B2(new_n461), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n491), .A2(new_n492), .ZN(new_n496));
  INV_X1    g310(.A(new_n481), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT95), .ZN(new_n499));
  AOI21_X1  g313(.A(G902), .B1(new_n495), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(G210), .B1(G237), .B2(G902), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n478), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n501), .B1(new_n478), .B2(new_n500), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n431), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n430), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT73), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n314), .A2(G210), .ZN(new_n507));
  XOR2_X1   g321(.A(new_n507), .B(KEYINPUT27), .Z(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT26), .B(G101), .ZN(new_n509));
  XOR2_X1   g323(.A(new_n508), .B(new_n509), .Z(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n248), .A2(new_n282), .A3(new_n286), .A4(new_n250), .ZN(new_n512));
  INV_X1    g326(.A(new_n439), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n193), .A2(new_n194), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n198), .A2(new_n199), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n189), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n207), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n517), .A2(new_n242), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n208), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n512), .A2(new_n513), .A3(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT71), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n519), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n280), .B1(new_n208), .B2(new_n203), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n439), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n512), .A2(KEYINPUT71), .A3(new_n513), .A4(new_n519), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n522), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n527), .A2(KEYINPUT28), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT28), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n520), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n506), .B(new_n511), .C1(new_n528), .C2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n512), .A2(KEYINPUT30), .A3(new_n519), .ZN(new_n533));
  AOI22_X1  g347(.A1(new_n285), .A2(new_n209), .B1(new_n518), .B2(new_n208), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT67), .B1(new_n534), .B2(KEYINPUT30), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT67), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT30), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n536), .B(new_n537), .C1(new_n523), .C2(new_n524), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n533), .A2(new_n439), .A3(new_n535), .A4(new_n538), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n539), .A2(new_n510), .A3(new_n522), .A4(new_n526), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT72), .B1(new_n540), .B2(KEYINPUT31), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(KEYINPUT31), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n540), .A2(KEYINPUT72), .A3(KEYINPUT31), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n531), .B1(new_n527), .B2(KEYINPUT28), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT73), .B1(new_n545), .B2(new_n510), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n532), .A2(new_n543), .A3(new_n544), .A4(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(G472), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(new_n548), .A3(new_n188), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT32), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT32), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n547), .A2(new_n551), .A3(new_n548), .A4(new_n188), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n539), .A2(new_n522), .A3(new_n526), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n555), .A2(new_n510), .ZN(new_n556));
  AOI211_X1 g370(.A(KEYINPUT29), .B(new_n556), .C1(new_n510), .C2(new_n545), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n512), .A2(new_n519), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n522), .B(new_n526), .C1(new_n513), .C2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n530), .B1(new_n560), .B2(new_n529), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n510), .A2(KEYINPUT29), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n188), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(G472), .B1(new_n557), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n553), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n333), .A2(new_n334), .ZN(new_n566));
  OR2_X1    g380(.A1(new_n240), .A2(G119), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n240), .A2(G119), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  XOR2_X1   g383(.A(KEYINPUT24), .B(G110), .Z(new_n570));
  INV_X1    g384(.A(KEYINPUT23), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n240), .A2(KEYINPUT23), .A3(G119), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n572), .A2(new_n567), .A3(new_n573), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n569), .A2(new_n570), .B1(new_n574), .B2(G110), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n566), .A2(new_n575), .ZN(new_n576));
  OAI22_X1  g390(.A1(new_n569), .A2(new_n570), .B1(new_n574), .B2(G110), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n333), .B(new_n577), .C1(new_n337), .C2(new_n339), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  XOR2_X1   g393(.A(KEYINPUT22), .B(G137), .Z(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(KEYINPUT76), .ZN(new_n581));
  INV_X1    g395(.A(G234), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n427), .A2(new_n582), .A3(G953), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n581), .B(new_n583), .ZN(new_n584));
  OR2_X1    g398(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n579), .A2(new_n584), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT77), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(KEYINPUT25), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n587), .A2(new_n188), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n585), .A2(new_n188), .A3(new_n586), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n591), .A2(new_n588), .A3(KEYINPUT25), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n593), .B1(new_n588), .B2(KEYINPUT25), .ZN(new_n594));
  OAI21_X1  g408(.A(G217), .B1(new_n582), .B2(G902), .ZN(new_n595));
  XOR2_X1   g409(.A(new_n595), .B(KEYINPUT74), .Z(new_n596));
  NAND2_X1  g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(G902), .B1(new_n582), .B2(G217), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n587), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n505), .A2(new_n565), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G101), .ZN(G3));
  INV_X1    g417(.A(new_n425), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n431), .B(new_n604), .C1(new_n502), .C2(new_n503), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n407), .A2(G478), .A3(G902), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT33), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n390), .A2(new_n398), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n607), .B1(new_n608), .B2(KEYINPUT102), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n407), .B(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n188), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n606), .B1(new_n612), .B2(G478), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n379), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n605), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n549), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n548), .B1(new_n547), .B2(new_n188), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n616), .A2(new_n617), .A3(new_n600), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n312), .A2(new_n429), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n615), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT34), .B(G104), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G6));
  NAND2_X1  g437(.A1(new_n362), .A2(new_n367), .ZN(new_n624));
  INV_X1    g438(.A(new_n372), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n370), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n418), .A2(new_n356), .A3(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n605), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n628), .A2(new_n618), .A3(new_n620), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT35), .B(G107), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G9));
  INV_X1    g445(.A(KEYINPUT103), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n616), .A2(new_n617), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT36), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n584), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n579), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n598), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n597), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n632), .B1(new_n633), .B2(new_n638), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n597), .A2(new_n637), .ZN(new_n640));
  NOR4_X1   g454(.A1(new_n616), .A2(new_n617), .A3(new_n640), .A4(KEYINPUT103), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n505), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT37), .B(G110), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G12));
  AOI21_X1  g458(.A(new_n619), .B1(new_n553), .B2(new_n564), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n418), .A2(new_n356), .ZN(new_n646));
  INV_X1    g460(.A(G900), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n420), .B1(new_n424), .B2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n646), .A2(KEYINPUT104), .A3(new_n626), .A4(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT104), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n651), .B1(new_n627), .B2(new_n648), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n650), .A2(new_n652), .A3(new_n638), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n504), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n645), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G128), .ZN(G30));
  XOR2_X1   g470(.A(new_n648), .B(KEYINPUT39), .Z(new_n657));
  NAND2_X1  g471(.A1(new_n620), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT40), .ZN(new_n659));
  INV_X1    g473(.A(new_n501), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n476), .A2(new_n477), .ZN(new_n661));
  INV_X1    g475(.A(new_n474), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n475), .B1(new_n462), .B2(new_n466), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n462), .B1(new_n498), .B2(KEYINPUT95), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n493), .A2(new_n494), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n188), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n660), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n478), .A2(new_n500), .A3(new_n501), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(KEYINPUT38), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT38), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n668), .A2(new_n672), .A3(new_n669), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n540), .B1(new_n560), .B2(new_n510), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n548), .B1(new_n675), .B2(new_n188), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n553), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n431), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n379), .A2(new_n418), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n638), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n674), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n659), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(new_n235), .ZN(G45));
  AOI21_X1  g498(.A(new_n375), .B1(new_n356), .B2(new_n374), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n377), .A2(new_n355), .A3(KEYINPUT98), .ZN(new_n686));
  OAI211_X1 g500(.A(new_n613), .B(new_n649), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n638), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n504), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n565), .A2(new_n690), .A3(new_n620), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G146), .ZN(G48));
  OR2_X1    g506(.A1(new_n294), .A2(new_n297), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n188), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(G469), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(new_n429), .A3(new_n298), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n615), .A2(new_n565), .A3(new_n601), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(KEYINPUT105), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT41), .B(G113), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G15));
  NAND4_X1  g515(.A1(new_n628), .A2(new_n565), .A3(new_n601), .A4(new_n697), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G116), .ZN(G18));
  NOR2_X1   g517(.A1(new_n504), .A2(new_n696), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n565), .A2(new_n704), .A3(new_n426), .A4(new_n638), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G119), .ZN(G21));
  NOR2_X1   g520(.A1(new_n504), .A2(new_n680), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n561), .A2(new_n511), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT31), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n540), .B(new_n709), .ZN(new_n710));
  AOI211_X1 g524(.A(G472), .B(G902), .C1(new_n708), .C2(new_n710), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n617), .A2(new_n711), .A3(new_n600), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n707), .A2(new_n604), .A3(new_n697), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT106), .B(G122), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G24));
  NAND2_X1  g529(.A1(new_n687), .A2(KEYINPUT107), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT107), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n379), .A2(new_n717), .A3(new_n613), .A4(new_n649), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NOR4_X1   g533(.A1(new_n719), .A2(new_n617), .A3(new_n640), .A4(new_n711), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n704), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G125), .ZN(G27));
  XOR2_X1   g536(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n723));
  OAI21_X1  g537(.A(new_n298), .B1(new_n310), .B2(new_n187), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n724), .A2(KEYINPUT108), .A3(new_n429), .ZN(new_n725));
  AOI21_X1  g539(.A(KEYINPUT108), .B1(new_n724), .B2(new_n429), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n668), .A2(new_n431), .A3(new_n669), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n565), .A2(new_n729), .A3(new_n601), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n723), .B1(new_n730), .B2(new_n719), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT110), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n553), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n550), .A2(KEYINPUT110), .A3(new_n552), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n564), .A3(new_n734), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n716), .A2(KEYINPUT42), .A3(new_n718), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n735), .A2(new_n601), .A3(new_n729), .A4(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n731), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G131), .ZN(G33));
  AND2_X1   g553(.A1(new_n650), .A2(new_n652), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n565), .A2(new_n729), .A3(new_n601), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G134), .ZN(G36));
  AND3_X1   g556(.A1(new_n613), .A2(new_n376), .A3(new_n378), .ZN(new_n743));
  XOR2_X1   g557(.A(KEYINPUT111), .B(KEYINPUT43), .Z(new_n744));
  OR2_X1    g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT43), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n743), .A2(KEYINPUT111), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(KEYINPUT112), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n745), .A2(new_n750), .A3(new_n747), .ZN(new_n751));
  AOI211_X1 g565(.A(new_n640), .B(new_n633), .C1(new_n749), .C2(new_n751), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n752), .A2(KEYINPUT44), .ZN(new_n753));
  INV_X1    g567(.A(new_n728), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n307), .B(KEYINPUT45), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(G469), .ZN(new_n756));
  NAND2_X1  g570(.A1(G469), .A2(G902), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(KEYINPUT46), .A3(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT46), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n759), .B(G469), .C1(new_n755), .C2(G902), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n758), .A2(new_n298), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n429), .A3(new_n657), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n752), .A2(KEYINPUT44), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n753), .A2(new_n754), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(KEYINPUT113), .B(G137), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n765), .B(new_n766), .ZN(G39));
  NAND2_X1  g581(.A1(new_n761), .A2(new_n429), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT47), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n761), .A2(KEYINPUT47), .A3(new_n429), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR4_X1   g586(.A1(new_n565), .A2(new_n601), .A3(new_n687), .A4(new_n728), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G140), .ZN(G42));
  NAND2_X1  g589(.A1(new_n695), .A2(new_n298), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(KEYINPUT49), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n601), .A2(new_n431), .A3(new_n429), .A4(new_n743), .ZN(new_n778));
  OR4_X1    g592(.A1(new_n674), .A2(new_n678), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n720), .A2(new_n729), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n416), .A2(new_n649), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n638), .A2(new_n356), .A3(new_n626), .A4(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n728), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n565), .A2(new_n620), .A3(new_n784), .ZN(new_n785));
  AND4_X1   g599(.A1(new_n780), .A2(new_n741), .A3(new_n781), .A4(new_n785), .ZN(new_n786));
  AOI22_X1  g600(.A1(new_n645), .A2(new_n784), .B1(new_n720), .B2(new_n729), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n780), .B1(new_n787), .B2(new_n741), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n698), .A2(new_n702), .A3(new_n713), .A4(new_n705), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n786), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n605), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n614), .B1(new_n379), .B2(new_n416), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n791), .A2(new_n618), .A3(new_n620), .A4(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n642), .A2(new_n602), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n794), .B1(new_n731), .B2(new_n737), .ZN(new_n795));
  AND4_X1   g609(.A1(new_n429), .A2(new_n640), .A3(new_n649), .A4(new_n724), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n678), .A2(new_n707), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n655), .A2(new_n691), .A3(new_n797), .A4(new_n721), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n801));
  AOI22_X1  g615(.A1(new_n645), .A2(new_n654), .B1(new_n720), .B2(new_n704), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n802), .A2(KEYINPUT52), .A3(new_n691), .A4(new_n797), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n800), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  OR3_X1    g618(.A1(new_n798), .A2(new_n801), .A3(new_n799), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n790), .A2(new_n795), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n800), .A2(new_n803), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n786), .A2(new_n788), .ZN(new_n810));
  AND4_X1   g624(.A1(new_n698), .A2(new_n702), .A3(new_n705), .A4(new_n713), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n809), .A2(new_n810), .A3(new_n795), .A4(new_n811), .ZN(new_n812));
  XOR2_X1   g626(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n813));
  OAI21_X1  g627(.A(new_n808), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT54), .ZN(new_n815));
  INV_X1    g629(.A(new_n420), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n678), .A2(new_n600), .A3(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n754), .A2(KEYINPUT117), .A3(new_n697), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n819), .B1(new_n728), .B2(new_n696), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n817), .A2(new_n821), .A3(new_n379), .A4(new_n613), .ZN(new_n822));
  INV_X1    g636(.A(G952), .ZN(new_n823));
  INV_X1    g637(.A(new_n712), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n745), .A2(new_n420), .A3(new_n747), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI211_X1 g640(.A(new_n823), .B(G953), .C1(new_n826), .C2(new_n704), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n735), .A2(new_n601), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n825), .B1(new_n818), .B2(new_n820), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n830), .A2(KEYINPUT119), .ZN(new_n831));
  OAI21_X1  g645(.A(KEYINPUT48), .B1(new_n830), .B2(KEYINPUT119), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n822), .B(new_n827), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT118), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n770), .B(new_n771), .C1(new_n429), .C2(new_n776), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n824), .A2(new_n728), .A3(new_n825), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(KEYINPUT51), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n838), .A2(new_n839), .ZN(new_n842));
  INV_X1    g656(.A(new_n674), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n696), .A2(new_n431), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n843), .A2(new_n826), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT50), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n843), .A2(new_n826), .A3(KEYINPUT50), .A4(new_n844), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n617), .A2(new_n640), .A3(new_n711), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n829), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n379), .A2(new_n613), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n817), .A2(new_n821), .A3(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n842), .A2(new_n849), .A3(new_n851), .A4(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n841), .B(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT120), .B1(new_n836), .B2(new_n855), .ZN(new_n856));
  XOR2_X1   g670(.A(new_n841), .B(new_n854), .Z(new_n857));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n857), .A2(new_n858), .A3(new_n835), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n741), .A2(new_n781), .A3(new_n785), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT114), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n787), .A2(new_n780), .A3(new_n741), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n811), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n794), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n738), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n866), .A2(KEYINPUT53), .A3(new_n805), .A4(new_n804), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n812), .A2(new_n813), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  AND4_X1   g684(.A1(new_n815), .A2(new_n856), .A3(new_n859), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n823), .A2(new_n401), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(KEYINPUT121), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n779), .B1(new_n871), .B2(new_n873), .ZN(G75));
  NOR2_X1   g688(.A1(new_n806), .A2(new_n807), .ZN(new_n875));
  INV_X1    g689(.A(new_n813), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n876), .B1(new_n866), .B2(new_n809), .ZN(new_n877));
  OAI211_X1 g691(.A(G210), .B(G902), .C1(new_n875), .C2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT56), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT122), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n662), .B1(new_n661), .B2(new_n663), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n478), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT55), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n878), .A2(KEYINPUT122), .A3(new_n879), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n880), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT122), .ZN(new_n886));
  INV_X1    g700(.A(G210), .ZN(new_n887));
  AOI211_X1 g701(.A(new_n887), .B(new_n188), .C1(new_n867), .C2(new_n868), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n886), .B(new_n883), .C1(new_n888), .C2(KEYINPUT56), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n823), .A2(G953), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT123), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n885), .A2(new_n892), .ZN(G51));
  INV_X1    g707(.A(new_n891), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n757), .B(KEYINPUT57), .Z(new_n895));
  INV_X1    g709(.A(new_n870), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n869), .B1(new_n867), .B2(new_n868), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n693), .ZN(new_n899));
  OAI21_X1  g713(.A(G902), .B1(new_n875), .B2(new_n877), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n900), .A2(new_n756), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n894), .B1(new_n899), .B2(new_n901), .ZN(G54));
  NAND2_X1  g716(.A1(KEYINPUT58), .A2(G475), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n904), .A2(new_n624), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n624), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n894), .B1(new_n905), .B2(new_n906), .ZN(G60));
  NAND2_X1  g721(.A1(new_n815), .A2(new_n870), .ZN(new_n908));
  NAND2_X1  g722(.A1(G478), .A2(G902), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT59), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n611), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n611), .B(new_n910), .C1(new_n896), .C2(new_n897), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n891), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n911), .A2(new_n913), .ZN(G63));
  NAND2_X1  g728(.A1(G217), .A2(G902), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT60), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(new_n867), .B2(new_n868), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n917), .A2(new_n587), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n894), .B1(new_n917), .B2(new_n636), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT124), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n917), .B2(new_n636), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n922), .A2(KEYINPUT61), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n918), .B(new_n919), .C1(new_n922), .C2(KEYINPUT61), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(G66));
  OAI21_X1  g740(.A(G953), .B1(new_n423), .B2(new_n472), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n789), .A2(new_n794), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n927), .B1(new_n928), .B2(G953), .ZN(new_n929));
  OAI22_X1  g743(.A1(new_n661), .A2(new_n663), .B1(G898), .B2(new_n401), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(G69));
  INV_X1    g745(.A(new_n658), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n754), .A2(new_n792), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n932), .A2(new_n933), .A3(new_n565), .A4(new_n601), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n765), .A2(new_n774), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n802), .A2(new_n691), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n683), .A2(new_n936), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n937), .A2(KEYINPUT62), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n937), .A2(KEYINPUT62), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(KEYINPUT125), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT125), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n935), .B(new_n942), .C1(new_n939), .C2(new_n938), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n533), .A2(new_n535), .A3(new_n538), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(new_n359), .Z(new_n946));
  NAND3_X1  g760(.A1(new_n944), .A2(new_n401), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n647), .B1(new_n946), .B2(new_n290), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n753), .A2(new_n754), .A3(new_n764), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n828), .A2(new_n707), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n762), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n951), .A2(G953), .ZN(new_n952));
  INV_X1    g766(.A(new_n738), .ZN(new_n953));
  INV_X1    g767(.A(new_n774), .ZN(new_n954));
  INV_X1    g768(.A(new_n741), .ZN(new_n955));
  NOR4_X1   g769(.A1(new_n953), .A2(new_n954), .A3(new_n955), .A4(new_n936), .ZN(new_n956));
  AOI22_X1  g770(.A1(new_n952), .A2(new_n956), .B1(G227), .B2(G953), .ZN(new_n957));
  OAI221_X1 g771(.A(new_n947), .B1(new_n401), .B2(new_n948), .C1(new_n946), .C2(new_n957), .ZN(G72));
  NAND2_X1  g772(.A1(new_n554), .A2(new_n510), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n941), .A2(new_n928), .A3(new_n943), .ZN(new_n960));
  XNOR2_X1  g774(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n548), .A2(new_n188), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT127), .Z(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n959), .B1(new_n960), .B2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n540), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n556), .A2(new_n967), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n814), .A2(new_n963), .A3(new_n968), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n951), .A2(new_n794), .A3(new_n789), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n964), .B1(new_n970), .B2(new_n956), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n555), .A2(new_n511), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n891), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NOR3_X1   g787(.A1(new_n966), .A2(new_n969), .A3(new_n973), .ZN(G57));
endmodule


