

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786;

  NOR2_X1 U381 ( .A1(n632), .A2(n611), .ZN(n730) );
  NOR2_X1 U382 ( .A1(n591), .A2(n365), .ZN(n364) );
  NAND2_X1 U383 ( .A1(n727), .A2(n714), .ZN(n658) );
  NAND2_X1 U384 ( .A1(n699), .A2(n652), .ZN(n653) );
  INV_X1 U385 ( .A(KEYINPUT31), .ZN(n368) );
  INV_X1 U386 ( .A(KEYINPUT78), .ZN(n370) );
  NAND2_X1 U387 ( .A1(n600), .A2(n677), .ZN(n680) );
  AND2_X1 U388 ( .A1(n690), .A2(n478), .ZN(n606) );
  XNOR2_X1 U389 ( .A(n767), .B(n490), .ZN(n523) );
  XOR2_X1 U390 ( .A(G146), .B(G125), .Z(n557) );
  XNOR2_X2 U391 ( .A(n362), .B(KEYINPUT22), .ZN(n635) );
  NAND2_X2 U392 ( .A1(n440), .A2(n467), .ZN(n362) );
  NAND2_X1 U393 ( .A1(n363), .A2(n577), .ZN(n602) );
  XNOR2_X1 U394 ( .A(n576), .B(KEYINPUT28), .ZN(n363) );
  NAND2_X1 U395 ( .A1(n366), .A2(n364), .ZN(n594) );
  INV_X1 U396 ( .A(n593), .ZN(n365) );
  INV_X1 U397 ( .A(n590), .ZN(n366) );
  NAND2_X1 U398 ( .A1(n367), .A2(n388), .ZN(n480) );
  NAND2_X1 U399 ( .A1(n623), .A2(n482), .ZN(n367) );
  XOR2_X2 U400 ( .A(n737), .B(n736), .Z(n390) );
  XNOR2_X2 U401 ( .A(n748), .B(n747), .ZN(n391) );
  NOR2_X2 U402 ( .A1(n680), .A2(n679), .ZN(n601) );
  OR2_X2 U403 ( .A1(n456), .A2(n708), .ZN(n453) );
  XNOR2_X2 U404 ( .A(n450), .B(KEYINPUT35), .ZN(n778) );
  OR2_X2 U405 ( .A1(n661), .A2(n712), .ZN(n375) );
  XNOR2_X2 U406 ( .A(n653), .B(n368), .ZN(n727) );
  AND2_X2 U407 ( .A1(n395), .A2(n630), .ZN(n440) );
  NAND2_X1 U408 ( .A1(n785), .A2(n780), .ZN(n639) );
  XNOR2_X1 U409 ( .A(n462), .B(KEYINPUT106), .ZN(n785) );
  AND2_X2 U410 ( .A1(n673), .A2(n622), .ZN(n482) );
  XNOR2_X1 U411 ( .A(n637), .B(KEYINPUT32), .ZN(n780) );
  OR2_X2 U412 ( .A1(n742), .A2(G902), .ZN(n461) );
  NOR2_X1 U413 ( .A1(n635), .A2(n369), .ZN(n636) );
  XNOR2_X2 U414 ( .A(n633), .B(n370), .ZN(n369) );
  XNOR2_X1 U415 ( .A(G110), .B(G128), .ZN(n517) );
  XOR2_X1 U416 ( .A(n693), .B(KEYINPUT6), .Z(n645) );
  OR2_X2 U417 ( .A1(n422), .A2(n378), .ZN(n395) );
  NOR2_X1 U418 ( .A1(n709), .A2(n602), .ZN(n603) );
  NAND2_X1 U419 ( .A1(n415), .A2(n382), .ZN(n693) );
  NOR2_X1 U420 ( .A1(G953), .A2(G237), .ZN(n549) );
  XNOR2_X1 U421 ( .A(n375), .B(n374), .ZN(n373) );
  NOR2_X1 U422 ( .A1(n645), .A2(n651), .ZN(n444) );
  OR2_X1 U423 ( .A1(n670), .A2(n412), .ZN(n411) );
  INV_X1 U424 ( .A(KEYINPUT86), .ZN(n374) );
  NAND2_X1 U425 ( .A1(n402), .A2(n476), .ZN(n662) );
  NAND2_X1 U426 ( .A1(n376), .A2(n373), .ZN(n372) );
  NOR2_X1 U427 ( .A1(n781), .A2(n783), .ZN(n433) );
  NAND2_X1 U428 ( .A1(n453), .A2(n451), .ZN(n450) );
  OR2_X1 U429 ( .A1(n655), .A2(KEYINPUT34), .ZN(n456) );
  NAND2_X1 U430 ( .A1(n395), .A2(n466), .ZN(n655) );
  AND2_X1 U431 ( .A1(n471), .A2(n384), .ZN(n466) );
  XNOR2_X1 U432 ( .A(n444), .B(n385), .ZN(n708) );
  BUF_X1 U433 ( .A(n579), .Z(n618) );
  INV_X1 U434 ( .A(n752), .ZN(n447) );
  XNOR2_X1 U435 ( .A(n523), .B(n524), .ZN(n565) );
  BUF_X1 U436 ( .A(n667), .Z(n439) );
  XNOR2_X1 U437 ( .A(n557), .B(n558), .ZN(n559) );
  XNOR2_X1 U438 ( .A(n455), .B(G953), .ZN(n667) );
  XNOR2_X1 U439 ( .A(G119), .B(KEYINPUT24), .ZN(n513) );
  NAND2_X1 U440 ( .A1(n371), .A2(n644), .ZN(n376) );
  XNOR2_X1 U441 ( .A(n639), .B(n638), .ZN(n371) );
  XNOR2_X2 U442 ( .A(n372), .B(KEYINPUT45), .ZN(n673) );
  XNOR2_X2 U443 ( .A(n618), .B(n595), .ZN(n600) );
  NOR2_X1 U444 ( .A1(n734), .A2(n477), .ZN(n476) );
  INV_X1 U445 ( .A(n732), .ZN(n477) );
  XNOR2_X1 U446 ( .A(n485), .B(KEYINPUT92), .ZN(n621) );
  XNOR2_X1 U447 ( .A(G902), .B(KEYINPUT15), .ZN(n485) );
  OR2_X1 U448 ( .A1(G902), .A2(G237), .ZN(n567) );
  XNOR2_X1 U449 ( .A(n408), .B(G119), .ZN(n562) );
  INV_X1 U450 ( .A(KEYINPUT3), .ZN(n408) );
  INV_X1 U451 ( .A(G122), .ZN(n398) );
  XNOR2_X1 U452 ( .A(n526), .B(G116), .ZN(n563) );
  XOR2_X1 U453 ( .A(KEYINPUT103), .B(G140), .Z(n543) );
  XNOR2_X1 U454 ( .A(G143), .B(G131), .ZN(n542) );
  XNOR2_X1 U455 ( .A(KEYINPUT12), .B(KEYINPUT102), .ZN(n544) );
  XOR2_X1 U456 ( .A(KEYINPUT101), .B(KEYINPUT11), .Z(n545) );
  XNOR2_X1 U457 ( .A(KEYINPUT68), .B(G101), .ZN(n490) );
  XNOR2_X1 U458 ( .A(G131), .B(G134), .ZN(n768) );
  INV_X1 U459 ( .A(KEYINPUT64), .ZN(n455) );
  NOR2_X1 U460 ( .A1(n469), .A2(n691), .ZN(n468) );
  XNOR2_X1 U461 ( .A(n532), .B(n460), .ZN(n459) );
  INV_X1 U462 ( .A(G469), .ZN(n460) );
  NAND2_X1 U463 ( .A1(n417), .A2(G902), .ZN(n414) );
  NAND2_X1 U464 ( .A1(n492), .A2(n413), .ZN(n412) );
  INV_X1 U465 ( .A(G902), .ZN(n413) );
  NAND2_X1 U466 ( .A1(n439), .A2(G227), .ZN(n457) );
  XNOR2_X1 U467 ( .A(n525), .B(n526), .ZN(n458) );
  XOR2_X1 U468 ( .A(G104), .B(KEYINPUT76), .Z(n525) );
  XOR2_X1 U469 ( .A(G137), .B(G140), .Z(n527) );
  INV_X1 U470 ( .A(KEYINPUT43), .ZN(n426) );
  XNOR2_X1 U471 ( .A(n420), .B(n597), .ZN(n619) );
  NOR2_X1 U472 ( .A1(n596), .A2(n676), .ZN(n420) );
  NAND2_X1 U473 ( .A1(n443), .A2(n642), .ZN(n452) );
  NAND2_X1 U474 ( .A1(n708), .A2(KEYINPUT34), .ZN(n443) );
  XNOR2_X1 U475 ( .A(n554), .B(n431), .ZN(n599) );
  XNOR2_X1 U476 ( .A(n555), .B(n432), .ZN(n431) );
  INV_X1 U477 ( .A(G475), .ZN(n432) );
  INV_X1 U478 ( .A(n693), .ZN(n575) );
  NAND2_X1 U479 ( .A1(n397), .A2(G475), .ZN(n449) );
  XNOR2_X1 U480 ( .A(n474), .B(KEYINPUT119), .ZN(n473) );
  NAND2_X1 U481 ( .A1(n475), .A2(n711), .ZN(n474) );
  INV_X1 U482 ( .A(n681), .ZN(n657) );
  XNOR2_X1 U483 ( .A(KEYINPUT98), .B(KEYINPUT20), .ZN(n501) );
  XNOR2_X1 U484 ( .A(n594), .B(n430), .ZN(n429) );
  NOR2_X1 U485 ( .A1(n612), .A2(n730), .ZN(n613) );
  INV_X1 U486 ( .A(KEYINPUT74), .ZN(n430) );
  NAND2_X1 U487 ( .A1(G234), .A2(G237), .ZN(n494) );
  NOR2_X1 U488 ( .A1(n722), .A2(n718), .ZN(n681) );
  XNOR2_X1 U489 ( .A(n406), .B(G116), .ZN(n405) );
  AND2_X1 U490 ( .A1(n549), .A2(G210), .ZN(n406) );
  XOR2_X1 U491 ( .A(G113), .B(KEYINPUT5), .Z(n488) );
  XNOR2_X1 U492 ( .A(n674), .B(KEYINPUT75), .ZN(n623) );
  XOR2_X1 U493 ( .A(KEYINPUT93), .B(KEYINPUT77), .Z(n558) );
  XOR2_X1 U494 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n556) );
  NOR2_X1 U495 ( .A1(n691), .A2(n381), .ZN(n478) );
  NOR2_X1 U496 ( .A1(n416), .A2(n410), .ZN(n409) );
  INV_X1 U497 ( .A(n677), .ZN(n416) );
  INV_X1 U498 ( .A(KEYINPUT0), .ZN(n470) );
  XNOR2_X1 U499 ( .A(n563), .B(KEYINPUT16), .ZN(n423) );
  INV_X1 U500 ( .A(KEYINPUT8), .ZN(n441) );
  XOR2_X1 U501 ( .A(G122), .B(G134), .Z(n539) );
  XNOR2_X1 U502 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U503 ( .A(n424), .B(G478), .ZN(n598) );
  NOR2_X1 U504 ( .A1(n664), .A2(G902), .ZN(n424) );
  XNOR2_X1 U505 ( .A(n565), .B(n531), .ZN(n742) );
  XNOR2_X1 U506 ( .A(n458), .B(n457), .ZN(n530) );
  XNOR2_X1 U507 ( .A(n616), .B(n425), .ZN(n617) );
  XNOR2_X1 U508 ( .A(n426), .B(KEYINPUT109), .ZN(n425) );
  XNOR2_X1 U509 ( .A(n419), .B(n418), .ZN(n783) );
  INV_X1 U510 ( .A(KEYINPUT40), .ZN(n418) );
  NOR2_X1 U511 ( .A1(n383), .A2(n452), .ZN(n451) );
  NOR2_X1 U512 ( .A1(n572), .A2(n599), .ZN(n722) );
  NOR2_X1 U513 ( .A1(n598), .A2(n573), .ZN(n718) );
  INV_X1 U514 ( .A(KEYINPUT60), .ZN(n445) );
  NAND2_X1 U515 ( .A1(n448), .A2(n447), .ZN(n446) );
  XNOR2_X1 U516 ( .A(n449), .B(n391), .ZN(n448) );
  INV_X1 U517 ( .A(G953), .ZN(n472) );
  OR2_X2 U518 ( .A1(n663), .A2(n662), .ZN(n377) );
  OR2_X1 U519 ( .A1(n628), .A2(KEYINPUT0), .ZN(n378) );
  OR2_X1 U520 ( .A1(KEYINPUT2), .A2(n675), .ZN(n379) );
  AND2_X1 U521 ( .A1(n411), .A2(n409), .ZN(n380) );
  AND2_X1 U522 ( .A1(n499), .A2(n624), .ZN(n381) );
  AND2_X1 U523 ( .A1(n411), .A2(n414), .ZN(n382) );
  AND2_X1 U524 ( .A1(n655), .A2(KEYINPUT34), .ZN(n383) );
  OR2_X1 U525 ( .A1(n629), .A2(n470), .ZN(n384) );
  INV_X1 U526 ( .A(G107), .ZN(n526) );
  XOR2_X1 U527 ( .A(n640), .B(KEYINPUT33), .Z(n385) );
  NOR2_X1 U528 ( .A1(n709), .A2(n708), .ZN(n386) );
  XOR2_X1 U529 ( .A(KEYINPUT48), .B(KEYINPUT70), .Z(n387) );
  XOR2_X1 U530 ( .A(n487), .B(KEYINPUT67), .Z(n388) );
  XOR2_X1 U531 ( .A(n670), .B(KEYINPUT62), .Z(n389) );
  XOR2_X1 U532 ( .A(n672), .B(KEYINPUT112), .Z(n392) );
  XOR2_X1 U533 ( .A(KEYINPUT84), .B(KEYINPUT56), .Z(n393) );
  XOR2_X1 U534 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n394) );
  XNOR2_X1 U535 ( .A(n401), .B(n562), .ZN(n400) );
  BUF_X1 U536 ( .A(n759), .Z(n396) );
  XNOR2_X1 U537 ( .A(n400), .B(n423), .ZN(n759) );
  AND2_X2 U538 ( .A1(n480), .A2(n377), .ZN(n397) );
  AND2_X1 U539 ( .A1(n480), .A2(n377), .ZN(n421) );
  INV_X1 U540 ( .A(n401), .ZN(n561) );
  XNOR2_X2 U541 ( .A(n399), .B(n398), .ZN(n401) );
  XNOR2_X2 U542 ( .A(G104), .B(G113), .ZN(n399) );
  XNOR2_X2 U543 ( .A(n662), .B(n620), .ZN(n674) );
  XNOR2_X1 U544 ( .A(n403), .B(n387), .ZN(n402) );
  NAND2_X1 U545 ( .A1(n613), .A2(n429), .ZN(n403) );
  XNOR2_X1 U546 ( .A(n489), .B(n404), .ZN(n491) );
  XNOR2_X1 U547 ( .A(n407), .B(n405), .ZN(n404) );
  XNOR2_X1 U548 ( .A(n488), .B(n562), .ZN(n407) );
  NAND2_X1 U549 ( .A1(n415), .A2(n380), .ZN(n493) );
  INV_X1 U550 ( .A(n414), .ZN(n410) );
  NAND2_X1 U551 ( .A1(n670), .A2(n417), .ZN(n415) );
  INV_X1 U552 ( .A(n492), .ZN(n417) );
  NAND2_X1 U553 ( .A1(n619), .A2(n722), .ZN(n419) );
  NAND2_X1 U554 ( .A1(n421), .A2(G478), .ZN(n666) );
  NAND2_X1 U555 ( .A1(n421), .A2(G472), .ZN(n671) );
  NAND2_X1 U556 ( .A1(n397), .A2(G210), .ZN(n738) );
  NAND2_X1 U557 ( .A1(n397), .A2(G217), .ZN(n749) );
  NAND2_X1 U558 ( .A1(n397), .A2(G469), .ZN(n743) );
  NAND2_X1 U559 ( .A1(n422), .A2(KEYINPUT0), .ZN(n471) );
  NOR2_X1 U560 ( .A1(n602), .A2(n422), .ZN(n587) );
  XNOR2_X2 U561 ( .A(n608), .B(n581), .ZN(n422) );
  XNOR2_X2 U562 ( .A(n603), .B(KEYINPUT42), .ZN(n781) );
  NOR2_X1 U563 ( .A1(n647), .A2(n575), .ZN(n463) );
  XNOR2_X1 U564 ( .A(n552), .B(n553), .ZN(n746) );
  NAND2_X1 U565 ( .A1(n428), .A2(KEYINPUT80), .ZN(n588) );
  NAND2_X1 U566 ( .A1(n657), .A2(n587), .ZN(n428) );
  XNOR2_X1 U567 ( .A(n446), .B(n445), .ZN(G60) );
  XNOR2_X1 U568 ( .A(n433), .B(n604), .ZN(n612) );
  XNOR2_X1 U569 ( .A(n434), .B(n393), .ZN(G51) );
  NAND2_X1 U570 ( .A1(n438), .A2(n447), .ZN(n434) );
  XNOR2_X1 U571 ( .A(n435), .B(n392), .ZN(G57) );
  NAND2_X1 U572 ( .A1(n437), .A2(n447), .ZN(n435) );
  NOR2_X2 U573 ( .A1(n635), .A2(n686), .ZN(n646) );
  NAND2_X1 U574 ( .A1(n377), .A2(n379), .ZN(n475) );
  XNOR2_X1 U575 ( .A(n436), .B(n394), .ZN(G75) );
  NAND2_X1 U576 ( .A1(n473), .A2(n472), .ZN(n436) );
  XNOR2_X1 U577 ( .A(n671), .B(n389), .ZN(n437) );
  XNOR2_X1 U578 ( .A(n738), .B(n390), .ZN(n438) );
  NOR2_X2 U579 ( .A1(n691), .A2(n690), .ZN(n687) );
  XNOR2_X1 U580 ( .A(n442), .B(n441), .ZN(n537) );
  NAND2_X1 U581 ( .A1(n667), .A2(G234), .ZN(n442) );
  NOR2_X1 U582 ( .A1(n750), .A2(G902), .ZN(n479) );
  XNOR2_X2 U583 ( .A(n534), .B(KEYINPUT4), .ZN(n767) );
  XNOR2_X1 U584 ( .A(n454), .B(n556), .ZN(n560) );
  NAND2_X1 U585 ( .A1(n667), .A2(G224), .ZN(n454) );
  XNOR2_X2 U586 ( .A(n605), .B(KEYINPUT1), .ZN(n686) );
  XNOR2_X2 U587 ( .A(n461), .B(n459), .ZN(n605) );
  NAND2_X1 U588 ( .A1(n464), .A2(n463), .ZN(n462) );
  XNOR2_X1 U589 ( .A(n646), .B(n465), .ZN(n464) );
  INV_X1 U590 ( .A(KEYINPUT105), .ZN(n465) );
  AND2_X1 U591 ( .A1(n471), .A2(n468), .ZN(n467) );
  INV_X1 U592 ( .A(n384), .ZN(n469) );
  XNOR2_X2 U593 ( .A(n479), .B(n522), .ZN(n690) );
  XNOR2_X2 U594 ( .A(n580), .B(KEYINPUT88), .ZN(n608) );
  XNOR2_X1 U595 ( .A(n759), .B(n564), .ZN(n566) );
  XNOR2_X1 U596 ( .A(n560), .B(n559), .ZN(n564) );
  XOR2_X2 U597 ( .A(G143), .B(G128), .Z(n534) );
  NOR2_X1 U598 ( .A1(n439), .A2(G952), .ZN(n752) );
  NOR2_X1 U599 ( .A1(n500), .A2(n381), .ZN(n483) );
  AND2_X1 U600 ( .A1(n549), .A2(G214), .ZN(n484) );
  INV_X1 U601 ( .A(n621), .ZN(n622) );
  INV_X1 U602 ( .A(KEYINPUT83), .ZN(n620) );
  AND2_X1 U603 ( .A1(n606), .A2(n575), .ZN(n576) );
  INV_X1 U604 ( .A(n654), .ZN(n533) );
  INV_X1 U605 ( .A(KEYINPUT39), .ZN(n597) );
  XNOR2_X1 U606 ( .A(KEYINPUT82), .B(n622), .ZN(n486) );
  NAND2_X1 U607 ( .A1(n486), .A2(KEYINPUT2), .ZN(n487) );
  XNOR2_X1 U608 ( .A(G146), .B(n768), .ZN(n528) );
  XNOR2_X1 U609 ( .A(n528), .B(G137), .ZN(n489) );
  XNOR2_X1 U610 ( .A(n491), .B(n523), .ZN(n670) );
  XNOR2_X1 U611 ( .A(KEYINPUT100), .B(G472), .ZN(n492) );
  NAND2_X1 U612 ( .A1(G214), .A2(n567), .ZN(n677) );
  XNOR2_X1 U613 ( .A(n493), .B(KEYINPUT30), .ZN(n500) );
  XNOR2_X1 U614 ( .A(n494), .B(KEYINPUT14), .ZN(n497) );
  NAND2_X1 U615 ( .A1(G902), .A2(n497), .ZN(n625) );
  NOR2_X1 U616 ( .A1(G900), .A2(n625), .ZN(n495) );
  INV_X1 U617 ( .A(n439), .ZN(n771) );
  NAND2_X1 U618 ( .A1(n495), .A2(n771), .ZN(n496) );
  XNOR2_X1 U619 ( .A(KEYINPUT108), .B(n496), .ZN(n499) );
  NAND2_X1 U620 ( .A1(n497), .A2(G952), .ZN(n707) );
  NOR2_X1 U621 ( .A1(G953), .A2(n707), .ZN(n498) );
  XOR2_X1 U622 ( .A(KEYINPUT94), .B(n498), .Z(n624) );
  NAND2_X1 U623 ( .A1(G234), .A2(n621), .ZN(n502) );
  XNOR2_X1 U624 ( .A(n502), .B(n501), .ZN(n504) );
  NAND2_X1 U625 ( .A1(G221), .A2(n504), .ZN(n503) );
  XNOR2_X1 U626 ( .A(KEYINPUT21), .B(n503), .ZN(n691) );
  NAND2_X1 U627 ( .A1(G217), .A2(n504), .ZN(n505) );
  XOR2_X1 U628 ( .A(n505), .B(KEYINPUT99), .Z(n507) );
  XNOR2_X1 U629 ( .A(KEYINPUT25), .B(KEYINPUT97), .ZN(n506) );
  XNOR2_X1 U630 ( .A(n507), .B(n506), .ZN(n522) );
  XOR2_X1 U631 ( .A(KEYINPUT10), .B(KEYINPUT69), .Z(n508) );
  XNOR2_X1 U632 ( .A(n557), .B(n508), .ZN(n548) );
  XNOR2_X1 U633 ( .A(n527), .B(n548), .ZN(n766) );
  INV_X1 U634 ( .A(KEYINPUT23), .ZN(n509) );
  NAND2_X1 U635 ( .A1(KEYINPUT96), .A2(n509), .ZN(n512) );
  INV_X1 U636 ( .A(KEYINPUT96), .ZN(n510) );
  NAND2_X1 U637 ( .A1(n510), .A2(KEYINPUT23), .ZN(n511) );
  NAND2_X1 U638 ( .A1(n512), .A2(n511), .ZN(n514) );
  XNOR2_X1 U639 ( .A(n514), .B(n513), .ZN(n516) );
  INV_X1 U640 ( .A(KEYINPUT81), .ZN(n515) );
  XNOR2_X1 U641 ( .A(n516), .B(n515), .ZN(n518) );
  XNOR2_X1 U642 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U643 ( .A(n766), .B(n519), .ZN(n521) );
  AND2_X1 U644 ( .A1(G221), .A2(n537), .ZN(n520) );
  XNOR2_X1 U645 ( .A(n521), .B(n520), .ZN(n750) );
  XNOR2_X1 U646 ( .A(G110), .B(KEYINPUT73), .ZN(n524) );
  XNOR2_X1 U647 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U648 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U649 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n532) );
  NAND2_X1 U650 ( .A1(n687), .A2(n605), .ZN(n654) );
  NAND2_X1 U651 ( .A1(n483), .A2(n533), .ZN(n596) );
  XOR2_X1 U652 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n536) );
  XNOR2_X1 U653 ( .A(n534), .B(n563), .ZN(n535) );
  XNOR2_X1 U654 ( .A(n536), .B(n535), .ZN(n541) );
  NAND2_X1 U655 ( .A1(G217), .A2(n537), .ZN(n538) );
  XNOR2_X1 U656 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U657 ( .A(n541), .B(n540), .ZN(n664) );
  INV_X1 U658 ( .A(n598), .ZN(n572) );
  XNOR2_X1 U659 ( .A(KEYINPUT13), .B(KEYINPUT104), .ZN(n555) );
  XNOR2_X1 U660 ( .A(n543), .B(n542), .ZN(n547) );
  XNOR2_X1 U661 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U662 ( .A(n547), .B(n546), .ZN(n553) );
  INV_X1 U663 ( .A(n548), .ZN(n551) );
  XNOR2_X1 U664 ( .A(n561), .B(n484), .ZN(n550) );
  NOR2_X1 U665 ( .A1(G902), .A2(n746), .ZN(n554) );
  INV_X1 U666 ( .A(n599), .ZN(n573) );
  NAND2_X1 U667 ( .A1(n572), .A2(n573), .ZN(n641) );
  NOR2_X1 U668 ( .A1(n596), .A2(n641), .ZN(n570) );
  XNOR2_X1 U669 ( .A(n566), .B(n565), .ZN(n735) );
  NOR2_X1 U670 ( .A1(n735), .A2(n622), .ZN(n569) );
  NAND2_X1 U671 ( .A1(G210), .A2(n567), .ZN(n568) );
  XNOR2_X1 U672 ( .A(n569), .B(n568), .ZN(n579) );
  NAND2_X1 U673 ( .A1(n570), .A2(n618), .ZN(n571) );
  XOR2_X1 U674 ( .A(KEYINPUT110), .B(n571), .Z(n784) );
  NOR2_X1 U675 ( .A1(KEYINPUT80), .A2(n681), .ZN(n574) );
  NOR2_X1 U676 ( .A1(n784), .A2(n574), .ZN(n593) );
  XOR2_X1 U677 ( .A(n605), .B(KEYINPUT111), .Z(n577) );
  NAND2_X1 U678 ( .A1(n579), .A2(n677), .ZN(n580) );
  INV_X1 U679 ( .A(KEYINPUT19), .ZN(n581) );
  BUF_X1 U680 ( .A(n587), .Z(n723) );
  NAND2_X1 U681 ( .A1(n723), .A2(KEYINPUT79), .ZN(n586) );
  OR2_X1 U682 ( .A1(KEYINPUT79), .A2(n587), .ZN(n583) );
  NAND2_X1 U683 ( .A1(n681), .A2(KEYINPUT80), .ZN(n582) );
  NAND2_X1 U684 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U685 ( .A1(n584), .A2(KEYINPUT47), .ZN(n585) );
  NAND2_X1 U686 ( .A1(n586), .A2(n585), .ZN(n591) );
  NOR2_X1 U687 ( .A1(KEYINPUT79), .A2(n588), .ZN(n589) );
  NOR2_X1 U688 ( .A1(KEYINPUT47), .A2(n589), .ZN(n590) );
  INV_X1 U689 ( .A(KEYINPUT38), .ZN(n595) );
  INV_X1 U690 ( .A(n600), .ZN(n676) );
  NAND2_X1 U691 ( .A1(n599), .A2(n598), .ZN(n679) );
  XNOR2_X1 U692 ( .A(KEYINPUT41), .B(n601), .ZN(n709) );
  XNOR2_X1 U693 ( .A(KEYINPUT46), .B(KEYINPUT85), .ZN(n604) );
  XOR2_X1 U694 ( .A(KEYINPUT90), .B(n686), .Z(n632) );
  NAND2_X1 U695 ( .A1(n722), .A2(n606), .ZN(n607) );
  NOR2_X1 U696 ( .A1(n645), .A2(n607), .ZN(n614) );
  INV_X1 U697 ( .A(n614), .ZN(n609) );
  NOR2_X1 U698 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U699 ( .A(KEYINPUT36), .B(n610), .Z(n611) );
  NAND2_X1 U700 ( .A1(n614), .A2(n677), .ZN(n615) );
  NOR2_X1 U701 ( .A1(n686), .A2(n615), .ZN(n616) );
  NOR2_X1 U702 ( .A1(n618), .A2(n617), .ZN(n734) );
  NAND2_X1 U703 ( .A1(n619), .A2(n718), .ZN(n732) );
  INV_X1 U704 ( .A(n690), .ZN(n647) );
  INV_X1 U705 ( .A(n679), .ZN(n630) );
  INV_X1 U706 ( .A(n624), .ZN(n627) );
  XNOR2_X1 U707 ( .A(G898), .B(KEYINPUT95), .ZN(n755) );
  NAND2_X1 U708 ( .A1(G953), .A2(n755), .ZN(n762) );
  NOR2_X1 U709 ( .A1(n625), .A2(n762), .ZN(n626) );
  NOR2_X1 U710 ( .A1(n627), .A2(n626), .ZN(n628) );
  INV_X1 U711 ( .A(n628), .ZN(n629) );
  NAND2_X1 U712 ( .A1(n645), .A2(n690), .ZN(n631) );
  NOR2_X1 U713 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U714 ( .A(n636), .B(KEYINPUT65), .ZN(n637) );
  OR2_X1 U715 ( .A1(KEYINPUT87), .A2(KEYINPUT44), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n686), .A2(n687), .ZN(n651) );
  XOR2_X1 U717 ( .A(KEYINPUT89), .B(KEYINPUT107), .Z(n640) );
  INV_X1 U718 ( .A(n641), .ZN(n642) );
  INV_X1 U719 ( .A(KEYINPUT44), .ZN(n643) );
  NAND2_X1 U720 ( .A1(n778), .A2(n643), .ZN(n644) );
  INV_X1 U721 ( .A(n645), .ZN(n650) );
  BUF_X1 U722 ( .A(n646), .Z(n648) );
  NAND2_X1 U723 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U724 ( .A1(n650), .A2(n649), .ZN(n712) );
  NAND2_X1 U725 ( .A1(n778), .A2(KEYINPUT44), .ZN(n660) );
  NOR2_X1 U726 ( .A1(n693), .A2(n651), .ZN(n699) );
  INV_X1 U727 ( .A(n655), .ZN(n652) );
  NOR2_X1 U728 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U729 ( .A1(n693), .A2(n656), .ZN(n714) );
  NAND2_X1 U730 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U731 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U732 ( .A1(n673), .A2(KEYINPUT2), .ZN(n663) );
  INV_X1 U733 ( .A(n664), .ZN(n665) );
  XNOR2_X1 U734 ( .A(n666), .B(n665), .ZN(n668) );
  NAND2_X1 U735 ( .A1(n668), .A2(n447), .ZN(n669) );
  XNOR2_X1 U736 ( .A(n669), .B(KEYINPUT123), .ZN(G63) );
  INV_X1 U737 ( .A(KEYINPUT63), .ZN(n672) );
  INV_X1 U738 ( .A(n673), .ZN(n756) );
  NOR2_X1 U739 ( .A1(n756), .A2(n674), .ZN(n675) );
  NOR2_X1 U740 ( .A1(n600), .A2(n677), .ZN(n678) );
  NOR2_X1 U741 ( .A1(n679), .A2(n678), .ZN(n683) );
  NOR2_X1 U742 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U743 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U744 ( .A(n684), .B(KEYINPUT118), .ZN(n685) );
  NOR2_X1 U745 ( .A1(n708), .A2(n685), .ZN(n704) );
  XNOR2_X1 U746 ( .A(KEYINPUT51), .B(KEYINPUT117), .ZN(n701) );
  XOR2_X1 U747 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n689) );
  OR2_X1 U748 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U749 ( .A(n689), .B(n688), .ZN(n697) );
  AND2_X1 U750 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U751 ( .A(KEYINPUT49), .B(n692), .ZN(n694) );
  NAND2_X1 U752 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U753 ( .A(KEYINPUT115), .B(n695), .Z(n696) );
  NOR2_X1 U754 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U755 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U756 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U757 ( .A1(n702), .A2(n709), .ZN(n703) );
  NOR2_X1 U758 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U759 ( .A(n705), .B(KEYINPUT52), .ZN(n706) );
  NOR2_X1 U760 ( .A1(n707), .A2(n706), .ZN(n710) );
  NOR2_X1 U761 ( .A1(n710), .A2(n386), .ZN(n711) );
  XOR2_X1 U762 ( .A(G101), .B(n712), .Z(G3) );
  INV_X1 U763 ( .A(n722), .ZN(n725) );
  NOR2_X1 U764 ( .A1(n725), .A2(n714), .ZN(n713) );
  XOR2_X1 U765 ( .A(G104), .B(n713), .Z(G6) );
  INV_X1 U766 ( .A(n718), .ZN(n728) );
  NOR2_X1 U767 ( .A1(n728), .A2(n714), .ZN(n716) );
  XNOR2_X1 U768 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n715) );
  XNOR2_X1 U769 ( .A(n716), .B(n715), .ZN(n717) );
  XNOR2_X1 U770 ( .A(G107), .B(n717), .ZN(G9) );
  XOR2_X1 U771 ( .A(KEYINPUT29), .B(KEYINPUT113), .Z(n720) );
  NAND2_X1 U772 ( .A1(n718), .A2(n723), .ZN(n719) );
  XNOR2_X1 U773 ( .A(n720), .B(n719), .ZN(n721) );
  XOR2_X1 U774 ( .A(G128), .B(n721), .Z(G30) );
  NAND2_X1 U775 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U776 ( .A(n724), .B(G146), .ZN(G48) );
  NOR2_X1 U777 ( .A1(n725), .A2(n727), .ZN(n726) );
  XOR2_X1 U778 ( .A(G113), .B(n726), .Z(G15) );
  NOR2_X1 U779 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U780 ( .A(G116), .B(n729), .Z(G18) );
  XNOR2_X1 U781 ( .A(G125), .B(n730), .ZN(n731) );
  XNOR2_X1 U782 ( .A(n731), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U783 ( .A(G134), .B(KEYINPUT114), .ZN(n733) );
  XNOR2_X1 U784 ( .A(n733), .B(n732), .ZN(G36) );
  XOR2_X1 U785 ( .A(G140), .B(n734), .Z(G42) );
  BUF_X1 U786 ( .A(n735), .Z(n737) );
  XOR2_X1 U787 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n736) );
  XOR2_X1 U788 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n740) );
  XNOR2_X1 U789 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n739) );
  XNOR2_X1 U790 ( .A(n740), .B(n739), .ZN(n741) );
  XOR2_X1 U791 ( .A(n742), .B(n741), .Z(n744) );
  XNOR2_X1 U792 ( .A(n744), .B(n743), .ZN(n745) );
  NOR2_X1 U793 ( .A1(n752), .A2(n745), .ZN(G54) );
  XOR2_X1 U794 ( .A(KEYINPUT59), .B(KEYINPUT66), .Z(n748) );
  XNOR2_X1 U795 ( .A(n746), .B(KEYINPUT91), .ZN(n747) );
  XNOR2_X1 U796 ( .A(n750), .B(n749), .ZN(n751) );
  NOR2_X1 U797 ( .A1(n752), .A2(n751), .ZN(G66) );
  NAND2_X1 U798 ( .A1(G953), .A2(G224), .ZN(n753) );
  XOR2_X1 U799 ( .A(KEYINPUT61), .B(n753), .Z(n754) );
  NOR2_X1 U800 ( .A1(n755), .A2(n754), .ZN(n758) );
  NOR2_X1 U801 ( .A1(G953), .A2(n756), .ZN(n757) );
  NOR2_X1 U802 ( .A1(n758), .A2(n757), .ZN(n765) );
  XNOR2_X1 U803 ( .A(n396), .B(G101), .ZN(n760) );
  XNOR2_X1 U804 ( .A(n760), .B(KEYINPUT124), .ZN(n761) );
  XNOR2_X1 U805 ( .A(n761), .B(G110), .ZN(n763) );
  NAND2_X1 U806 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U807 ( .A(n765), .B(n764), .ZN(G69) );
  XNOR2_X1 U808 ( .A(n766), .B(n767), .ZN(n769) );
  XNOR2_X1 U809 ( .A(n769), .B(n768), .ZN(n773) );
  XOR2_X1 U810 ( .A(n773), .B(n674), .Z(n770) );
  NOR2_X1 U811 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U812 ( .A(n772), .B(KEYINPUT125), .ZN(n777) );
  XNOR2_X1 U813 ( .A(G227), .B(n773), .ZN(n774) );
  NAND2_X1 U814 ( .A1(n774), .A2(G900), .ZN(n775) );
  NAND2_X1 U815 ( .A1(n775), .A2(G953), .ZN(n776) );
  NAND2_X1 U816 ( .A1(n777), .A2(n776), .ZN(G72) );
  XOR2_X1 U817 ( .A(G122), .B(n778), .Z(n779) );
  XNOR2_X1 U818 ( .A(KEYINPUT126), .B(n779), .ZN(G24) );
  XNOR2_X1 U819 ( .A(G119), .B(n780), .ZN(G21) );
  XNOR2_X1 U820 ( .A(G137), .B(KEYINPUT127), .ZN(n782) );
  XNOR2_X1 U821 ( .A(n782), .B(n781), .ZN(G39) );
  XOR2_X1 U822 ( .A(n783), .B(G131), .Z(G33) );
  XOR2_X1 U823 ( .A(G143), .B(n784), .Z(G45) );
  BUF_X1 U824 ( .A(n785), .Z(n786) );
  XNOR2_X1 U825 ( .A(G110), .B(n786), .ZN(G12) );
endmodule

