

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721;

  OR2_X1 U365 ( .A1(n649), .A2(n444), .ZN(n447) );
  XNOR2_X1 U366 ( .A(n386), .B(G125), .ZN(n421) );
  INV_X1 U367 ( .A(G146), .ZN(n386) );
  INV_X1 U368 ( .A(G953), .ZN(n712) );
  BUF_X1 U369 ( .A(n630), .Z(n705) );
  AND2_X1 U370 ( .A1(n353), .A2(n599), .ZN(n510) );
  NAND2_X1 U371 ( .A1(n536), .A2(n491), .ZN(n404) );
  BUF_X1 U372 ( .A(n532), .Z(n575) );
  XNOR2_X2 U373 ( .A(n347), .B(n344), .ZN(n631) );
  AND2_X2 U374 ( .A1(n510), .A2(n517), .ZN(n509) );
  AND2_X1 U375 ( .A1(n350), .A2(n368), .ZN(n349) );
  XNOR2_X1 U376 ( .A(n560), .B(n559), .ZN(n721) );
  AND2_X1 U377 ( .A1(n578), .A2(n363), .ZN(n560) );
  AND2_X1 U378 ( .A1(n485), .A2(n484), .ZN(n641) );
  NOR2_X1 U379 ( .A1(n707), .A2(G902), .ZN(n400) );
  INV_X1 U380 ( .A(n352), .ZN(n341) );
  XNOR2_X1 U381 ( .A(n354), .B(n346), .ZN(n662) );
  XNOR2_X1 U382 ( .A(n522), .B(n521), .ZN(n342) );
  XNOR2_X1 U383 ( .A(n522), .B(n521), .ZN(n618) );
  BUF_X1 U384 ( .A(n617), .Z(n343) );
  AND2_X1 U385 ( .A1(n565), .A2(n345), .ZN(n367) );
  NOR2_X1 U386 ( .A1(n448), .A2(n449), .ZN(n351) );
  XNOR2_X1 U387 ( .A(n359), .B(n357), .ZN(n490) );
  XNOR2_X1 U388 ( .A(n461), .B(n358), .ZN(n357) );
  OR2_X1 U389 ( .A1(n702), .A2(G902), .ZN(n359) );
  XNOR2_X1 U390 ( .A(n455), .B(n454), .ZN(n458) );
  XNOR2_X1 U391 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U392 ( .A(n356), .B(n355), .ZN(n455) );
  NAND2_X1 U393 ( .A1(n488), .A2(n667), .ZN(n353) );
  INV_X1 U394 ( .A(KEYINPUT102), .ZN(n358) );
  XNOR2_X1 U395 ( .A(G101), .B(G146), .ZN(n406) );
  XNOR2_X1 U396 ( .A(n451), .B(KEYINPUT100), .ZN(n356) );
  XNOR2_X1 U397 ( .A(G107), .B(KEYINPUT7), .ZN(n451) );
  XNOR2_X1 U398 ( .A(KEYINPUT9), .B(KEYINPUT101), .ZN(n355) );
  XNOR2_X1 U399 ( .A(n385), .B(n384), .ZN(n482) );
  NAND2_X2 U400 ( .A1(n364), .A2(n374), .ZN(n711) );
  XNOR2_X1 U401 ( .A(n366), .B(n365), .ZN(n364) );
  INV_X1 U402 ( .A(KEYINPUT48), .ZN(n365) );
  XNOR2_X1 U403 ( .A(G119), .B(G116), .ZN(n410) );
  XNOR2_X1 U404 ( .A(G119), .B(G128), .ZN(n388) );
  XNOR2_X1 U405 ( .A(G140), .B(KEYINPUT10), .ZN(n387) );
  XNOR2_X1 U406 ( .A(n380), .B(n379), .ZN(n429) );
  XNOR2_X1 U407 ( .A(G104), .B(G101), .ZN(n380) );
  XNOR2_X1 U408 ( .A(G110), .B(G107), .ZN(n379) );
  XNOR2_X1 U409 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U410 ( .A(n360), .B(KEYINPUT108), .ZN(n571) );
  NAND2_X1 U411 ( .A1(n363), .A2(n361), .ZN(n360) );
  AND2_X1 U412 ( .A1(n362), .A2(n548), .ZN(n361) );
  NAND2_X1 U413 ( .A1(n352), .A2(n351), .ZN(n348) );
  NAND2_X1 U414 ( .A1(n448), .A2(n449), .ZN(n368) );
  NOR2_X1 U415 ( .A1(n480), .A2(n484), .ZN(n686) );
  XNOR2_X1 U416 ( .A(n459), .B(n460), .ZN(n702) );
  XOR2_X1 U417 ( .A(n429), .B(n383), .Z(n344) );
  OR2_X1 U418 ( .A1(n490), .A2(n487), .ZN(n558) );
  INV_X1 U419 ( .A(n558), .ZN(n363) );
  XOR2_X1 U420 ( .A(n569), .B(KEYINPUT73), .Z(n345) );
  XOR2_X1 U421 ( .A(KEYINPUT106), .B(KEYINPUT33), .Z(n346) );
  XNOR2_X1 U422 ( .A(n347), .B(n710), .ZN(n714) );
  XNOR2_X2 U423 ( .A(n415), .B(n391), .ZN(n347) );
  NAND2_X1 U424 ( .A1(n349), .A2(n348), .ZN(n370) );
  NAND2_X1 U425 ( .A1(n662), .A2(n449), .ZN(n350) );
  INV_X1 U426 ( .A(n662), .ZN(n352) );
  NAND2_X1 U427 ( .A1(n510), .A2(n515), .ZN(n511) );
  NAND2_X1 U428 ( .A1(n418), .A2(n362), .ZN(n354) );
  NOR2_X1 U429 ( .A1(n571), .A2(n549), .ZN(n550) );
  INV_X1 U430 ( .A(n547), .ZN(n362) );
  NAND2_X1 U431 ( .A1(n566), .A2(n367), .ZN(n366) );
  XNOR2_X2 U432 ( .A(n369), .B(n479), .ZN(n617) );
  NAND2_X1 U433 ( .A1(n370), .A2(n478), .ZN(n369) );
  XNOR2_X2 U434 ( .A(n405), .B(KEYINPUT75), .ZN(n480) );
  BUF_X1 U435 ( .A(n482), .Z(n541) );
  NOR2_X2 U436 ( .A1(n496), .A2(n675), .ZN(n405) );
  BUF_X1 U437 ( .A(n660), .Z(n661) );
  OR2_X1 U438 ( .A1(n603), .A2(G902), .ZN(n371) );
  XOR2_X1 U439 ( .A(n399), .B(n398), .Z(n372) );
  XOR2_X1 U440 ( .A(n591), .B(n590), .Z(n373) );
  AND2_X1 U441 ( .A1(n600), .A2(n659), .ZN(n374) );
  INV_X1 U442 ( .A(KEYINPUT76), .ZN(n581) );
  XNOR2_X1 U443 ( .A(n711), .B(n581), .ZN(n583) );
  XNOR2_X1 U444 ( .A(n423), .B(n422), .ZN(n426) );
  XNOR2_X1 U445 ( .A(n421), .B(n387), .ZN(n710) );
  INV_X1 U446 ( .A(n709), .ZN(n594) );
  XNOR2_X2 U447 ( .A(G128), .B(KEYINPUT83), .ZN(n375) );
  XNOR2_X2 U448 ( .A(n375), .B(G143), .ZN(n456) );
  INV_X1 U449 ( .A(KEYINPUT64), .ZN(n376) );
  XNOR2_X1 U450 ( .A(n376), .B(KEYINPUT4), .ZN(n377) );
  XNOR2_X2 U451 ( .A(n456), .B(n377), .ZN(n424) );
  XNOR2_X1 U452 ( .A(G134), .B(G131), .ZN(n378) );
  XNOR2_X2 U453 ( .A(n424), .B(n378), .ZN(n415) );
  XNOR2_X1 U454 ( .A(G137), .B(KEYINPUT70), .ZN(n391) );
  NAND2_X1 U455 ( .A1(G227), .A2(n712), .ZN(n382) );
  XOR2_X1 U456 ( .A(G146), .B(G140), .Z(n381) );
  XNOR2_X1 U457 ( .A(n382), .B(n381), .ZN(n383) );
  INV_X1 U458 ( .A(G902), .ZN(n434) );
  NAND2_X1 U459 ( .A1(n631), .A2(n434), .ZN(n385) );
  INV_X1 U460 ( .A(G469), .ZN(n384) );
  XNOR2_X1 U461 ( .A(n482), .B(KEYINPUT1), .ZN(n496) );
  XOR2_X1 U462 ( .A(KEYINPUT23), .B(G110), .Z(n389) );
  XNOR2_X1 U463 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U464 ( .A(n710), .B(n390), .ZN(n396) );
  XNOR2_X1 U465 ( .A(n391), .B(KEYINPUT24), .ZN(n394) );
  NAND2_X1 U466 ( .A1(G234), .A2(n712), .ZN(n392) );
  XOR2_X1 U467 ( .A(KEYINPUT8), .B(n392), .Z(n450) );
  NAND2_X1 U468 ( .A1(G221), .A2(n450), .ZN(n393) );
  XNOR2_X1 U469 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U470 ( .A(n396), .B(n395), .ZN(n707) );
  XNOR2_X1 U471 ( .A(KEYINPUT15), .B(G902), .ZN(n579) );
  NAND2_X1 U472 ( .A1(G234), .A2(n579), .ZN(n397) );
  XNOR2_X1 U473 ( .A(KEYINPUT20), .B(n397), .ZN(n401) );
  NAND2_X1 U474 ( .A1(G217), .A2(n401), .ZN(n399) );
  XOR2_X1 U475 ( .A(KEYINPUT25), .B(KEYINPUT78), .Z(n398) );
  XNOR2_X2 U476 ( .A(n400), .B(n372), .ZN(n536) );
  NAND2_X1 U477 ( .A1(G221), .A2(n401), .ZN(n403) );
  INV_X1 U478 ( .A(KEYINPUT21), .ZN(n402) );
  XNOR2_X1 U479 ( .A(n403), .B(n402), .ZN(n677) );
  XNOR2_X1 U480 ( .A(n677), .B(KEYINPUT92), .ZN(n491) );
  XNOR2_X2 U481 ( .A(n404), .B(KEYINPUT68), .ZN(n675) );
  XNOR2_X1 U482 ( .A(n480), .B(KEYINPUT105), .ZN(n418) );
  XOR2_X1 U483 ( .A(G137), .B(KEYINPUT5), .Z(n407) );
  XNOR2_X1 U484 ( .A(n407), .B(n406), .ZN(n409) );
  NOR2_X1 U485 ( .A1(G953), .A2(G237), .ZN(n470) );
  NAND2_X1 U486 ( .A1(n470), .A2(G210), .ZN(n408) );
  XNOR2_X1 U487 ( .A(n409), .B(n408), .ZN(n413) );
  XNOR2_X1 U488 ( .A(n410), .B(KEYINPUT3), .ZN(n412) );
  XNOR2_X1 U489 ( .A(G113), .B(KEYINPUT71), .ZN(n411) );
  XNOR2_X1 U490 ( .A(n412), .B(n411), .ZN(n430) );
  XNOR2_X1 U491 ( .A(n413), .B(n430), .ZN(n414) );
  XNOR2_X1 U492 ( .A(n415), .B(n414), .ZN(n591) );
  OR2_X2 U493 ( .A1(n591), .A2(G902), .ZN(n416) );
  XNOR2_X2 U494 ( .A(n416), .B(G472), .ZN(n681) );
  XNOR2_X1 U495 ( .A(KEYINPUT104), .B(KEYINPUT6), .ZN(n417) );
  XNOR2_X1 U496 ( .A(n681), .B(n417), .ZN(n547) );
  NAND2_X1 U497 ( .A1(n712), .A2(G224), .ZN(n419) );
  XNOR2_X1 U498 ( .A(n419), .B(KEYINPUT79), .ZN(n423) );
  XNOR2_X1 U499 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n420) );
  INV_X1 U500 ( .A(n424), .ZN(n425) );
  XNOR2_X1 U501 ( .A(n426), .B(n425), .ZN(n432) );
  XNOR2_X1 U502 ( .A(KEYINPUT72), .B(KEYINPUT16), .ZN(n427) );
  XNOR2_X1 U503 ( .A(n427), .B(G122), .ZN(n428) );
  XNOR2_X1 U504 ( .A(n429), .B(n428), .ZN(n431) );
  XNOR2_X1 U505 ( .A(n431), .B(n430), .ZN(n627) );
  XNOR2_X1 U506 ( .A(n432), .B(n627), .ZN(n611) );
  INV_X1 U507 ( .A(n579), .ZN(n585) );
  OR2_X2 U508 ( .A1(n611), .A2(n585), .ZN(n437) );
  INV_X1 U509 ( .A(G237), .ZN(n433) );
  NAND2_X1 U510 ( .A1(n434), .A2(n433), .ZN(n438) );
  NAND2_X1 U511 ( .A1(n438), .A2(G210), .ZN(n435) );
  XNOR2_X1 U512 ( .A(n435), .B(KEYINPUT89), .ZN(n436) );
  XNOR2_X2 U513 ( .A(n437), .B(n436), .ZN(n532) );
  NAND2_X1 U514 ( .A1(n438), .A2(G214), .ZN(n663) );
  NAND2_X1 U515 ( .A1(n532), .A2(n663), .ZN(n549) );
  INV_X1 U516 ( .A(KEYINPUT19), .ZN(n439) );
  XNOR2_X2 U517 ( .A(n549), .B(n439), .ZN(n649) );
  NAND2_X1 U518 ( .A1(G234), .A2(G237), .ZN(n440) );
  XNOR2_X1 U519 ( .A(n440), .B(KEYINPUT14), .ZN(n441) );
  NAND2_X1 U520 ( .A1(G952), .A2(n441), .ZN(n694) );
  NOR2_X1 U521 ( .A1(G953), .A2(n694), .ZN(n526) );
  NAND2_X1 U522 ( .A1(G902), .A2(n441), .ZN(n523) );
  XOR2_X1 U523 ( .A(G898), .B(KEYINPUT90), .Z(n623) );
  NAND2_X1 U524 ( .A1(G953), .A2(n623), .ZN(n626) );
  NOR2_X1 U525 ( .A1(n523), .A2(n626), .ZN(n442) );
  OR2_X1 U526 ( .A1(n526), .A2(n442), .ZN(n443) );
  XNOR2_X1 U527 ( .A(n443), .B(KEYINPUT91), .ZN(n444) );
  INV_X1 U528 ( .A(KEYINPUT66), .ZN(n445) );
  XNOR2_X1 U529 ( .A(n445), .B(KEYINPUT0), .ZN(n446) );
  XNOR2_X2 U530 ( .A(n447), .B(n446), .ZN(n494) );
  INV_X1 U531 ( .A(n494), .ZN(n448) );
  INV_X1 U532 ( .A(KEYINPUT34), .ZN(n449) );
  NAND2_X1 U533 ( .A1(n450), .A2(G217), .ZN(n460) );
  XNOR2_X1 U534 ( .A(G116), .B(G122), .ZN(n453) );
  INV_X1 U535 ( .A(KEYINPUT99), .ZN(n452) );
  XNOR2_X1 U536 ( .A(n456), .B(G134), .ZN(n457) );
  XNOR2_X1 U537 ( .A(n458), .B(n457), .ZN(n459) );
  INV_X1 U538 ( .A(G478), .ZN(n461) );
  XOR2_X1 U539 ( .A(KEYINPUT98), .B(KEYINPUT13), .Z(n463) );
  XNOR2_X1 U540 ( .A(KEYINPUT97), .B(G475), .ZN(n462) );
  XNOR2_X1 U541 ( .A(n463), .B(n462), .ZN(n476) );
  XOR2_X1 U542 ( .A(G122), .B(G104), .Z(n465) );
  XNOR2_X1 U543 ( .A(G113), .B(G143), .ZN(n464) );
  XNOR2_X1 U544 ( .A(n465), .B(n464), .ZN(n469) );
  XOR2_X1 U545 ( .A(KEYINPUT96), .B(KEYINPUT12), .Z(n467) );
  XNOR2_X1 U546 ( .A(KEYINPUT11), .B(KEYINPUT95), .ZN(n466) );
  XNOR2_X1 U547 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U548 ( .A(n469), .B(n468), .ZN(n474) );
  XOR2_X1 U549 ( .A(G131), .B(KEYINPUT94), .Z(n472) );
  NAND2_X1 U550 ( .A1(G214), .A2(n470), .ZN(n471) );
  XNOR2_X1 U551 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U552 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U553 ( .A(n710), .B(n475), .ZN(n603) );
  XNOR2_X1 U554 ( .A(n476), .B(n371), .ZN(n487) );
  INV_X1 U555 ( .A(n487), .ZN(n489) );
  NAND2_X1 U556 ( .A1(n490), .A2(n489), .ZN(n477) );
  XNOR2_X1 U557 ( .A(n477), .B(KEYINPUT107), .ZN(n533) );
  XNOR2_X1 U558 ( .A(n533), .B(KEYINPUT80), .ZN(n478) );
  INV_X1 U559 ( .A(KEYINPUT35), .ZN(n479) );
  INV_X1 U560 ( .A(n681), .ZN(n484) );
  NAND2_X1 U561 ( .A1(n686), .A2(n494), .ZN(n481) );
  XNOR2_X1 U562 ( .A(n481), .B(KEYINPUT31), .ZN(n655) );
  NOR2_X2 U563 ( .A1(n675), .A2(n541), .ZN(n529) );
  NAND2_X1 U564 ( .A1(n494), .A2(n529), .ZN(n483) );
  XNOR2_X1 U565 ( .A(n483), .B(KEYINPUT93), .ZN(n485) );
  OR2_X2 U566 ( .A1(n655), .A2(n641), .ZN(n488) );
  NAND2_X1 U567 ( .A1(n490), .A2(n487), .ZN(n486) );
  XOR2_X1 U568 ( .A(n486), .B(KEYINPUT103), .Z(n577) );
  NAND2_X1 U569 ( .A1(n577), .A2(n558), .ZN(n667) );
  OR2_X1 U570 ( .A1(n490), .A2(n489), .ZN(n666) );
  INV_X1 U571 ( .A(n491), .ZN(n492) );
  NOR2_X1 U572 ( .A1(n666), .A2(n492), .ZN(n493) );
  NAND2_X1 U573 ( .A1(n494), .A2(n493), .ZN(n495) );
  XNOR2_X1 U574 ( .A(n495), .B(KEYINPUT22), .ZN(n508) );
  BUF_X1 U575 ( .A(n496), .Z(n497) );
  INV_X1 U576 ( .A(n497), .ZN(n570) );
  AND2_X1 U577 ( .A1(n497), .A2(n536), .ZN(n498) );
  NAND2_X1 U578 ( .A1(n498), .A2(n547), .ZN(n499) );
  OR2_X1 U579 ( .A1(n508), .A2(n499), .ZN(n599) );
  NOR2_X1 U580 ( .A1(n497), .A2(n536), .ZN(n500) );
  NAND2_X1 U581 ( .A1(n500), .A2(n547), .ZN(n501) );
  XNOR2_X1 U582 ( .A(n501), .B(KEYINPUT82), .ZN(n502) );
  OR2_X2 U583 ( .A1(n502), .A2(n508), .ZN(n505) );
  INV_X1 U584 ( .A(KEYINPUT81), .ZN(n503) );
  XNOR2_X1 U585 ( .A(n503), .B(KEYINPUT32), .ZN(n504) );
  XNOR2_X2 U586 ( .A(n505), .B(n504), .ZN(n608) );
  NOR2_X1 U587 ( .A1(n536), .A2(n681), .ZN(n506) );
  NAND2_X1 U588 ( .A1(n497), .A2(n506), .ZN(n507) );
  OR2_X1 U589 ( .A1(n508), .A2(n507), .ZN(n597) );
  AND2_X2 U590 ( .A1(n608), .A2(n597), .ZN(n517) );
  NAND2_X1 U591 ( .A1(n617), .A2(n509), .ZN(n512) );
  NAND2_X1 U592 ( .A1(n512), .A2(n511), .ZN(n514) );
  INV_X1 U593 ( .A(KEYINPUT87), .ZN(n513) );
  XNOR2_X1 U594 ( .A(n514), .B(n513), .ZN(n520) );
  INV_X1 U595 ( .A(KEYINPUT44), .ZN(n515) );
  NAND2_X1 U596 ( .A1(n617), .A2(n515), .ZN(n516) );
  XNOR2_X1 U597 ( .A(n516), .B(KEYINPUT67), .ZN(n518) );
  NAND2_X1 U598 ( .A1(n518), .A2(n517), .ZN(n519) );
  NAND2_X1 U599 ( .A1(n520), .A2(n519), .ZN(n522) );
  XNOR2_X1 U600 ( .A(KEYINPUT85), .B(KEYINPUT45), .ZN(n521) );
  OR2_X1 U601 ( .A1(n712), .A2(n523), .ZN(n524) );
  NOR2_X1 U602 ( .A1(G900), .A2(n524), .ZN(n525) );
  NOR2_X1 U603 ( .A1(n526), .A2(n525), .ZN(n539) );
  NAND2_X1 U604 ( .A1(n681), .A2(n663), .ZN(n527) );
  XNOR2_X1 U605 ( .A(n527), .B(KEYINPUT30), .ZN(n528) );
  NOR2_X1 U606 ( .A1(n539), .A2(n528), .ZN(n530) );
  NAND2_X1 U607 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X2 U608 ( .A(n531), .B(KEYINPUT77), .ZN(n556) );
  NAND2_X1 U609 ( .A1(n556), .A2(n575), .ZN(n535) );
  INV_X1 U610 ( .A(n533), .ZN(n534) );
  OR2_X1 U611 ( .A1(n535), .A2(n534), .ZN(n647) );
  XNOR2_X1 U612 ( .A(n647), .B(KEYINPUT84), .ZN(n546) );
  INV_X1 U613 ( .A(n536), .ZN(n537) );
  NAND2_X1 U614 ( .A1(n677), .A2(n537), .ZN(n538) );
  NOR2_X1 U615 ( .A1(n539), .A2(n538), .ZN(n548) );
  AND2_X1 U616 ( .A1(n681), .A2(n548), .ZN(n540) );
  XOR2_X1 U617 ( .A(KEYINPUT28), .B(n540), .Z(n542) );
  NOR2_X1 U618 ( .A1(n542), .A2(n541), .ZN(n648) );
  NAND2_X1 U619 ( .A1(n667), .A2(n648), .ZN(n543) );
  NOR2_X1 U620 ( .A1(n543), .A2(n649), .ZN(n567) );
  INV_X1 U621 ( .A(n567), .ZN(n544) );
  NAND2_X1 U622 ( .A1(KEYINPUT47), .A2(n544), .ZN(n545) );
  NAND2_X1 U623 ( .A1(n546), .A2(n545), .ZN(n554) );
  INV_X1 U624 ( .A(KEYINPUT36), .ZN(n551) );
  XNOR2_X1 U625 ( .A(n551), .B(n550), .ZN(n552) );
  NOR2_X1 U626 ( .A1(n552), .A2(n497), .ZN(n657) );
  XNOR2_X1 U627 ( .A(n657), .B(KEYINPUT86), .ZN(n553) );
  NOR2_X1 U628 ( .A1(n554), .A2(n553), .ZN(n566) );
  XNOR2_X1 U629 ( .A(KEYINPUT74), .B(KEYINPUT38), .ZN(n555) );
  XOR2_X1 U630 ( .A(n555), .B(n575), .Z(n664) );
  NAND2_X1 U631 ( .A1(n556), .A2(n664), .ZN(n557) );
  XNOR2_X1 U632 ( .A(n557), .B(KEYINPUT39), .ZN(n578) );
  XNOR2_X1 U633 ( .A(KEYINPUT110), .B(KEYINPUT40), .ZN(n559) );
  NAND2_X1 U634 ( .A1(n664), .A2(n663), .ZN(n668) );
  NOR2_X1 U635 ( .A1(n668), .A2(n666), .ZN(n561) );
  XNOR2_X1 U636 ( .A(n561), .B(KEYINPUT41), .ZN(n695) );
  INV_X1 U637 ( .A(n648), .ZN(n562) );
  NOR2_X1 U638 ( .A1(n695), .A2(n562), .ZN(n563) );
  XNOR2_X1 U639 ( .A(n563), .B(KEYINPUT42), .ZN(n720) );
  NOR2_X2 U640 ( .A1(n721), .A2(n720), .ZN(n564) );
  XNOR2_X1 U641 ( .A(n564), .B(KEYINPUT46), .ZN(n565) );
  XNOR2_X1 U642 ( .A(KEYINPUT47), .B(KEYINPUT69), .ZN(n568) );
  NAND2_X1 U643 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U644 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U645 ( .A1(n663), .A2(n572), .ZN(n573) );
  XNOR2_X1 U646 ( .A(n573), .B(KEYINPUT109), .ZN(n574) );
  XNOR2_X1 U647 ( .A(n574), .B(KEYINPUT43), .ZN(n576) );
  OR2_X1 U648 ( .A1(n576), .A2(n575), .ZN(n600) );
  INV_X1 U649 ( .A(n577), .ZN(n654) );
  NAND2_X1 U650 ( .A1(n578), .A2(n654), .ZN(n659) );
  NOR2_X1 U651 ( .A1(n618), .A2(n711), .ZN(n660) );
  INV_X1 U652 ( .A(KEYINPUT2), .ZN(n582) );
  OR2_X1 U653 ( .A1(n582), .A2(n579), .ZN(n580) );
  OR2_X2 U654 ( .A1(n660), .A2(n580), .ZN(n588) );
  NAND2_X1 U655 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U656 ( .A1(n584), .A2(n342), .ZN(n586) );
  NAND2_X1 U657 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X2 U658 ( .A1(n588), .A2(n587), .ZN(n630) );
  NAND2_X1 U659 ( .A1(n630), .A2(G472), .ZN(n592) );
  XOR2_X1 U660 ( .A(KEYINPUT88), .B(KEYINPUT111), .Z(n589) );
  XNOR2_X1 U661 ( .A(n589), .B(KEYINPUT62), .ZN(n590) );
  XNOR2_X1 U662 ( .A(n592), .B(n373), .ZN(n595) );
  INV_X1 U663 ( .A(G952), .ZN(n593) );
  AND2_X1 U664 ( .A1(n593), .A2(G953), .ZN(n709) );
  NAND2_X1 U665 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U666 ( .A(n596), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U667 ( .A(n597), .B(G110), .ZN(G12) );
  XNOR2_X1 U668 ( .A(G101), .B(KEYINPUT112), .ZN(n598) );
  XNOR2_X1 U669 ( .A(n599), .B(n598), .ZN(G3) );
  XNOR2_X1 U670 ( .A(n600), .B(G140), .ZN(G42) );
  NAND2_X1 U671 ( .A1(n630), .A2(G475), .ZN(n605) );
  XOR2_X1 U672 ( .A(KEYINPUT65), .B(KEYINPUT123), .Z(n601) );
  XNOR2_X1 U673 ( .A(n601), .B(KEYINPUT59), .ZN(n602) );
  XNOR2_X1 U674 ( .A(n603), .B(n602), .ZN(n604) );
  XNOR2_X1 U675 ( .A(n605), .B(n604), .ZN(n606) );
  NOR2_X2 U676 ( .A1(n606), .A2(n709), .ZN(n607) );
  XNOR2_X1 U677 ( .A(n607), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U678 ( .A(n608), .B(G119), .ZN(G21) );
  NAND2_X1 U679 ( .A1(n630), .A2(G210), .ZN(n613) );
  XOR2_X1 U680 ( .A(KEYINPUT122), .B(KEYINPUT54), .Z(n609) );
  XNOR2_X1 U681 ( .A(n609), .B(KEYINPUT55), .ZN(n610) );
  XNOR2_X1 U682 ( .A(n611), .B(n610), .ZN(n612) );
  XNOR2_X1 U683 ( .A(n613), .B(n612), .ZN(n614) );
  NOR2_X2 U684 ( .A1(n614), .A2(n709), .ZN(n615) );
  XNOR2_X1 U685 ( .A(n615), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U686 ( .A(G122), .B(KEYINPUT125), .Z(n616) );
  XNOR2_X1 U687 ( .A(n343), .B(n616), .ZN(G24) );
  BUF_X1 U688 ( .A(n342), .Z(n619) );
  NOR2_X1 U689 ( .A1(n619), .A2(G953), .ZN(n620) );
  XNOR2_X1 U690 ( .A(n620), .B(KEYINPUT124), .ZN(n625) );
  NAND2_X1 U691 ( .A1(G953), .A2(G224), .ZN(n621) );
  XOR2_X1 U692 ( .A(KEYINPUT61), .B(n621), .Z(n622) );
  NOR2_X1 U693 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U694 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U695 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U696 ( .A(n629), .B(n628), .ZN(G69) );
  NAND2_X1 U697 ( .A1(n705), .A2(G469), .ZN(n634) );
  XNOR2_X1 U698 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n632) );
  XNOR2_X1 U699 ( .A(n631), .B(n632), .ZN(n633) );
  XNOR2_X1 U700 ( .A(n634), .B(n633), .ZN(n635) );
  NOR2_X1 U701 ( .A1(n635), .A2(n709), .ZN(G54) );
  XOR2_X1 U702 ( .A(G104), .B(KEYINPUT113), .Z(n637) );
  NAND2_X1 U703 ( .A1(n641), .A2(n363), .ZN(n636) );
  XNOR2_X1 U704 ( .A(n637), .B(n636), .ZN(G6) );
  XOR2_X1 U705 ( .A(KEYINPUT115), .B(KEYINPUT27), .Z(n639) );
  XNOR2_X1 U706 ( .A(G107), .B(KEYINPUT26), .ZN(n638) );
  XNOR2_X1 U707 ( .A(n639), .B(n638), .ZN(n640) );
  XOR2_X1 U708 ( .A(KEYINPUT114), .B(n640), .Z(n643) );
  NAND2_X1 U709 ( .A1(n641), .A2(n654), .ZN(n642) );
  XNOR2_X1 U710 ( .A(n643), .B(n642), .ZN(G9) );
  NAND2_X1 U711 ( .A1(n654), .A2(n648), .ZN(n644) );
  NOR2_X1 U712 ( .A1(n644), .A2(n649), .ZN(n646) );
  XNOR2_X1 U713 ( .A(G128), .B(KEYINPUT29), .ZN(n645) );
  XNOR2_X1 U714 ( .A(n646), .B(n645), .ZN(G30) );
  XNOR2_X1 U715 ( .A(G143), .B(n647), .ZN(G45) );
  NAND2_X1 U716 ( .A1(n648), .A2(n363), .ZN(n650) );
  NOR2_X1 U717 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U718 ( .A(G146), .B(n651), .Z(G48) );
  NAND2_X1 U719 ( .A1(n655), .A2(n363), .ZN(n652) );
  XNOR2_X1 U720 ( .A(n652), .B(KEYINPUT116), .ZN(n653) );
  XNOR2_X1 U721 ( .A(G113), .B(n653), .ZN(G15) );
  NAND2_X1 U722 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U723 ( .A(n656), .B(G116), .ZN(G18) );
  XNOR2_X1 U724 ( .A(G125), .B(n657), .ZN(n658) );
  XNOR2_X1 U725 ( .A(n658), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U726 ( .A(G134), .B(n659), .ZN(G36) );
  XNOR2_X1 U727 ( .A(n661), .B(KEYINPUT2), .ZN(n699) );
  NOR2_X1 U728 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U729 ( .A1(n666), .A2(n665), .ZN(n671) );
  INV_X1 U730 ( .A(n667), .ZN(n669) );
  NOR2_X1 U731 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U732 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U733 ( .A(n672), .B(KEYINPUT120), .ZN(n673) );
  NOR2_X1 U734 ( .A1(n341), .A2(n673), .ZN(n674) );
  XOR2_X1 U735 ( .A(KEYINPUT121), .B(n674), .Z(n691) );
  XNOR2_X1 U736 ( .A(KEYINPUT119), .B(KEYINPUT51), .ZN(n688) );
  NAND2_X1 U737 ( .A1(n675), .A2(n497), .ZN(n676) );
  XOR2_X1 U738 ( .A(KEYINPUT50), .B(n676), .Z(n684) );
  NOR2_X1 U739 ( .A1(n536), .A2(n677), .ZN(n679) );
  XNOR2_X1 U740 ( .A(KEYINPUT117), .B(KEYINPUT49), .ZN(n678) );
  XNOR2_X1 U741 ( .A(n679), .B(n678), .ZN(n680) );
  NOR2_X1 U742 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U743 ( .A(KEYINPUT118), .B(n682), .Z(n683) );
  NOR2_X1 U744 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U745 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U746 ( .A(n688), .B(n687), .ZN(n689) );
  NOR2_X1 U747 ( .A1(n689), .A2(n695), .ZN(n690) );
  NOR2_X1 U748 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U749 ( .A(n692), .B(KEYINPUT52), .ZN(n693) );
  NOR2_X1 U750 ( .A1(n694), .A2(n693), .ZN(n697) );
  NOR2_X1 U751 ( .A1(n341), .A2(n695), .ZN(n696) );
  NOR2_X1 U752 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U753 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U754 ( .A1(n700), .A2(G953), .ZN(n701) );
  XNOR2_X1 U755 ( .A(n701), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U756 ( .A1(n705), .A2(G478), .ZN(n703) );
  XNOR2_X1 U757 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U758 ( .A1(n709), .A2(n704), .ZN(G63) );
  NAND2_X1 U759 ( .A1(n705), .A2(G217), .ZN(n706) );
  XNOR2_X1 U760 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U761 ( .A1(n709), .A2(n708), .ZN(G66) );
  XNOR2_X1 U762 ( .A(n711), .B(n714), .ZN(n713) );
  NAND2_X1 U763 ( .A1(n713), .A2(n712), .ZN(n718) );
  XNOR2_X1 U764 ( .A(G227), .B(n714), .ZN(n715) );
  NAND2_X1 U765 ( .A1(n715), .A2(G900), .ZN(n716) );
  NAND2_X1 U766 ( .A1(n716), .A2(G953), .ZN(n717) );
  NAND2_X1 U767 ( .A1(n718), .A2(n717), .ZN(G72) );
  XOR2_X1 U768 ( .A(G137), .B(KEYINPUT126), .Z(n719) );
  XNOR2_X1 U769 ( .A(n720), .B(n719), .ZN(G39) );
  XOR2_X1 U770 ( .A(n721), .B(G131), .Z(G33) );
endmodule

