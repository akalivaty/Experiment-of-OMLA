//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 1 1 0 1 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT81), .B1(new_n190), .B2(G104), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT81), .ZN(new_n192));
  INV_X1    g006(.A(G104), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G107), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT82), .B(G101), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT3), .B1(new_n193), .B2(G107), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(new_n190), .A3(G104), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n195), .A2(new_n196), .A3(new_n197), .A4(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n202), .B(new_n204), .C1(KEYINPUT1), .C2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT1), .B1(new_n203), .B2(G146), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n203), .A2(G146), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n201), .A2(G143), .ZN(new_n209));
  OAI211_X1 g023(.A(G128), .B(new_n207), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n190), .A2(G104), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n193), .A2(G107), .ZN(new_n212));
  OAI21_X1  g026(.A(G101), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n200), .A2(new_n206), .A3(new_n210), .A4(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n214), .B(KEYINPUT10), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT11), .ZN(new_n216));
  INV_X1    g030(.A(G134), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n216), .B1(new_n217), .B2(G137), .ZN(new_n218));
  INV_X1    g032(.A(G137), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(KEYINPUT11), .A3(G134), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(G137), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n218), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G131), .ZN(new_n223));
  INV_X1    g037(.A(G131), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n218), .A2(new_n220), .A3(new_n224), .A4(new_n221), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(G143), .B(G146), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT0), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(new_n205), .ZN(new_n230));
  NAND2_X1  g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(KEYINPUT64), .A3(new_n231), .ZN(new_n232));
  NOR3_X1   g046(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n228), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  NOR3_X1   g049(.A1(new_n208), .A2(new_n209), .A3(new_n231), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n192), .B1(new_n193), .B2(G107), .ZN(new_n238));
  NOR3_X1   g052(.A1(new_n190), .A2(KEYINPUT81), .A3(G104), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n197), .B(new_n199), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G101), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(KEYINPUT4), .A3(new_n200), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT83), .ZN(new_n243));
  INV_X1    g057(.A(G101), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n197), .A2(new_n199), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n244), .B1(new_n245), .B2(new_n195), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n243), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  AND4_X1   g062(.A1(new_n243), .A2(new_n240), .A3(new_n247), .A4(G101), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n237), .B(new_n242), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n215), .A2(new_n227), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n227), .B1(new_n215), .B2(new_n250), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT69), .ZN(new_n253));
  INV_X1    g067(.A(G953), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(KEYINPUT69), .A2(G953), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G227), .ZN(new_n258));
  XNOR2_X1  g072(.A(G110), .B(G140), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n258), .B(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  OR3_X1    g075(.A1(new_n251), .A2(new_n252), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT85), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n200), .A2(new_n213), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n210), .A2(new_n206), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI211_X1 g080(.A(new_n263), .B(new_n227), .C1(new_n266), .C2(new_n214), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n227), .B1(new_n266), .B2(new_n214), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT85), .B1(new_n268), .B2(KEYINPUT84), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT12), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n267), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n214), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n200), .A2(new_n213), .B1(new_n206), .B2(new_n210), .ZN(new_n273));
  OAI211_X1 g087(.A(KEYINPUT84), .B(new_n226), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n270), .B1(new_n274), .B2(new_n263), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n251), .B1(new_n271), .B2(new_n276), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n262), .B(G469), .C1(new_n277), .C2(new_n260), .ZN(new_n278));
  NAND2_X1  g092(.A1(G469), .A2(G902), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  XOR2_X1   g094(.A(KEYINPUT73), .B(G902), .Z(new_n281));
  NAND3_X1  g095(.A1(new_n215), .A2(new_n250), .A3(new_n227), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n274), .A2(new_n263), .A3(new_n270), .ZN(new_n283));
  INV_X1    g097(.A(new_n267), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n282), .B(new_n260), .C1(new_n285), .C2(new_n275), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n261), .B1(new_n251), .B2(new_n252), .ZN(new_n287));
  AOI211_X1 g101(.A(G469), .B(new_n281), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n189), .B1(new_n280), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n254), .A2(G952), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n290), .B1(G234), .B2(G237), .ZN(new_n291));
  INV_X1    g105(.A(new_n281), .ZN(new_n292));
  AOI211_X1 g106(.A(new_n257), .B(new_n292), .C1(G234), .C2(G237), .ZN(new_n293));
  XOR2_X1   g107(.A(KEYINPUT21), .B(G898), .Z(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n291), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(G214), .B1(G237), .B2(G902), .ZN(new_n298));
  INV_X1    g112(.A(G119), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G116), .ZN(new_n300));
  INV_X1    g114(.A(G116), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G119), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT2), .B(G113), .ZN(new_n304));
  XOR2_X1   g118(.A(new_n303), .B(new_n304), .Z(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n306), .B(new_n242), .C1(new_n248), .C2(new_n249), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n200), .A2(new_n213), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n303), .A2(new_n304), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n300), .A2(new_n302), .A3(KEYINPUT5), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n300), .A2(KEYINPUT5), .ZN(new_n311));
  INV_X1    g125(.A(G113), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n309), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n308), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n307), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(G110), .B(G122), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n307), .A2(new_n317), .A3(new_n315), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(KEYINPUT6), .A3(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n228), .A2(KEYINPUT0), .A3(G128), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n233), .B1(new_n324), .B2(new_n231), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n322), .B1(new_n325), .B2(new_n228), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n326), .A2(KEYINPUT86), .A3(G125), .ZN(new_n327));
  INV_X1    g141(.A(G125), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n237), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT86), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n330), .B1(new_n265), .B2(new_n328), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n327), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT87), .B(G224), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n254), .ZN(new_n334));
  XOR2_X1   g148(.A(new_n332), .B(new_n334), .Z(new_n335));
  INV_X1    g149(.A(KEYINPUT6), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n316), .A2(new_n336), .A3(new_n318), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n321), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(G210), .B1(G237), .B2(G902), .ZN(new_n339));
  XOR2_X1   g153(.A(KEYINPUT88), .B(KEYINPUT7), .Z(new_n340));
  NAND2_X1  g154(.A1(new_n334), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n332), .A2(new_n341), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n210), .A2(new_n206), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT86), .B1(new_n343), .B2(G125), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n326), .A2(G125), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n346), .A2(KEYINPUT7), .A3(new_n327), .A4(new_n334), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n317), .B(KEYINPUT8), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n308), .A2(new_n314), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n308), .A2(new_n314), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n342), .A2(new_n347), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(G902), .B1(new_n352), .B2(new_n320), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n338), .A2(new_n339), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n339), .B1(new_n338), .B2(new_n353), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n297), .B(new_n298), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G237), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n257), .A2(G214), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n203), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n257), .A2(G143), .A3(G214), .A4(new_n357), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G131), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT17), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n359), .A2(new_n224), .A3(new_n360), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G140), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G125), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT16), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n328), .A2(G140), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT77), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n371), .B1(new_n366), .B2(G125), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n328), .A2(KEYINPUT77), .A3(G140), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n370), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n369), .B1(new_n374), .B2(new_n368), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G146), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n201), .B(new_n369), .C1(new_n374), .C2(new_n368), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT89), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n224), .B1(new_n359), .B2(new_n360), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT17), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n376), .A2(KEYINPUT89), .A3(new_n377), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n365), .A2(new_n380), .A3(new_n382), .A4(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT18), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n359), .B(new_n360), .C1(new_n385), .C2(new_n224), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n328), .A2(G140), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n367), .A2(new_n387), .A3(new_n201), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n388), .B1(new_n374), .B2(new_n201), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n386), .B(new_n389), .C1(new_n362), .C2(new_n385), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n384), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(G113), .B(G122), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n392), .B(new_n193), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n384), .A2(new_n393), .A3(new_n390), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G902), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  XOR2_X1   g213(.A(KEYINPUT90), .B(G475), .Z(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G478), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(KEYINPUT15), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n301), .A2(G122), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT14), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n407), .B1(new_n301), .B2(G122), .ZN(new_n408));
  OAI22_X1  g222(.A1(new_n408), .A2(KEYINPUT92), .B1(KEYINPUT14), .B2(new_n406), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n408), .A2(KEYINPUT92), .ZN(new_n410));
  OAI21_X1  g224(.A(G107), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(G116), .B(G122), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n190), .ZN(new_n413));
  XNOR2_X1  g227(.A(G128), .B(G143), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n413), .B1(new_n414), .B2(G134), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n415), .B1(G134), .B2(new_n414), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(KEYINPUT13), .B1(new_n205), .B2(G143), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n418), .A2(new_n217), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(new_n414), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n412), .B(new_n190), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT91), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n422), .B1(new_n420), .B2(new_n421), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n417), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G217), .ZN(new_n427));
  NOR3_X1   g241(.A1(new_n188), .A2(new_n427), .A3(G953), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n417), .B(new_n428), .C1(new_n424), .C2(new_n425), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n405), .B1(new_n432), .B2(new_n292), .ZN(new_n433));
  AOI211_X1 g247(.A(new_n281), .B(new_n404), .C1(new_n430), .C2(new_n431), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(G475), .A2(G902), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n367), .A2(new_n387), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n438), .A2(KEYINPUT19), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n328), .A2(KEYINPUT77), .A3(G140), .ZN(new_n440));
  AOI21_X1  g254(.A(KEYINPUT77), .B1(new_n328), .B2(G140), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n367), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n439), .B1(KEYINPUT19), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n201), .ZN(new_n444));
  INV_X1    g258(.A(new_n364), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n376), .B(new_n444), .C1(new_n445), .C2(new_n381), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n390), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n394), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n437), .B1(new_n396), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT20), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI211_X1 g265(.A(KEYINPUT20), .B(new_n437), .C1(new_n396), .C2(new_n448), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n402), .B(new_n435), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  NOR3_X1   g267(.A1(new_n289), .A2(new_n356), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT67), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT65), .ZN(new_n456));
  AOI22_X1  g270(.A1(new_n326), .A2(new_n456), .B1(new_n223), .B2(new_n225), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n322), .B(KEYINPUT65), .C1(new_n325), .C2(new_n228), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n217), .A2(G137), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n219), .A2(G134), .ZN(new_n460));
  OAI21_X1  g274(.A(G131), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n225), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n343), .A2(new_n462), .A3(KEYINPUT66), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n210), .A2(new_n225), .A3(new_n461), .A4(new_n206), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT66), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI22_X1  g280(.A1(new_n457), .A2(new_n458), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n455), .B1(new_n467), .B2(KEYINPUT30), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT30), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n464), .B(KEYINPUT66), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n456), .B1(new_n235), .B2(new_n236), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n471), .A2(new_n226), .A3(new_n458), .ZN(new_n472));
  OAI211_X1 g286(.A(KEYINPUT67), .B(new_n469), .C1(new_n470), .C2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n237), .A2(new_n226), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n343), .A2(new_n462), .A3(KEYINPUT68), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT68), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n464), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n474), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  OR2_X1    g292(.A1(new_n478), .A2(new_n469), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n468), .A2(new_n306), .A3(new_n473), .A4(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n257), .A2(G210), .A3(new_n357), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(G101), .ZN(new_n482));
  XNOR2_X1  g296(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n482), .B(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n478), .A2(new_n306), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n480), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT31), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n474), .A2(new_n464), .A3(new_n305), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT28), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(KEYINPUT71), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT70), .B(KEYINPUT28), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n467), .A2(new_n305), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n493), .B1(new_n494), .B2(new_n485), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n484), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT31), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n480), .A2(new_n499), .A3(new_n484), .A4(new_n486), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n488), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(G472), .A2(G902), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT32), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n501), .A2(KEYINPUT32), .A3(new_n502), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n496), .A2(new_n497), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n484), .B1(new_n480), .B2(new_n486), .ZN(new_n508));
  NOR3_X1   g322(.A1(new_n507), .A2(KEYINPUT29), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT72), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n478), .A2(new_n306), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n486), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n478), .A2(KEYINPUT72), .A3(new_n306), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(KEYINPUT28), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n492), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n484), .A2(KEYINPUT29), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n292), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(G472), .B1(new_n509), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n505), .A2(new_n506), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n257), .A2(G221), .A3(G234), .ZN(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT22), .B(G137), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n520), .B(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT23), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(new_n205), .A3(G119), .ZN(new_n525));
  OAI21_X1  g339(.A(KEYINPUT23), .B1(new_n299), .B2(G128), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n205), .A2(G119), .ZN(new_n527));
  OAI211_X1 g341(.A(G110), .B(new_n525), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT76), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(KEYINPUT24), .A2(G110), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT75), .ZN(new_n533));
  NAND2_X1  g347(.A1(KEYINPUT24), .A2(G110), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(KEYINPUT74), .B1(new_n205), .B2(G119), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT74), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(new_n299), .A3(G128), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AND2_X1   g353(.A1(KEYINPUT24), .A2(G110), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT75), .B1(new_n540), .B2(new_n531), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n205), .A2(G119), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n535), .A2(new_n539), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n299), .A2(G128), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n544), .A2(new_n542), .A3(KEYINPUT23), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n545), .A2(KEYINPUT76), .A3(G110), .A4(new_n525), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n530), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n547), .B1(new_n377), .B2(new_n376), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n535), .A2(new_n541), .B1(new_n539), .B2(new_n542), .ZN(new_n549));
  AOI21_X1  g363(.A(G110), .B1(new_n545), .B2(new_n525), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n388), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n442), .A2(KEYINPUT16), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n201), .B1(new_n552), .B2(new_n369), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n523), .B1(new_n548), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n547), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n378), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n376), .B(new_n388), .C1(new_n550), .C2(new_n549), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n557), .A2(new_n558), .A3(new_n522), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n555), .A2(new_n292), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT78), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n560), .A2(new_n561), .A3(KEYINPUT25), .ZN(new_n562));
  AOI21_X1  g376(.A(KEYINPUT25), .B1(new_n560), .B2(new_n561), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n427), .B1(new_n292), .B2(G234), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n564), .A2(G902), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n555), .A2(new_n559), .A3(new_n567), .ZN(new_n568));
  XOR2_X1   g382(.A(new_n568), .B(KEYINPUT79), .Z(new_n569));
  OAI21_X1  g383(.A(KEYINPUT80), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n563), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n560), .A2(new_n561), .A3(KEYINPUT25), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(new_n572), .A3(new_n564), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT80), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n568), .B(KEYINPUT79), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n454), .A2(new_n519), .A3(new_n577), .ZN(new_n578));
  XOR2_X1   g392(.A(new_n578), .B(new_n196), .Z(G3));
  NAND2_X1  g393(.A1(new_n501), .A2(new_n292), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G472), .ZN(new_n581));
  INV_X1    g395(.A(new_n189), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n251), .A2(new_n252), .A3(new_n261), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n282), .B1(new_n285), .B2(new_n275), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n583), .B1(new_n584), .B2(new_n261), .ZN(new_n585));
  OAI21_X1  g399(.A(G469), .B1(new_n585), .B2(G902), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n286), .A2(new_n287), .ZN(new_n587));
  INV_X1    g401(.A(G469), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(new_n588), .A3(new_n292), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n582), .B1(new_n586), .B2(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n581), .A2(new_n590), .A3(new_n577), .A4(new_n503), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n298), .B1(new_n354), .B2(new_n355), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT93), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT93), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n594), .B(new_n298), .C1(new_n354), .C2(new_n355), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n593), .A2(new_n297), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(G902), .B1(new_n395), .B2(new_n396), .ZN(new_n597));
  OAI22_X1  g411(.A1(new_n451), .A2(new_n452), .B1(new_n597), .B2(new_n400), .ZN(new_n598));
  AOI211_X1 g412(.A(G478), .B(new_n281), .C1(new_n430), .C2(new_n431), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT33), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n432), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n430), .A2(KEYINPUT33), .A3(new_n431), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n292), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n599), .B1(new_n603), .B2(G478), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n598), .A2(new_n604), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n591), .A2(new_n596), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT34), .B(G104), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G6));
  NAND2_X1  g422(.A1(new_n449), .A2(new_n450), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(KEYINPUT95), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT95), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n452), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n451), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT94), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n614), .A2(new_n610), .A3(new_n612), .A4(new_n615), .ZN(new_n618));
  INV_X1    g432(.A(new_n435), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n617), .A2(new_n618), .A3(new_n402), .A4(new_n619), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n591), .A2(new_n596), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT35), .B(G107), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G9));
  AOI22_X1  g437(.A1(new_n580), .A2(G472), .B1(new_n501), .B2(new_n502), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n557), .A2(new_n558), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n523), .A2(KEYINPUT36), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n567), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n573), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n454), .A2(new_n624), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT37), .B(G110), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G12));
  INV_X1    g446(.A(G900), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n291), .B1(new_n293), .B2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n620), .A2(new_n634), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n593), .A2(new_n595), .ZN(new_n636));
  INV_X1    g450(.A(new_n629), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n289), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n635), .A2(new_n636), .A3(new_n519), .A4(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G128), .ZN(G30));
  AND3_X1   g454(.A1(new_n501), .A2(KEYINPUT32), .A3(new_n502), .ZN(new_n641));
  AOI21_X1  g455(.A(KEYINPUT32), .B1(new_n501), .B2(new_n502), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n480), .A2(new_n486), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(new_n497), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n512), .A2(new_n513), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n398), .B1(new_n647), .B2(new_n484), .ZN(new_n648));
  OAI21_X1  g462(.A(G472), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n643), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(new_n650), .B(KEYINPUT96), .Z(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(new_n634), .B(KEYINPUT39), .Z(new_n653));
  NAND2_X1  g467(.A1(new_n590), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT97), .B(KEYINPUT40), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n354), .A2(new_n355), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT38), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n598), .A2(new_n619), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n659), .A2(new_n298), .A3(new_n637), .ZN(new_n660));
  OR4_X1    g474(.A1(new_n652), .A2(new_n656), .A3(new_n658), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G143), .ZN(G45));
  NOR2_X1   g476(.A1(new_n605), .A2(new_n634), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n636), .A2(new_n519), .A3(new_n638), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G146), .ZN(G48));
  INV_X1    g479(.A(new_n577), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n666), .B1(new_n643), .B2(new_n518), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n598), .A2(new_n604), .ZN(new_n668));
  AND4_X1   g482(.A1(new_n297), .A2(new_n593), .A3(new_n668), .A4(new_n595), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n587), .A2(new_n292), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(G469), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n589), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n582), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n667), .A2(new_n669), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT41), .B(G113), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G15));
  NOR2_X1   g490(.A1(new_n596), .A2(new_n620), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n673), .A2(new_n593), .A3(new_n595), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n677), .A2(new_n667), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G116), .ZN(G18));
  NOR3_X1   g494(.A1(new_n453), .A2(new_n637), .A3(new_n296), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n678), .A2(new_n519), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT98), .B(G119), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G21));
  NAND3_X1  g498(.A1(new_n593), .A2(new_n595), .A3(new_n659), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT99), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n593), .A2(KEYINPUT99), .A3(new_n659), .A4(new_n595), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n673), .A2(new_n297), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n573), .A2(new_n575), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n515), .A2(new_n497), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n692), .A2(new_n488), .A3(new_n500), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n502), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n581), .A2(new_n694), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n690), .A2(new_n691), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n689), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT100), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT100), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n689), .A2(new_n696), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G122), .ZN(G24));
  INV_X1    g516(.A(new_n634), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n668), .A2(new_n703), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n695), .A2(new_n704), .A3(new_n637), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n678), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G125), .ZN(G27));
  INV_X1    g521(.A(KEYINPUT102), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n262), .A2(new_n708), .ZN(new_n709));
  OAI211_X1 g523(.A(G469), .B(new_n709), .C1(new_n585), .C2(new_n708), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n279), .B(KEYINPUT101), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(new_n589), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n189), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT42), .ZN(new_n714));
  INV_X1    g528(.A(new_n298), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n354), .A2(new_n355), .A3(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NOR4_X1   g531(.A1(new_n713), .A2(new_n704), .A3(new_n714), .A4(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n691), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n643), .A2(KEYINPUT104), .ZN(new_n720));
  OAI21_X1  g534(.A(KEYINPUT104), .B1(new_n505), .B2(KEYINPUT32), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n518), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n718), .B(new_n719), .C1(new_n720), .C2(new_n722), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n712), .A2(new_n189), .A3(new_n716), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n724), .A2(new_n519), .A3(new_n577), .A4(new_n663), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT103), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n725), .A2(new_n726), .A3(new_n714), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n726), .B1(new_n725), .B2(new_n714), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n723), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G131), .ZN(G33));
  NAND3_X1  g544(.A1(new_n667), .A2(new_n635), .A3(new_n724), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G134), .ZN(G36));
  OAI211_X1 g546(.A(KEYINPUT45), .B(new_n709), .C1(new_n585), .C2(new_n708), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n733), .B(G469), .C1(KEYINPUT45), .C2(new_n585), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n734), .A2(new_n711), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n288), .B1(new_n735), .B2(KEYINPUT46), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n736), .A2(KEYINPUT105), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(KEYINPUT105), .ZN(new_n738));
  OAI21_X1  g552(.A(KEYINPUT106), .B1(new_n735), .B2(KEYINPUT46), .ZN(new_n739));
  OR3_X1    g553(.A1(new_n735), .A2(KEYINPUT106), .A3(KEYINPUT46), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n737), .A2(new_n738), .A3(new_n739), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n189), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n598), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n604), .ZN(new_n745));
  XOR2_X1   g559(.A(new_n745), .B(KEYINPUT43), .Z(new_n746));
  INV_X1    g560(.A(new_n624), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n747), .A3(new_n629), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n748), .A2(new_n749), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n750), .A2(new_n751), .A3(new_n717), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n743), .A2(new_n653), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G137), .ZN(G39));
  OR2_X1    g568(.A1(new_n742), .A2(KEYINPUT47), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n742), .A2(KEYINPUT47), .ZN(new_n756));
  NOR4_X1   g570(.A1(new_n519), .A2(new_n704), .A3(new_n577), .A4(new_n717), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n755), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT107), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n758), .B(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G140), .ZN(G42));
  NOR4_X1   g575(.A1(new_n745), .A2(new_n691), .A3(new_n715), .A4(new_n582), .ZN(new_n762));
  XOR2_X1   g576(.A(new_n672), .B(KEYINPUT49), .Z(new_n763));
  NAND4_X1  g577(.A1(new_n652), .A2(new_n658), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n746), .A2(new_n291), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n695), .A2(new_n691), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n755), .A2(new_n756), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n671), .A2(new_n582), .A3(new_n589), .ZN(new_n770));
  AOI211_X1 g584(.A(new_n717), .B(new_n768), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n673), .A2(new_n716), .ZN(new_n772));
  XOR2_X1   g586(.A(new_n772), .B(KEYINPUT115), .Z(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n765), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT116), .ZN(new_n775));
  OR3_X1    g589(.A1(new_n775), .A2(new_n637), .A3(new_n695), .ZN(new_n776));
  AND4_X1   g590(.A1(new_n577), .A2(new_n652), .A3(new_n291), .A4(new_n773), .ZN(new_n777));
  INV_X1    g591(.A(new_n604), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n744), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n658), .A2(new_n715), .A3(new_n673), .ZN(new_n780));
  XOR2_X1   g594(.A(new_n780), .B(KEYINPUT114), .Z(new_n781));
  NAND2_X1  g595(.A1(new_n767), .A2(new_n781), .ZN(new_n782));
  XOR2_X1   g596(.A(new_n782), .B(KEYINPUT50), .Z(new_n783));
  NAND3_X1  g597(.A1(new_n776), .A2(new_n779), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(KEYINPUT113), .B1(new_n771), .B2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n706), .A2(new_n639), .A3(new_n664), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT111), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n712), .A2(new_n189), .A3(new_n637), .A4(new_n703), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n791), .B1(new_n649), .B2(new_n643), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n790), .B1(new_n689), .B2(new_n792), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n689), .A2(new_n790), .A3(new_n792), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n789), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT53), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n679), .A2(new_n674), .A3(new_n682), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n799), .B1(new_n698), .B2(new_n700), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT109), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n356), .A2(new_n605), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n802), .A2(new_n624), .A3(new_n577), .A4(new_n590), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n578), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT108), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n578), .A2(KEYINPUT108), .A3(new_n803), .ZN(new_n807));
  INV_X1    g621(.A(new_n356), .ZN(new_n808));
  INV_X1    g622(.A(new_n453), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n808), .A2(new_n809), .A3(new_n590), .A4(new_n629), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n598), .A2(new_n435), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  OAI22_X1  g626(.A1(new_n810), .A2(new_n747), .B1(new_n591), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  AND4_X1   g628(.A1(new_n801), .A2(new_n806), .A3(new_n807), .A4(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n813), .B1(new_n804), .B2(new_n805), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n801), .B1(new_n816), .B2(new_n807), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n800), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n617), .A2(new_n618), .A3(new_n402), .ZN(new_n820));
  NOR4_X1   g634(.A1(new_n820), .A2(new_n717), .A3(new_n619), .A4(new_n634), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n519), .A2(new_n638), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n821), .A2(new_n822), .B1(new_n705), .B2(new_n724), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n729), .A2(new_n731), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n819), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n798), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT110), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n729), .A2(new_n731), .A3(new_n823), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n828), .B1(new_n818), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n806), .A2(new_n807), .A3(new_n814), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(KEYINPUT109), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n816), .A2(new_n801), .A3(new_n807), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n824), .A2(new_n834), .A3(KEYINPUT110), .A4(new_n800), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n830), .A2(new_n835), .A3(new_n797), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT112), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n837), .B1(new_n836), .B2(new_n838), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n788), .B(new_n827), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n836), .A2(new_n838), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n836), .A2(new_n838), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT54), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n290), .B(KEYINPUT117), .ZN(new_n847));
  INV_X1    g661(.A(new_n678), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n847), .B1(new_n768), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n719), .B1(new_n722), .B2(new_n720), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n775), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT48), .ZN(new_n852));
  AOI211_X1 g666(.A(new_n849), .B(new_n852), .C1(new_n668), .C2(new_n777), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n787), .A2(new_n846), .A3(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OR2_X1    g670(.A1(G952), .A2(G953), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n854), .A2(new_n855), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n764), .B1(new_n858), .B2(new_n859), .ZN(G75));
  NOR2_X1   g674(.A1(new_n257), .A2(G952), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT56), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n827), .B1(new_n839), .B2(new_n840), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n281), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n863), .B1(new_n865), .B2(new_n339), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n321), .A2(new_n337), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(new_n335), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n868), .B(KEYINPUT55), .Z(new_n869));
  AOI21_X1  g683(.A(new_n869), .B1(KEYINPUT119), .B2(new_n863), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n862), .B1(new_n866), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n871), .B1(new_n866), .B2(new_n870), .ZN(G51));
  XNOR2_X1  g686(.A(new_n587), .B(KEYINPUT120), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n864), .A2(KEYINPUT54), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n841), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n711), .B(KEYINPUT57), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n873), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OR2_X1    g692(.A1(new_n865), .A2(new_n734), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n861), .B1(new_n878), .B2(new_n879), .ZN(G54));
  AND4_X1   g694(.A1(KEYINPUT58), .A2(new_n864), .A3(G475), .A4(new_n281), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n396), .A2(new_n448), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n862), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n883), .B1(new_n882), .B2(new_n881), .ZN(G60));
  NAND2_X1  g698(.A1(new_n601), .A2(new_n602), .ZN(new_n885));
  XNOR2_X1  g699(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n403), .A2(new_n398), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n886), .B(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n861), .B1(new_n875), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n885), .B1(new_n846), .B2(new_n888), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT122), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n890), .A2(new_n891), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n893), .A2(new_n895), .ZN(G63));
  INV_X1    g710(.A(KEYINPUT124), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT61), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n862), .B1(new_n897), .B2(KEYINPUT61), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n842), .A2(KEYINPUT112), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n826), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(G217), .A2(G902), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT60), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n900), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n905), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n864), .A2(KEYINPUT123), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n899), .B1(new_n909), .B2(new_n627), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n555), .A2(new_n559), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n906), .A2(new_n911), .A3(new_n908), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n898), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n864), .A2(KEYINPUT123), .A3(new_n907), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT123), .B1(new_n864), .B2(new_n907), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n627), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n899), .ZN(new_n917));
  AND4_X1   g731(.A1(new_n898), .A2(new_n916), .A3(new_n912), .A4(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n913), .A2(new_n918), .ZN(G66));
  INV_X1    g733(.A(new_n333), .ZN(new_n920));
  OAI21_X1  g734(.A(G953), .B1(new_n295), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n257), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n921), .B1(new_n819), .B2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(G898), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n867), .B1(new_n924), .B2(new_n922), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n923), .B(new_n925), .Z(G69));
  NAND3_X1  g740(.A1(new_n468), .A2(new_n473), .A3(new_n479), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(new_n443), .Z(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n850), .B1(new_n687), .B2(new_n688), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n743), .A2(new_n653), .A3(new_n930), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n729), .A2(new_n731), .ZN(new_n932));
  AND4_X1   g746(.A1(new_n753), .A2(new_n931), .A3(new_n932), .A4(new_n789), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n922), .B1(new_n760), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT126), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n257), .A2(G900), .ZN(new_n936));
  OR3_X1    g750(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n935), .B1(new_n934), .B2(new_n936), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n929), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n257), .B1(G227), .B2(G900), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT127), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n760), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT125), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(KEYINPUT62), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n661), .A2(new_n789), .A3(new_n946), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n947), .A2(new_n945), .A3(KEYINPUT62), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n947), .B1(new_n945), .B2(KEYINPUT62), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n716), .B1(new_n668), .B2(new_n811), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n950), .A2(new_n654), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n667), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n949), .A2(new_n753), .A3(new_n952), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n944), .A2(new_n948), .A3(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n928), .A2(new_n922), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  OAI22_X1  g770(.A1(new_n954), .A2(new_n956), .B1(KEYINPUT127), .B2(new_n940), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n939), .A2(new_n943), .A3(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n943), .ZN(new_n959));
  INV_X1    g773(.A(new_n938), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n928), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n957), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n959), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n958), .A2(new_n964), .ZN(G72));
  NAND2_X1  g779(.A1(G472), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT63), .Z(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(new_n954), .B2(new_n819), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n969), .A2(new_n497), .A3(new_n645), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n843), .A2(new_n844), .ZN(new_n971));
  INV_X1    g785(.A(new_n508), .ZN(new_n972));
  AOI211_X1 g786(.A(new_n968), .B(new_n971), .C1(new_n487), .C2(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n760), .A2(new_n819), .A3(new_n933), .ZN(new_n974));
  AOI211_X1 g788(.A(new_n484), .B(new_n644), .C1(new_n974), .C2(new_n967), .ZN(new_n975));
  NOR4_X1   g789(.A1(new_n970), .A2(new_n973), .A3(new_n861), .A4(new_n975), .ZN(G57));
endmodule


