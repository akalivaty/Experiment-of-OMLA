//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1206, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1267, new_n1268, new_n1269;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  NAND2_X1  g0004(.A1(G87), .A2(G250), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT66), .ZN(new_n207));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  INV_X1    g0009(.A(G77), .ZN(new_n210));
  INV_X1    g0010(.A(G244), .ZN(new_n211));
  OAI22_X1  g0011(.A1(new_n208), .A2(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n207), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n205), .B1(new_n214), .B2(KEYINPUT67), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(KEYINPUT67), .B2(new_n214), .ZN(new_n216));
  INV_X1    g0016(.A(G58), .ZN(new_n217));
  INV_X1    g0017(.A(G232), .ZN(new_n218));
  INV_X1    g0018(.A(G97), .ZN(new_n219));
  INV_X1    g0019(.A(G257), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G107), .ZN(new_n222));
  INV_X1    g0022(.A(G264), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n204), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n204), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT0), .Z(new_n229));
  NOR2_X1   g0029(.A1(G58), .A2(G68), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(KEYINPUT65), .ZN(new_n233));
  INV_X1    g0033(.A(G20), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(KEYINPUT65), .A2(G20), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g0037(.A1(G1), .A2(G13), .ZN(new_n238));
  NOR3_X1   g0038(.A1(new_n232), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NOR3_X1   g0039(.A1(new_n226), .A2(new_n229), .A3(new_n239), .ZN(G361));
  XOR2_X1   g0040(.A(G238), .B(G244), .Z(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G226), .B(G232), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G250), .B(G257), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n223), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G270), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G358));
  XOR2_X1   g0049(.A(G68), .B(G77), .Z(new_n250));
  XNOR2_X1  g0050(.A(G50), .B(G58), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(G107), .B(G116), .Z(new_n253));
  XNOR2_X1  g0053(.A(G87), .B(G97), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n252), .B(new_n255), .ZN(G351));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n258));
  INV_X1    g0058(.A(G274), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n238), .B1(G33), .B2(G41), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n258), .ZN(new_n264));
  INV_X1    g0064(.A(G226), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n261), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(KEYINPUT3), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT3), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G33), .ZN(new_n270));
  AND2_X1   g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n271), .A2(G222), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n268), .A2(new_n270), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(new_n272), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n275), .B(KEYINPUT69), .ZN(new_n276));
  INV_X1    g0076(.A(G223), .ZN(new_n277));
  OAI221_X1 g0077(.A(new_n273), .B1(new_n210), .B2(new_n271), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n262), .B(KEYINPUT70), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n266), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  XOR2_X1   g0080(.A(KEYINPUT71), .B(G179), .Z(new_n281));
  AND2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(G20), .B1(new_n231), .B2(G50), .ZN(new_n283));
  INV_X1    g0083(.A(G150), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n237), .A2(G33), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT8), .B(G58), .ZN(new_n288));
  OAI221_X1 g0088(.A(new_n283), .B1(new_n284), .B2(new_n286), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n238), .ZN(new_n291));
  INV_X1    g0091(.A(G50), .ZN(new_n292));
  INV_X1    g0092(.A(G13), .ZN(new_n293));
  NOR3_X1   g0093(.A1(new_n293), .A2(new_n234), .A3(G1), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n289), .A2(new_n291), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n291), .B1(new_n257), .B2(G20), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n295), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n298), .B1(new_n280), .B2(G169), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n282), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n298), .B(KEYINPUT9), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n280), .A2(G190), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G200), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n280), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(KEYINPUT10), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n305), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT10), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n307), .A2(new_n301), .A3(new_n308), .A4(new_n302), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n300), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT70), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n262), .B(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(G33), .A2(G97), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n218), .A2(G1698), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n271), .B(new_n314), .C1(G226), .C2(G1698), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n312), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n261), .B1(new_n264), .B2(new_n209), .ZN(new_n317));
  NOR3_X1   g0117(.A1(new_n316), .A2(KEYINPUT13), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT13), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n315), .A2(new_n313), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n279), .ZN(new_n321));
  INV_X1    g0121(.A(new_n317), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n319), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(G169), .B1(new_n318), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT14), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n318), .A2(new_n323), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G179), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT14), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n328), .B(G169), .C1(new_n318), .C2(new_n323), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n325), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n257), .A2(new_n208), .A3(G13), .A4(G20), .ZN(new_n331));
  XOR2_X1   g0131(.A(new_n331), .B(KEYINPUT12), .Z(new_n332));
  AOI21_X1  g0132(.A(new_n332), .B1(G68), .B2(new_n296), .ZN(new_n333));
  OAI22_X1  g0133(.A1(new_n287), .A2(new_n210), .B1(new_n234), .B2(G68), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT74), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI221_X1 g0136(.A(KEYINPUT74), .B1(new_n234), .B2(G68), .C1(new_n287), .C2(new_n210), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n336), .B(new_n337), .C1(new_n292), .C2(new_n286), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT11), .ZN(new_n339));
  AND3_X1   g0139(.A1(new_n338), .A2(new_n339), .A3(new_n291), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n339), .B1(new_n338), .B2(new_n291), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n333), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n330), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(KEYINPUT13), .B1(new_n316), .B2(new_n317), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n321), .A2(new_n322), .A3(new_n319), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n344), .A2(G190), .A3(new_n345), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n333), .B(new_n346), .C1(new_n340), .C2(new_n341), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n326), .A2(new_n304), .ZN(new_n348));
  OR2_X1    g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NOR3_X1   g0149(.A1(new_n274), .A2(new_n218), .A3(G1698), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n350), .B(KEYINPUT72), .ZN(new_n351));
  OAI221_X1 g0151(.A(new_n351), .B1(new_n222), .B2(new_n271), .C1(new_n276), .C2(new_n209), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n279), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n261), .B1(new_n264), .B2(new_n211), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n353), .A2(G190), .A3(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n288), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n235), .A2(new_n236), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n357), .A2(new_n285), .B1(new_n358), .B2(G77), .ZN(new_n359));
  XOR2_X1   g0159(.A(KEYINPUT15), .B(G87), .Z(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n359), .B1(new_n287), .B2(new_n361), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n362), .A2(new_n291), .B1(G77), .B2(new_n296), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n294), .A2(new_n210), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n364), .B(KEYINPUT73), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n356), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n354), .B1(new_n352), .B2(new_n279), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n369), .A2(new_n304), .ZN(new_n370));
  OR2_X1    g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  AND4_X1   g0171(.A1(new_n310), .A2(new_n343), .A3(new_n349), .A4(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT75), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(new_n267), .B2(KEYINPUT3), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n269), .A2(KEYINPUT75), .A3(G33), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n268), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT7), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(new_n378), .A3(new_n237), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n374), .A2(new_n375), .B1(KEYINPUT3), .B2(new_n267), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT7), .B1(new_n380), .B2(G20), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n379), .A2(new_n381), .A3(G68), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n285), .A2(G159), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n383), .B(KEYINPUT76), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n217), .A2(new_n208), .ZN(new_n385));
  OAI21_X1  g0185(.A(G20), .B1(new_n385), .B2(new_n230), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n382), .A2(KEYINPUT16), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT16), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n378), .B1(new_n271), .B2(G20), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n237), .A2(new_n274), .A3(KEYINPUT7), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n208), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n384), .A2(new_n386), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n389), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n388), .A2(new_n394), .A3(new_n291), .ZN(new_n395));
  INV_X1    g0195(.A(new_n294), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n288), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n296), .B2(new_n288), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n277), .A2(new_n272), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n265), .A2(G1698), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n376), .A2(new_n268), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT77), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G33), .A2(G87), .ZN(new_n404));
  AND3_X1   g0204(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n403), .B1(new_n402), .B2(new_n404), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n279), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n263), .A2(G232), .A3(new_n258), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT78), .ZN(new_n409));
  XNOR2_X1  g0209(.A(new_n408), .B(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n407), .A2(new_n261), .A3(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(G169), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n407), .A2(new_n261), .A3(new_n281), .A4(new_n410), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n399), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT18), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT18), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n399), .A2(new_n413), .A3(new_n417), .A4(new_n414), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT17), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n411), .A2(G200), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n407), .A2(G190), .A3(new_n261), .A4(new_n410), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n424), .A2(new_n395), .A3(new_n398), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n421), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n395), .A2(new_n398), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n427), .A2(KEYINPUT17), .A3(new_n422), .A4(new_n424), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n366), .B1(new_n369), .B2(G169), .ZN(new_n431));
  INV_X1    g0231(.A(new_n281), .ZN(new_n432));
  AOI211_X1 g0232(.A(new_n432), .B(new_n354), .C1(new_n352), .C2(new_n279), .ZN(new_n433));
  OR2_X1    g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n372), .A2(new_n420), .A3(new_n430), .A4(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n376), .A2(G244), .A3(G1698), .A4(new_n268), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT80), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n209), .A2(G1698), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n380), .A2(new_n439), .B1(G33), .B2(G116), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n380), .A2(KEYINPUT80), .A3(G244), .A4(G1698), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n279), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT79), .ZN(new_n444));
  INV_X1    g0244(.A(G45), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(G1), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n444), .B1(new_n447), .B2(new_n259), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n446), .A2(KEYINPUT79), .A3(G274), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n263), .A2(G250), .A3(new_n447), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n443), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT81), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n452), .B1(new_n442), .B2(new_n279), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT81), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n455), .A2(G200), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n457), .B1(new_n443), .B2(new_n453), .ZN(new_n460));
  AOI211_X1 g0260(.A(KEYINPUT81), .B(new_n452), .C1(new_n442), .C2(new_n279), .ZN(new_n461));
  OAI21_X1  g0261(.A(G190), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n396), .A2(new_n360), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n380), .A2(G68), .A3(new_n237), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n237), .A2(G33), .A3(G97), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT19), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G87), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(new_n219), .A3(new_n222), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n313), .A2(new_n466), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n469), .B1(new_n358), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n464), .A2(new_n467), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n463), .B1(new_n472), .B2(new_n291), .ZN(new_n473));
  AOI211_X1 g0273(.A(new_n291), .B(new_n294), .C1(new_n257), .C2(G33), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G87), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n459), .A2(new_n462), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n455), .A2(new_n412), .A3(new_n458), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n281), .B1(new_n460), .B2(new_n461), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n472), .A2(new_n291), .ZN(new_n480));
  INV_X1    g0280(.A(new_n463), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n474), .A2(new_n360), .ZN(new_n482));
  AND4_X1   g0282(.A1(KEYINPUT82), .A2(new_n480), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(KEYINPUT82), .B1(new_n473), .B2(new_n482), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n478), .A2(new_n479), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n477), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT83), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n222), .B1(new_n390), .B2(new_n391), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT6), .ZN(new_n490));
  NOR3_X1   g0290(.A1(new_n490), .A2(new_n219), .A3(G107), .ZN(new_n491));
  XNOR2_X1  g0291(.A(G97), .B(G107), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n491), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  OAI22_X1  g0293(.A1(new_n493), .A2(new_n237), .B1(new_n210), .B2(new_n286), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n291), .B1(new_n489), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n474), .A2(G97), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n294), .A2(new_n219), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  AND2_X1   g0298(.A1(KEYINPUT5), .A2(G41), .ZN(new_n499));
  NOR2_X1   g0299(.A1(KEYINPUT5), .A2(G41), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n446), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OR2_X1    g0301(.A1(new_n501), .A2(new_n259), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n263), .A2(new_n501), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(new_n220), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n268), .A2(new_n270), .A3(G250), .A4(G1698), .ZN(new_n506));
  AND2_X1   g0306(.A1(KEYINPUT4), .A2(G244), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n268), .A2(new_n270), .A3(new_n507), .A4(new_n272), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G33), .A2(G283), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n506), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT4), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n376), .A2(G244), .A3(new_n272), .A4(new_n268), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n502), .B(new_n505), .C1(new_n513), .C2(new_n312), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G200), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n512), .A2(new_n511), .ZN(new_n516));
  INV_X1    g0316(.A(new_n510), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n279), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n519), .A2(G190), .A3(new_n502), .A4(new_n505), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n498), .A2(new_n515), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n514), .A2(new_n412), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n519), .A2(new_n281), .A3(new_n502), .A4(new_n505), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n267), .A2(G97), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n237), .A2(new_n509), .A3(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(G116), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n290), .A2(new_n238), .B1(G20), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT20), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n528), .A2(KEYINPUT20), .A3(new_n530), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n533), .A2(new_n534), .B1(new_n474), .B2(G116), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n294), .A2(new_n529), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n220), .A2(new_n272), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n223), .A2(G1698), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n376), .A2(new_n268), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n274), .A2(G303), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT84), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n540), .A2(KEYINPUT84), .A3(new_n541), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n544), .A2(new_n279), .A3(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n502), .ZN(new_n547));
  INV_X1    g0347(.A(new_n503), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n547), .B1(G270), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n537), .B1(new_n550), .B2(G190), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n304), .B2(new_n550), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT24), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT85), .ZN(new_n554));
  OAI21_X1  g0354(.A(KEYINPUT23), .B1(new_n234), .B2(G107), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT86), .ZN(new_n556));
  NOR2_X1   g0356(.A1(KEYINPUT23), .A2(G107), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n235), .A2(new_n236), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT86), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n559), .B(KEYINPUT23), .C1(new_n234), .C2(G107), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n234), .A2(G33), .A3(G116), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n556), .A2(new_n558), .A3(new_n560), .A4(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT22), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n271), .A2(G87), .A3(new_n237), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n380), .A2(KEYINPUT22), .A3(G87), .A4(new_n237), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n554), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n562), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n237), .A2(G87), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n563), .B1(new_n569), .B2(new_n274), .ZN(new_n570));
  AND4_X1   g0370(.A1(new_n554), .A2(new_n568), .A3(new_n570), .A4(new_n566), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n553), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n568), .A2(new_n570), .A3(new_n566), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT85), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n565), .A2(new_n554), .A3(new_n566), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n574), .A2(new_n575), .A3(KEYINPUT24), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n572), .A2(new_n291), .A3(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n503), .A2(new_n223), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n376), .B(new_n268), .C1(G257), .C2(new_n272), .ZN(new_n579));
  NOR2_X1   g0379(.A1(G250), .A2(G1698), .ZN(new_n580));
  INV_X1    g0380(.A(G294), .ZN(new_n581));
  OAI22_X1  g0381(.A1(new_n579), .A2(new_n580), .B1(new_n267), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n578), .B1(new_n582), .B2(new_n279), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n583), .A2(new_n502), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(G190), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT25), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n396), .B2(G107), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n587), .A2(KEYINPUT87), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n294), .A2(KEYINPUT25), .A3(new_n222), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n587), .A2(KEYINPUT87), .A3(new_n589), .ZN(new_n590));
  AOI211_X1 g0390(.A(new_n588), .B(new_n590), .C1(G107), .C2(new_n474), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n583), .A2(new_n502), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G200), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n577), .A2(new_n585), .A3(new_n591), .A4(new_n593), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n526), .A2(new_n552), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n550), .A2(G179), .A3(new_n537), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n412), .B1(new_n535), .B2(new_n536), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n546), .A2(new_n549), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT21), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n599), .B1(new_n597), .B2(new_n598), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n596), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n592), .A2(new_n412), .ZN(new_n603));
  INV_X1    g0403(.A(G179), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n577), .A2(new_n591), .B1(new_n604), .B2(new_n584), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n602), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT83), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n477), .A2(new_n486), .A3(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n488), .A2(new_n595), .A3(new_n606), .A4(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n435), .A2(new_n609), .ZN(G372));
  INV_X1    g0410(.A(new_n300), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n347), .A2(new_n348), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n612), .B1(new_n434), .B2(new_n343), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n419), .B1(new_n613), .B2(new_n430), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n306), .A2(new_n309), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n611), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n525), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n488), .A2(new_n619), .A3(new_n608), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(KEYINPUT26), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n473), .A2(new_n482), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n454), .A2(new_n412), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n479), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g0424(.A(new_n624), .B(KEYINPUT88), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n526), .A2(new_n594), .ZN(new_n626));
  INV_X1    g0426(.A(new_n537), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n627), .A2(new_n598), .A3(new_n604), .ZN(new_n628));
  INV_X1    g0428(.A(new_n601), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n597), .A2(new_n599), .A3(new_n598), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n577), .A2(new_n591), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n584), .A2(new_n604), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(new_n603), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n626), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n462), .B(new_n476), .C1(new_n304), .C2(new_n456), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n636), .A2(new_n624), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n625), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n636), .A2(new_n639), .A3(new_n619), .A4(new_n624), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n621), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n618), .B1(new_n435), .B2(new_n642), .ZN(G369));
  NAND2_X1  g0443(.A1(new_n237), .A2(G13), .ZN(new_n644));
  OR3_X1    g0444(.A1(new_n644), .A2(KEYINPUT27), .A3(G1), .ZN(new_n645));
  OAI21_X1  g0445(.A(KEYINPUT27), .B1(new_n644), .B2(G1), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(G213), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(G343), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n631), .A2(new_n537), .A3(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n649), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n602), .B1(new_n627), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n650), .A2(new_n552), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(G330), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n634), .A2(new_n649), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n594), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n651), .B1(new_n577), .B2(new_n591), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n634), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT89), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n631), .A2(new_n649), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n658), .B1(new_n662), .B2(new_n666), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n664), .A2(new_n667), .ZN(G399));
  AND3_X1   g0468(.A1(new_n477), .A2(new_n486), .A3(new_n607), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n607), .B1(new_n477), .B2(new_n486), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n671), .A2(new_n606), .A3(new_n595), .A4(new_n651), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n456), .A2(KEYINPUT90), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT90), .ZN(new_n674));
  AOI211_X1 g0474(.A(new_n674), .B(new_n452), .C1(new_n442), .C2(new_n279), .ZN(new_n675));
  INV_X1    g0475(.A(new_n514), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n673), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n677), .A2(new_n281), .A3(new_n598), .A4(new_n592), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT30), .ZN(new_n679));
  OAI21_X1  g0479(.A(G179), .B1(new_n460), .B2(new_n461), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n550), .A2(new_n583), .A3(new_n676), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n455), .A2(new_n458), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n583), .A2(new_n546), .A3(new_n549), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(new_n514), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n683), .A2(KEYINPUT30), .A3(new_n685), .A4(G179), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n678), .A2(new_n682), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n649), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT31), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT91), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AND3_X1   g0492(.A1(new_n687), .A2(KEYINPUT31), .A3(new_n649), .ZN(new_n693));
  AOI21_X1  g0493(.A(KEYINPUT31), .B1(new_n687), .B2(new_n649), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n672), .B(new_n692), .C1(new_n695), .C2(new_n691), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n488), .A2(new_n639), .A3(new_n619), .A4(new_n608), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT88), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n624), .B(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n636), .A2(new_n619), .A3(new_n624), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(KEYINPUT26), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n634), .A2(new_n631), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n526), .A2(new_n594), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n637), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n699), .A2(new_n701), .A3(new_n703), .A4(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n651), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT29), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT29), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n641), .A2(new_n710), .A3(new_n651), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n698), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n257), .ZN(new_n713));
  INV_X1    g0513(.A(new_n227), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G41), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n469), .A2(G116), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(G1), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n232), .B2(new_n716), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT28), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n713), .A2(new_n720), .ZN(G364));
  AOI21_X1  g0521(.A(new_n238), .B1(G20), .B2(new_n412), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n237), .A2(G190), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT96), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G179), .A2(G200), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n281), .A2(new_n237), .ZN(new_n728));
  INV_X1    g0528(.A(G190), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n728), .A2(new_n729), .A3(G200), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  XNOR2_X1  g0531(.A(KEYINPUT33), .B(G317), .ZN(new_n732));
  AOI22_X1  g0532(.A1(new_n727), .A2(G329), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(G311), .ZN(new_n734));
  XOR2_X1   g0534(.A(new_n728), .B(KEYINPUT94), .Z(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(new_n729), .A3(new_n304), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n733), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n304), .A2(G179), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT98), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n724), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g0540(.A(new_n740), .B(KEYINPUT99), .Z(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n737), .B1(new_n742), .B2(G283), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n739), .A2(G20), .A3(G190), .ZN(new_n744));
  INV_X1    g0544(.A(G303), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n274), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n728), .A2(G190), .A3(G200), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT95), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n747), .A2(new_n748), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n746), .B1(new_n751), .B2(G326), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n725), .A2(G190), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n358), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n743), .B(new_n752), .C1(new_n581), .C2(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n735), .A2(G190), .A3(new_n304), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n756), .B1(G322), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n736), .ZN(new_n760));
  INV_X1    g0560(.A(new_n744), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n760), .A2(G77), .B1(G87), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n727), .A2(G159), .ZN(new_n763));
  XOR2_X1   g0563(.A(KEYINPUT97), .B(KEYINPUT32), .Z(new_n764));
  OR2_X1    g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n274), .B1(new_n763), .B2(new_n764), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n755), .A2(new_n219), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n762), .A2(new_n765), .A3(new_n766), .A4(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n741), .A2(new_n222), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n757), .A2(new_n217), .ZN(new_n771));
  INV_X1    g0571(.A(new_n751), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n772), .A2(new_n292), .B1(new_n208), .B2(new_n730), .ZN(new_n773));
  NOR4_X1   g0573(.A1(new_n769), .A2(new_n770), .A3(new_n771), .A4(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n722), .B1(new_n759), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n227), .A2(G355), .A3(new_n271), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n714), .A2(new_n380), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(G45), .B2(new_n232), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n252), .A2(new_n445), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n776), .B1(G116), .B2(new_n227), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G13), .A2(G33), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(G20), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT93), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n722), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n780), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n644), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n257), .B1(new_n788), .B2(G45), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n716), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT92), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n784), .B(KEYINPUT100), .Z(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n653), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n775), .A2(new_n787), .A3(new_n791), .A4(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n791), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n653), .A2(new_n654), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n656), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n795), .A2(new_n798), .ZN(G396));
  NAND2_X1  g0599(.A1(new_n742), .A2(G87), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n800), .B1(new_n529), .B2(new_n736), .C1(new_n745), .C2(new_n772), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(G107), .B2(new_n761), .ZN(new_n802));
  INV_X1    g0602(.A(G283), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n274), .B1(new_n730), .B2(new_n803), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n767), .B(new_n804), .C1(new_n727), .C2(G311), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n802), .B(new_n805), .C1(new_n581), .C2(new_n757), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT101), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n751), .A2(G137), .B1(G150), .B2(new_n731), .ZN(new_n808));
  INV_X1    g0608(.A(G143), .ZN(new_n809));
  INV_X1    g0609(.A(G159), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n808), .B1(new_n809), .B2(new_n757), .C1(new_n810), .C2(new_n736), .ZN(new_n811));
  XOR2_X1   g0611(.A(KEYINPUT102), .B(KEYINPUT34), .Z(new_n812));
  XNOR2_X1  g0612(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n741), .A2(new_n208), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n727), .A2(G132), .B1(G58), .B2(new_n754), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n292), .B2(new_n744), .ZN(new_n816));
  NOR4_X1   g0616(.A1(new_n813), .A2(new_n377), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n722), .B1(new_n807), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n818), .A2(new_n791), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n722), .A2(new_n781), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NOR3_X1   g0621(.A1(new_n431), .A2(new_n433), .A3(new_n649), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n368), .A2(new_n370), .B1(new_n367), .B2(new_n651), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n822), .B1(new_n823), .B2(new_n434), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n819), .B1(G77), .B2(new_n821), .C1(new_n782), .C2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n824), .B1(new_n641), .B2(new_n651), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n639), .B1(new_n671), .B2(new_n619), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n706), .A2(new_n640), .A3(new_n701), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n651), .B(new_n824), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT103), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n641), .A2(KEYINPUT103), .A3(new_n651), .A4(new_n824), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n826), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(new_n698), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(new_n796), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n825), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(G384));
  NAND4_X1  g0637(.A1(new_n416), .A2(new_n426), .A3(new_n428), .A4(new_n418), .ZN(new_n838));
  INV_X1    g0638(.A(new_n647), .ZN(new_n839));
  INV_X1    g0639(.A(new_n398), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n388), .A2(new_n291), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n382), .A2(new_n387), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n389), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n840), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n838), .A2(new_n839), .A3(new_n845), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n422), .A2(new_n395), .A3(new_n398), .A4(new_n424), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n839), .B1(new_n413), .B2(new_n414), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n847), .B1(new_n848), .B2(new_n844), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(KEYINPUT37), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT37), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n851), .B(new_n847), .C1(new_n848), .C2(new_n427), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  AND3_X1   g0653(.A1(new_n846), .A2(KEYINPUT38), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT38), .B1(new_n846), .B2(new_n853), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(KEYINPUT39), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT38), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n847), .B1(new_n848), .B2(new_n427), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT37), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT104), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n860), .A2(new_n861), .A3(new_n852), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n838), .A2(new_n399), .A3(new_n839), .ZN(new_n863));
  OR2_X1    g0663(.A1(new_n848), .A2(new_n427), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n864), .A2(KEYINPUT104), .A3(new_n851), .A4(new_n847), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n862), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n854), .B1(new_n858), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n857), .B1(KEYINPUT39), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n343), .A2(new_n649), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  OAI22_X1  g0670(.A1(new_n868), .A2(new_n870), .B1(new_n420), .B2(new_n839), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n822), .B1(new_n831), .B2(new_n832), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n342), .A2(new_n649), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n343), .A2(new_n349), .A3(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n342), .B(new_n649), .C1(new_n612), .C2(new_n330), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n872), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n856), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n871), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n435), .B1(new_n709), .B2(new_n711), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n881), .A2(new_n617), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n880), .B(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT40), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n876), .A2(new_n824), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n609), .A2(new_n649), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n687), .A2(KEYINPUT31), .A3(new_n649), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n690), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n885), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n884), .B1(new_n889), .B2(new_n856), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n866), .A2(new_n858), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n846), .A2(new_n853), .A3(KEYINPUT38), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n876), .A2(new_n824), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(new_n695), .B2(new_n672), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n893), .A2(new_n895), .A3(KEYINPUT40), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n890), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n886), .A2(new_n888), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n435), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n897), .B(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n900), .A2(new_n654), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n883), .B(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n257), .B2(new_n788), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT35), .ZN(new_n904));
  AOI211_X1 g0704(.A(new_n238), .B(new_n237), .C1(new_n493), .C2(new_n904), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n905), .B(G116), .C1(new_n904), .C2(new_n493), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n906), .B(KEYINPUT36), .ZN(new_n907));
  OAI21_X1  g0707(.A(G77), .B1(new_n217), .B2(new_n208), .ZN(new_n908));
  OAI22_X1  g0708(.A1(new_n232), .A2(new_n908), .B1(G50), .B2(new_n208), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(G1), .A3(new_n293), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n903), .A2(new_n907), .A3(new_n910), .ZN(G367));
  XNOR2_X1  g0711(.A(new_n715), .B(KEYINPUT41), .ZN(new_n912));
  INV_X1    g0712(.A(new_n667), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n526), .B1(new_n498), .B2(new_n651), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n619), .A2(new_n649), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT45), .ZN(new_n918));
  OR3_X1    g0718(.A1(new_n913), .A2(KEYINPUT44), .A3(new_n916), .ZN(new_n919));
  OAI21_X1  g0719(.A(KEYINPUT44), .B1(new_n913), .B2(new_n916), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(new_n664), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n662), .B(new_n666), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(new_n656), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n712), .A2(new_n925), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n912), .B1(new_n927), .B2(new_n712), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n789), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n662), .A2(new_n666), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n916), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT42), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n930), .A2(KEYINPUT42), .A3(new_n916), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n525), .B1(new_n914), .B2(new_n634), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n933), .A2(new_n934), .B1(new_n651), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n476), .A2(new_n651), .ZN(new_n937));
  MUX2_X1   g0737(.A(new_n637), .B(new_n625), .S(new_n937), .Z(new_n938));
  NOR2_X1   g0738(.A1(new_n938), .A2(KEYINPUT43), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT105), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n940), .B(new_n941), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n938), .A2(KEYINPUT43), .ZN(new_n943));
  OR3_X1    g0743(.A1(new_n936), .A2(new_n939), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n945), .A2(KEYINPUT106), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(KEYINPUT106), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n946), .A2(new_n664), .A3(new_n916), .A4(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n946), .A2(new_n947), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n664), .A2(new_n916), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n929), .A2(new_n948), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n757), .A2(new_n284), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n760), .A2(G50), .B1(G159), .B2(new_n731), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n208), .B2(new_n755), .ZN(new_n955));
  AOI211_X1 g0755(.A(new_n953), .B(new_n955), .C1(G143), .C2(new_n751), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n761), .A2(G58), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n727), .A2(G137), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n274), .B1(new_n740), .B2(G77), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n956), .A2(new_n957), .A3(new_n958), .A4(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n772), .A2(new_n734), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n757), .A2(new_n745), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n736), .A2(new_n803), .B1(new_n222), .B2(new_n755), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n962), .B(new_n963), .C1(G317), .C2(new_n727), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT46), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n744), .B2(new_n529), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n740), .A2(G97), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n744), .A2(new_n965), .A3(new_n529), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n380), .B(new_n968), .C1(G294), .C2(new_n731), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n964), .A2(new_n966), .A3(new_n967), .A4(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n960), .B1(new_n961), .B2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT47), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n722), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n938), .A2(new_n792), .ZN(new_n974));
  INV_X1    g0774(.A(new_n777), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n786), .B1(new_n227), .B2(new_n361), .C1(new_n248), .C2(new_n975), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n973), .A2(new_n791), .A3(new_n974), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n952), .A2(new_n977), .ZN(G387));
  AND2_X1   g0778(.A1(new_n245), .A2(G45), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n227), .A2(new_n271), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n979), .A2(new_n975), .B1(new_n717), .B2(new_n980), .ZN(new_n981));
  OR3_X1    g0781(.A1(new_n288), .A2(KEYINPUT50), .A3(G50), .ZN(new_n982));
  AOI21_X1  g0782(.A(G45), .B1(G68), .B2(G77), .ZN(new_n983));
  OAI21_X1  g0783(.A(KEYINPUT50), .B1(new_n288), .B2(G50), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n982), .A2(new_n717), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n981), .A2(new_n985), .B1(new_n222), .B2(new_n714), .ZN(new_n986));
  INV_X1    g0786(.A(new_n786), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n791), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n722), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n751), .A2(G322), .B1(G311), .B2(new_n731), .ZN(new_n990));
  INV_X1    g0790(.A(G317), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n990), .B1(new_n745), .B2(new_n736), .C1(new_n991), .C2(new_n757), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT48), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n993), .B1(new_n803), .B2(new_n755), .C1(new_n581), .C2(new_n744), .ZN(new_n994));
  XOR2_X1   g0794(.A(KEYINPUT107), .B(KEYINPUT49), .Z(new_n995));
  XNOR2_X1  g0795(.A(new_n994), .B(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n740), .A2(G116), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n380), .B1(new_n727), .B2(G326), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n380), .B1(new_n757), .B2(new_n292), .C1(new_n208), .C2(new_n736), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n730), .A2(new_n288), .B1(new_n361), .B2(new_n755), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n744), .A2(new_n210), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n726), .A2(new_n284), .ZN(new_n1003));
  NOR4_X1   g0803(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n219), .B2(new_n741), .C1(new_n810), .C2(new_n772), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n989), .B1(new_n999), .B2(new_n1005), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n988), .B(new_n1006), .C1(new_n662), .C2(new_n793), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n789), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n925), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n712), .A2(new_n925), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n715), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1010), .B1(new_n926), .B2(new_n1012), .ZN(G393));
  OAI221_X1 g0813(.A(new_n786), .B1(new_n219), .B2(new_n227), .C1(new_n975), .C2(new_n255), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n791), .B(new_n1014), .C1(new_n916), .C2(new_n784), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n760), .A2(G294), .B1(G116), .B2(new_n754), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n745), .B2(new_n730), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT108), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1018), .A2(new_n770), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n727), .A2(G322), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n772), .A2(new_n991), .B1(new_n757), .B2(new_n734), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT52), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n271), .B1(new_n761), .B2(G283), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1019), .A2(new_n1020), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n758), .A2(G159), .B1(G150), .B2(new_n751), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT51), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n377), .B(new_n1026), .C1(new_n357), .C2(new_n760), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n754), .A2(G77), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n761), .A2(G68), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n727), .A2(G143), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n800), .B1(new_n292), .B2(new_n730), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1024), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT109), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1015), .B1(new_n1034), .B2(new_n722), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n923), .B2(new_n1008), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n715), .B1(new_n923), .B2(new_n926), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1036), .B1(new_n927), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT110), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(G390));
  NAND2_X1  g0842(.A1(new_n823), .A2(new_n434), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n707), .A2(new_n651), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n822), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n696), .A2(G330), .A3(new_n824), .A4(new_n876), .ZN(new_n1047));
  OAI211_X1 g0847(.A(G330), .B(new_n824), .C1(new_n886), .C2(new_n888), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n877), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1046), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n609), .A2(new_n649), .B1(new_n694), .B2(KEYINPUT91), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n691), .B1(new_n690), .B2(new_n887), .ZN(new_n1052));
  OAI211_X1 g0852(.A(G330), .B(new_n824), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n654), .B1(new_n695), .B2(new_n672), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n1053), .A2(new_n877), .B1(new_n885), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1050), .B1(new_n872), .B2(new_n1055), .ZN(new_n1056));
  NOR3_X1   g0856(.A1(new_n435), .A2(new_n898), .A3(new_n654), .ZN(new_n1057));
  NOR3_X1   g0857(.A1(new_n881), .A2(new_n1057), .A3(new_n617), .ZN(new_n1058));
  AND3_X1   g0858(.A1(new_n1056), .A2(KEYINPUT112), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(KEYINPUT112), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n870), .B1(new_n872), .B2(new_n877), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n868), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n867), .A2(new_n869), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1064), .B(KEYINPUT111), .C1(new_n1046), .C2(new_n877), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT111), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n877), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n893), .A2(new_n870), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1065), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1047), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1063), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n1062), .A2(new_n868), .B1(new_n1069), .B2(new_n1065), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1054), .A2(new_n885), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1072), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n716), .B1(new_n1061), .B2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n1076), .B2(new_n1061), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1076), .A2(new_n1008), .ZN(new_n1079));
  XOR2_X1   g0879(.A(KEYINPUT54), .B(G143), .Z(new_n1080));
  AOI22_X1  g0880(.A1(new_n760), .A2(new_n1080), .B1(G159), .B2(new_n754), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n740), .A2(G50), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n758), .A2(G132), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G125), .B2(new_n727), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n751), .A2(G128), .ZN(new_n1086));
  OAI21_X1  g0886(.A(KEYINPUT53), .B1(new_n744), .B2(new_n284), .ZN(new_n1087));
  NOR3_X1   g0887(.A1(new_n744), .A2(KEYINPUT53), .A3(new_n284), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n274), .B(new_n1088), .C1(G137), .C2(new_n731), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .A4(new_n1089), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n751), .A2(G283), .B1(G107), .B2(new_n731), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n219), .B2(new_n736), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT113), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n274), .B(new_n1028), .C1(new_n757), .C2(new_n529), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(G294), .B2(new_n727), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1093), .B(new_n1095), .C1(new_n468), .C2(new_n744), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1090), .B1(new_n1096), .B2(new_n814), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT114), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n791), .B1(new_n357), .B2(new_n821), .C1(new_n1098), .C2(new_n989), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n1099), .A2(KEYINPUT115), .B1(new_n781), .B2(new_n868), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(KEYINPUT115), .B2(new_n1099), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1078), .A2(new_n1079), .A3(new_n1101), .ZN(G378));
  INV_X1    g0902(.A(KEYINPUT122), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n890), .A2(new_n896), .A3(G330), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT120), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n890), .A2(new_n896), .A3(KEYINPUT120), .A4(G330), .ZN(new_n1107));
  XOR2_X1   g0907(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n310), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n310), .A2(new_n1109), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n298), .A2(new_n839), .ZN(new_n1112));
  OR3_X1    g0912(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1112), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1106), .A2(new_n1107), .A3(new_n1116), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n897), .A2(KEYINPUT120), .A3(G330), .A4(new_n1115), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n878), .A2(new_n879), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n871), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n880), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1123), .A2(KEYINPUT57), .A3(new_n1124), .ZN(new_n1125));
  AOI221_X4 g0925(.A(new_n1047), .B1(new_n1065), .B2(new_n1069), .C1(new_n1062), .C2(new_n868), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1075), .B1(new_n1063), .B2(new_n1070), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n1126), .A2(new_n1127), .B1(new_n1060), .B2(new_n1059), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1125), .B1(new_n1058), .B2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1103), .B1(new_n1129), .B2(new_n716), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT57), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1058), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n1061), .B2(new_n1076), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT121), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1117), .A2(new_n1134), .A3(new_n1118), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(new_n1122), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1131), .B1(new_n1133), .B2(new_n1136), .ZN(new_n1137));
  OAI211_X1 g0937(.A(KEYINPUT122), .B(new_n715), .C1(new_n1133), .C2(new_n1125), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1130), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1136), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n1008), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n736), .A2(new_n361), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n740), .A2(G58), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT116), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n1002), .A2(G41), .A3(new_n380), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1144), .B(new_n1145), .C1(new_n803), .C2(new_n726), .ZN(new_n1146));
  XOR2_X1   g0946(.A(new_n1146), .B(KEYINPUT117), .Z(new_n1147));
  AOI211_X1 g0947(.A(new_n1142), .B(new_n1147), .C1(G97), .C2(new_n731), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n751), .A2(G116), .B1(G68), .B2(new_n754), .ZN(new_n1149));
  XOR2_X1   g0949(.A(new_n1149), .B(KEYINPUT118), .Z(new_n1150));
  OAI211_X1 g0950(.A(new_n1148), .B(new_n1150), .C1(new_n222), .C2(new_n757), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT58), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n758), .A2(G128), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n760), .A2(G137), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n751), .A2(G125), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n761), .A2(new_n1080), .B1(G150), .B2(new_n754), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(G132), .B2(new_n731), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT59), .ZN(new_n1159));
  AOI21_X1  g0959(.A(G33), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n740), .A2(G159), .ZN(new_n1161));
  AOI21_X1  g0961(.A(G41), .B1(new_n727), .B2(G124), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1164));
  AOI21_X1  g0964(.A(G41), .B1(new_n376), .B2(G33), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n1163), .A2(new_n1164), .B1(G50), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n989), .B1(new_n1152), .B2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1116), .A2(new_n782), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n791), .B1(G50), .B2(new_n821), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT119), .ZN(new_n1171));
  OR3_X1    g0971(.A1(new_n1168), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n1141), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1139), .A2(new_n1173), .ZN(G375));
  NAND2_X1  g0974(.A1(new_n1144), .A2(new_n380), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1175), .A2(KEYINPUT123), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1175), .A2(KEYINPUT123), .B1(G137), .B2(new_n758), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n760), .A2(G150), .B1(new_n731), .B2(new_n1080), .ZN(new_n1178));
  INV_X1    g0978(.A(G128), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1178), .B1(new_n1179), .B2(new_n726), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(G50), .B2(new_n754), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1177), .B(new_n1181), .C1(new_n810), .C2(new_n744), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1176), .B(new_n1182), .C1(G132), .C2(new_n751), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n274), .B1(new_n529), .B2(new_n730), .C1(new_n741), .C2(new_n210), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(G294), .B2(new_n751), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n803), .B2(new_n757), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n744), .A2(new_n219), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n726), .A2(new_n745), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n736), .A2(new_n222), .B1(new_n361), .B2(new_n755), .ZN(new_n1189));
  NOR4_X1   g0989(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n722), .B1(new_n1183), .B2(new_n1190), .ZN(new_n1191));
  AND2_X1   g0991(.A1(new_n1191), .A2(new_n791), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1192), .B1(G68), .B2(new_n821), .C1(new_n782), .C2(new_n876), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n1056), .B2(new_n1008), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1196));
  OR2_X1    g0996(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n912), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1195), .B1(new_n1198), .B2(new_n1199), .ZN(G381));
  XNOR2_X1  g1000(.A(G375), .B(KEYINPUT124), .ZN(new_n1201));
  INV_X1    g1001(.A(G378), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n952), .A2(new_n977), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1203));
  NOR4_X1   g1003(.A1(new_n1203), .A2(G396), .A3(G393), .A4(G381), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1201), .A2(new_n836), .A3(new_n1202), .A4(new_n1204), .ZN(G407));
  NAND3_X1  g1005(.A1(new_n1201), .A2(new_n648), .A3(new_n1202), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(G407), .A2(G213), .A3(new_n1206), .ZN(G409));
  XOR2_X1   g1007(.A(G393), .B(G396), .Z(new_n1208));
  INV_X1    g1008(.A(new_n1203), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n952), .A2(new_n977), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1208), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1210), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1208), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1212), .A2(new_n1203), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1211), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(G213), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1216), .A2(G343), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1139), .A2(G378), .A3(new_n1173), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1133), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1219), .A2(new_n912), .A3(new_n1140), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1123), .A2(new_n1008), .A3(new_n1124), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1220), .A2(new_n1172), .A3(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1202), .A2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1217), .B1(new_n1218), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1198), .A2(KEYINPUT60), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT60), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1197), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1225), .A2(new_n715), .A3(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n1195), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(new_n836), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1228), .A2(G384), .A3(new_n1195), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT63), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1215), .B1(new_n1224), .B2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT61), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1218), .A2(new_n1223), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT125), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1217), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1218), .A2(KEYINPUT125), .A3(new_n1223), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1217), .A2(G2897), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1232), .A2(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1232), .A2(new_n1243), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1233), .B1(new_n1242), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1232), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1239), .A2(new_n1240), .A3(new_n1249), .A4(new_n1241), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1235), .B(new_n1236), .C1(new_n1248), .C2(new_n1251), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1211), .A2(new_n1214), .A3(KEYINPUT126), .ZN(new_n1253));
  AOI21_X1  g1053(.A(KEYINPUT126), .B1(new_n1211), .B2(new_n1214), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT62), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1232), .A2(new_n1256), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1224), .A2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(new_n1250), .B2(new_n1256), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1236), .B1(new_n1246), .B2(new_n1224), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1255), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1252), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT127), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1252), .A2(new_n1261), .A3(KEYINPUT127), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(G405));
  NAND2_X1  g1066(.A1(G375), .A2(new_n1202), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1218), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(new_n1268), .B(new_n1249), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(new_n1255), .B(new_n1269), .ZN(G402));
endmodule


