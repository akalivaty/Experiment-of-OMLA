//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1 0 0 1 0 0 0 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1204, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  AND2_X1   g0010(.A1(G116), .A2(G270), .ZN(new_n211));
  AND2_X1   g0011(.A1(KEYINPUT64), .A2(G68), .ZN(new_n212));
  NOR2_X1   g0012(.A1(KEYINPUT64), .A2(G68), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(new_n214), .A2(G238), .B1(G50), .B2(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  INV_X1    g0017(.A(G77), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI211_X1 g0020(.A(new_n211), .B(new_n220), .C1(G107), .C2(G264), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT65), .ZN(new_n223));
  AOI22_X1  g0023(.A1(new_n221), .A2(new_n223), .B1(G1), .B2(G20), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT1), .Z(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n207), .ZN(new_n227));
  INV_X1    g0027(.A(new_n201), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n210), .B(new_n225), .C1(new_n227), .C2(new_n230), .ZN(G361));
  XOR2_X1   g0031(.A(G226), .B(G232), .Z(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G58), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  AND2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  OAI211_X1 g0050(.A(G250), .B(new_n248), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  OAI211_X1 g0051(.A(G257), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G294), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n251), .B(new_n252), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G45), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G1), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT5), .B(G41), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n256), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G264), .ZN(new_n262));
  AND2_X1   g0062(.A1(new_n260), .A2(new_n259), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G274), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n257), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G179), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n255), .A2(new_n256), .B1(new_n261), .B2(G264), .ZN(new_n267));
  AOI21_X1  g0067(.A(G169), .B1(new_n267), .B2(new_n264), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n207), .B(G87), .C1(new_n249), .C2(new_n250), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT81), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(KEYINPUT22), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT23), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n273), .B1(new_n207), .B2(G107), .ZN(new_n274));
  INV_X1    g0074(.A(G107), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(KEYINPUT23), .A3(G20), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n270), .A2(new_n272), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  OR2_X1    g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT81), .B(KEYINPUT22), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n280), .A2(new_n281), .A3(new_n207), .A4(G87), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n277), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT24), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n226), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n277), .A2(KEYINPUT24), .A3(new_n282), .A4(new_n283), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n286), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n288), .B(KEYINPUT67), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n207), .A2(G1), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n292), .A2(G13), .B1(new_n206), .B2(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G107), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n292), .A2(G13), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(G107), .ZN(new_n298));
  XNOR2_X1  g0098(.A(KEYINPUT82), .B(KEYINPUT25), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n298), .B(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n290), .A2(new_n296), .A3(new_n300), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n269), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(G200), .B1(new_n267), .B2(new_n264), .ZN(new_n303));
  INV_X1    g0103(.A(G190), .ZN(new_n304));
  INV_X1    g0104(.A(new_n265), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n306), .A2(new_n301), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT83), .B1(new_n302), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G200), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n265), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(G190), .B2(new_n265), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n311), .A2(new_n296), .A3(new_n290), .A4(new_n300), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT83), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n269), .A2(new_n301), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n308), .A2(new_n315), .ZN(new_n316));
  XOR2_X1   g0116(.A(new_n288), .B(KEYINPUT67), .Z(new_n317));
  NOR2_X1   g0117(.A1(new_n317), .A2(new_n292), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n203), .A2(G20), .ZN(new_n319));
  INV_X1    g0119(.A(G150), .ZN(new_n320));
  NOR2_X1   g0120(.A1(G20), .A2(G33), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(KEYINPUT68), .A2(G58), .ZN(new_n323));
  XOR2_X1   g0123(.A(new_n323), .B(KEYINPUT8), .Z(new_n324));
  NAND2_X1  g0124(.A1(new_n207), .A2(G33), .ZN(new_n325));
  OAI221_X1 g0125(.A(new_n319), .B1(new_n320), .B2(new_n322), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n318), .A2(G50), .B1(new_n326), .B2(new_n317), .ZN(new_n327));
  INV_X1    g0127(.A(new_n297), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n202), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n331));
  INV_X1    g0131(.A(G274), .ZN(new_n332));
  OR2_X1    g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G226), .ZN(new_n334));
  INV_X1    g0134(.A(G41), .ZN(new_n335));
  OAI211_X1 g0135(.A(G1), .B(G13), .C1(new_n253), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n331), .ZN(new_n337));
  MUX2_X1   g0137(.A(G222), .B(G223), .S(G1698), .Z(new_n338));
  NOR2_X1   g0138(.A1(new_n249), .A2(new_n250), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n256), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n280), .A2(G77), .ZN(new_n341));
  OAI221_X1 g0141(.A(new_n333), .B1(new_n334), .B2(new_n337), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  OR2_X1    g0142(.A1(new_n342), .A2(G179), .ZN(new_n343));
  INV_X1    g0143(.A(G169), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n330), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n342), .A2(new_n304), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n348), .B1(G200), .B2(new_n342), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n327), .B(new_n329), .C1(KEYINPUT69), .C2(KEYINPUT9), .ZN(new_n350));
  AND2_X1   g0150(.A1(KEYINPUT69), .A2(KEYINPUT9), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n350), .A2(new_n351), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n349), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT10), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT10), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n356), .B(new_n349), .C1(new_n352), .C2(new_n353), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n347), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  XOR2_X1   g0158(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n359));
  OAI211_X1 g0159(.A(G226), .B(new_n248), .C1(new_n249), .C2(new_n250), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n360), .B(KEYINPUT70), .ZN(new_n361));
  OAI211_X1 g0161(.A(G232), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n362));
  NAND2_X1  g0162(.A1(G33), .A2(G97), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n336), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n336), .A2(G238), .A3(new_n331), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n367), .A2(new_n333), .A3(KEYINPUT71), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(KEYINPUT71), .B1(new_n367), .B2(new_n333), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n359), .B1(new_n366), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n367), .A2(new_n333), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT71), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n368), .ZN(new_n376));
  INV_X1    g0176(.A(new_n359), .ZN(new_n377));
  OR2_X1    g0177(.A1(new_n360), .A2(KEYINPUT70), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n360), .A2(KEYINPUT70), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n364), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n376), .B(new_n377), .C1(new_n380), .C2(new_n336), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n372), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G169), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT14), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT73), .B1(new_n366), .B2(new_n371), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT73), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n376), .B(new_n386), .C1(new_n380), .C2(new_n336), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n385), .A2(KEYINPUT13), .A3(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n388), .A2(G179), .A3(new_n381), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT14), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n382), .A2(new_n390), .A3(G169), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n384), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n321), .A2(G50), .ZN(new_n393));
  OAI221_X1 g0193(.A(new_n393), .B1(new_n218), .B2(new_n325), .C1(new_n214), .C2(new_n207), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n317), .A2(new_n394), .ZN(new_n395));
  XOR2_X1   g0195(.A(new_n395), .B(KEYINPUT11), .Z(new_n396));
  NOR2_X1   g0196(.A1(new_n288), .A2(new_n292), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT12), .ZN(new_n398));
  OAI21_X1  g0198(.A(G68), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n214), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n328), .A2(new_n400), .A3(KEYINPUT12), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n399), .B(new_n401), .C1(KEYINPUT12), .C2(new_n328), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n396), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n392), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n388), .A2(G190), .A3(new_n381), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n382), .A2(G200), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n406), .A2(new_n407), .A3(new_n403), .ZN(new_n408));
  AND2_X1   g0208(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  XOR2_X1   g0209(.A(KEYINPUT8), .B(G58), .Z(new_n410));
  AOI22_X1  g0210(.A1(new_n410), .A2(new_n321), .B1(G20), .B2(G77), .ZN(new_n411));
  XOR2_X1   g0211(.A(KEYINPUT15), .B(G87), .Z(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n411), .B1(new_n413), .B2(new_n325), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(new_n288), .B1(G77), .B2(new_n397), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(G77), .B2(new_n297), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n280), .A2(G238), .A3(G1698), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n280), .A2(G232), .A3(new_n248), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n417), .B(new_n418), .C1(new_n275), .C2(new_n280), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n256), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n336), .A2(new_n331), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(G244), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n420), .A2(new_n333), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n416), .B1(G200), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n423), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(G190), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n358), .A2(new_n409), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n324), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n429), .A2(new_n328), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n291), .B1(G1), .B2(new_n207), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n430), .B1(new_n431), .B2(new_n429), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT74), .ZN(new_n434));
  OR2_X1    g0234(.A1(KEYINPUT64), .A2(G68), .ZN(new_n435));
  NAND2_X1  g0235(.A1(KEYINPUT64), .A2(G68), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(G58), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n207), .B1(new_n437), .B2(new_n228), .ZN(new_n438));
  INV_X1    g0238(.A(G159), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n322), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n434), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n440), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n201), .B1(new_n214), .B2(G58), .ZN(new_n443));
  OAI211_X1 g0243(.A(KEYINPUT74), .B(new_n442), .C1(new_n443), .C2(new_n207), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n278), .A2(new_n207), .A3(new_n279), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT7), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n278), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n279), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(KEYINPUT75), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT75), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n446), .A2(new_n451), .A3(new_n447), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n450), .A2(new_n214), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT16), .B1(new_n445), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT7), .B1(new_n339), .B2(new_n207), .ZN(new_n455));
  INV_X1    g0255(.A(new_n449), .ZN(new_n456));
  OAI21_X1  g0256(.A(G68), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n441), .A2(new_n444), .A3(KEYINPUT16), .A4(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n288), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n433), .B1(new_n454), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n334), .A2(G1698), .ZN(new_n461));
  OAI221_X1 g0261(.A(new_n461), .B1(G223), .B2(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G33), .A2(G87), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n336), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n333), .B1(new_n337), .B2(new_n217), .ZN(new_n465));
  INV_X1    g0265(.A(G179), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n462), .A2(new_n463), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n256), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n331), .A2(new_n332), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n470), .B1(new_n421), .B2(G232), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n467), .B1(G169), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n460), .A2(KEYINPUT18), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(KEYINPUT18), .B1(new_n460), .B2(new_n474), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n458), .A2(new_n288), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n453), .A2(new_n441), .A3(new_n444), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT16), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(G200), .B1(new_n469), .B2(new_n471), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n464), .A2(new_n465), .A3(G190), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n483), .A2(new_n433), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT17), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n483), .A2(KEYINPUT17), .A3(new_n433), .A4(new_n487), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n425), .A2(new_n466), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n492), .B(new_n416), .C1(G169), .C2(new_n425), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n478), .A2(new_n490), .A3(new_n491), .A4(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n428), .A2(new_n494), .ZN(new_n495));
  AND2_X1   g0295(.A1(G33), .A2(G283), .ZN(new_n496));
  OAI211_X1 g0296(.A(G244), .B(new_n248), .C1(new_n249), .C2(new_n250), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT4), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n280), .A2(KEYINPUT4), .A3(G244), .A4(new_n248), .ZN(new_n500));
  OAI211_X1 g0300(.A(G250), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT76), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT76), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n280), .A2(new_n503), .A3(G250), .A4(G1698), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n499), .A2(new_n500), .A3(new_n502), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n256), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n261), .A2(G257), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n506), .A2(new_n264), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G169), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n505), .A2(new_n256), .B1(G257), .B2(new_n261), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(G179), .A3(new_n264), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT78), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n297), .A2(G97), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n450), .A2(G107), .A3(new_n452), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n275), .A2(KEYINPUT6), .A3(G97), .ZN(new_n516));
  XOR2_X1   g0316(.A(G97), .B(G107), .Z(new_n517));
  OAI21_X1  g0317(.A(new_n516), .B1(new_n517), .B2(KEYINPUT6), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n518), .A2(G20), .B1(G77), .B2(new_n321), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n514), .B1(new_n520), .B2(new_n288), .ZN(new_n521));
  INV_X1    g0321(.A(G97), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n294), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n513), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n515), .A2(new_n519), .B1(new_n226), .B2(new_n287), .ZN(new_n526));
  NOR4_X1   g0326(.A1(new_n526), .A2(KEYINPUT78), .A3(new_n523), .A4(new_n514), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n512), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n506), .A2(G190), .A3(new_n264), .A4(new_n507), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n521), .A2(new_n529), .A3(new_n524), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT77), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n508), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n510), .A2(KEYINPUT77), .A3(new_n264), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n532), .A2(G200), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n528), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT21), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n261), .A2(G270), .B1(new_n263), .B2(G274), .ZN(new_n538));
  OAI211_X1 g0338(.A(G264), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n539));
  OAI211_X1 g0339(.A(G257), .B(new_n248), .C1(new_n249), .C2(new_n250), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n278), .A2(G303), .A3(new_n279), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT79), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n542), .A2(new_n543), .A3(new_n256), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n543), .B1(new_n542), .B2(new_n256), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n538), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G169), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n293), .A2(G116), .ZN(new_n548));
  OAI22_X1  g0348(.A1(new_n548), .A2(new_n288), .B1(G116), .B2(new_n297), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n496), .A2(G20), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n550), .B1(G33), .B2(new_n522), .ZN(new_n551));
  INV_X1    g0351(.A(G116), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G20), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n288), .A2(KEYINPUT80), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(KEYINPUT80), .B1(new_n288), .B2(new_n553), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n551), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT20), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(KEYINPUT20), .B(new_n551), .C1(new_n554), .C2(new_n555), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n549), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n537), .B1(new_n547), .B2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n560), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n562), .A2(KEYINPUT21), .A3(G169), .A4(new_n546), .ZN(new_n563));
  OAI211_X1 g0363(.A(G179), .B(new_n538), .C1(new_n544), .C2(new_n545), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n562), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n561), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n546), .A2(G200), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n568), .B(new_n560), .C1(new_n304), .C2(new_n546), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(G238), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n248), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n219), .A2(G1698), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n572), .B(new_n573), .C1(new_n249), .C2(new_n250), .ZN(new_n574));
  NAND2_X1  g0374(.A1(G33), .A2(G116), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n576), .A2(new_n256), .B1(G274), .B2(new_n259), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n336), .B(G250), .C1(G1), .C2(new_n258), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n309), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT19), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n207), .B1(new_n363), .B2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(G87), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n582), .A2(new_n522), .A3(new_n275), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n207), .B(G68), .C1(new_n249), .C2(new_n250), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n580), .B1(new_n325), .B2(new_n522), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n587), .A2(new_n288), .B1(new_n328), .B2(new_n413), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n291), .A2(G87), .A3(new_n293), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n579), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n576), .A2(new_n256), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n259), .A2(G274), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n592), .A2(new_n593), .A3(new_n578), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(G190), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n291), .A2(new_n293), .A3(new_n412), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n594), .A2(new_n344), .B1(new_n588), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n577), .A2(new_n466), .A3(new_n578), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n591), .A2(new_n596), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NOR3_X1   g0401(.A1(new_n567), .A2(new_n570), .A3(new_n601), .ZN(new_n602));
  AND4_X1   g0402(.A1(new_n316), .A2(new_n495), .A3(new_n536), .A4(new_n602), .ZN(G372));
  INV_X1    g0403(.A(new_n405), .ZN(new_n604));
  INV_X1    g0404(.A(new_n493), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n408), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n490), .A2(new_n491), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n478), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n355), .A2(new_n357), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n347), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n495), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n598), .A2(new_n599), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n591), .A2(KEYINPUT84), .B1(G190), .B2(new_n595), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT84), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n579), .B2(new_n590), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n613), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  AND4_X1   g0417(.A1(new_n312), .A2(new_n528), .A3(new_n617), .A4(new_n535), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n567), .A2(KEYINPUT85), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT85), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n561), .A2(new_n563), .A3(new_n620), .A4(new_n566), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n619), .A2(new_n314), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n512), .B(new_n600), .C1(new_n525), .C2(new_n527), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(KEYINPUT26), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n614), .A2(new_n616), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n509), .A2(new_n511), .B1(new_n521), .B2(new_n524), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT26), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n626), .A2(new_n627), .A3(new_n628), .A4(new_n612), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n625), .A2(new_n612), .A3(new_n629), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n623), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n610), .B1(new_n611), .B2(new_n631), .ZN(G369));
  INV_X1    g0432(.A(G13), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n633), .A2(G20), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n206), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n635), .A2(KEYINPUT27), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(KEYINPUT27), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(G213), .A3(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(G343), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n560), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n643), .B1(new_n619), .B2(new_n621), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n567), .A2(new_n570), .A3(new_n642), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(G330), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n301), .A2(new_n640), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n316), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n269), .A2(new_n301), .A3(new_n640), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n651), .B(KEYINPUT86), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n314), .A2(new_n640), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n567), .A2(new_n641), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT87), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n656), .B(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n655), .B1(new_n653), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n654), .A2(new_n659), .ZN(G399));
  NAND2_X1  g0460(.A1(new_n208), .A2(new_n335), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n583), .A2(G116), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(new_n662), .A3(G1), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n229), .B2(new_n661), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n664), .B(KEYINPUT28), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT29), .ZN(new_n666));
  INV_X1    g0466(.A(new_n617), .ZN(new_n667));
  INV_X1    g0467(.A(new_n627), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT26), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n624), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n613), .B1(new_n670), .B2(new_n628), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n314), .A2(new_n561), .A3(new_n566), .A4(new_n563), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT88), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n528), .A2(new_n617), .A3(new_n535), .A4(new_n312), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n669), .B(new_n671), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n666), .B1(new_n676), .B2(new_n641), .ZN(new_n677));
  AOI211_X1 g0477(.A(KEYINPUT29), .B(new_n640), .C1(new_n623), .C2(new_n630), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n316), .A2(new_n536), .A3(new_n602), .A4(new_n641), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT30), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n261), .A2(G270), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n264), .ZN(new_n683));
  INV_X1    g0483(.A(new_n545), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n542), .A2(new_n543), .A3(new_n256), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n686), .A2(G179), .A3(new_n510), .A4(new_n595), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n681), .B1(new_n687), .B2(new_n265), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n686), .A2(new_n305), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n689), .A2(new_n466), .A3(new_n508), .A4(new_n594), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n510), .A2(new_n595), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n691), .A2(KEYINPUT30), .A3(new_n305), .A4(new_n565), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n688), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n640), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT31), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n693), .A2(KEYINPUT31), .A3(new_n640), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n680), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G330), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n679), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n665), .B1(new_n701), .B2(G1), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT89), .ZN(G364));
  NAND2_X1  g0503(.A1(new_n634), .A2(G45), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n661), .A2(G1), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n646), .ZN(new_n707));
  NOR2_X1   g0507(.A1(G13), .A2(G33), .ZN(new_n708));
  XOR2_X1   g0508(.A(new_n708), .B(KEYINPUT92), .Z(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(G20), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n707), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n243), .A2(G45), .ZN(new_n714));
  XOR2_X1   g0514(.A(new_n714), .B(KEYINPUT90), .Z(new_n715));
  NAND2_X1  g0515(.A1(new_n339), .A2(new_n208), .ZN(new_n716));
  XOR2_X1   g0516(.A(new_n716), .B(KEYINPUT91), .Z(new_n717));
  OAI211_X1 g0517(.A(new_n715), .B(new_n717), .C1(G45), .C2(new_n229), .ZN(new_n718));
  INV_X1    g0518(.A(G355), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n280), .A2(new_n208), .ZN(new_n720));
  OAI221_X1 g0520(.A(new_n718), .B1(G116), .B2(new_n208), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n226), .B1(G20), .B2(new_n344), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n711), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n207), .A2(G190), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(new_n466), .A3(new_n309), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n726), .A2(KEYINPUT93), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(KEYINPUT93), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n309), .A2(G179), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n725), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AOI22_X1  g0533(.A1(new_n730), .A2(G329), .B1(G283), .B2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(G326), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n207), .A2(new_n304), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n736), .A2(G179), .A3(G200), .ZN(new_n737));
  INV_X1    g0537(.A(new_n725), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n738), .A2(new_n466), .A3(new_n309), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  XOR2_X1   g0540(.A(KEYINPUT33), .B(G317), .Z(new_n741));
  OAI221_X1 g0541(.A(new_n734), .B1(new_n735), .B2(new_n737), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n466), .A2(new_n309), .ZN(new_n743));
  OAI21_X1  g0543(.A(G20), .B1(new_n743), .B2(new_n304), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT95), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n744), .A2(new_n745), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n254), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n736), .A2(new_n731), .ZN(new_n751));
  INV_X1    g0551(.A(G303), .ZN(new_n752));
  INV_X1    g0552(.A(G322), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n736), .A2(G179), .A3(new_n309), .ZN(new_n754));
  OAI221_X1 g0554(.A(new_n339), .B1(new_n751), .B2(new_n752), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n725), .A2(G179), .A3(new_n309), .ZN(new_n756));
  INV_X1    g0556(.A(G311), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR4_X1   g0558(.A1(new_n742), .A2(new_n750), .A3(new_n755), .A4(new_n758), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n748), .A2(G97), .B1(G68), .B2(new_n739), .ZN(new_n760));
  OAI221_X1 g0560(.A(new_n760), .B1(new_n218), .B2(new_n756), .C1(new_n275), .C2(new_n732), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n729), .A2(new_n439), .ZN(new_n762));
  XNOR2_X1  g0562(.A(KEYINPUT94), .B(KEYINPUT32), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n762), .B(new_n763), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n737), .A2(new_n202), .B1(new_n751), .B2(new_n582), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n280), .B1(new_n754), .B2(new_n216), .ZN(new_n766));
  NOR4_X1   g0566(.A1(new_n761), .A2(new_n764), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n722), .B1(new_n759), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n724), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n706), .B1(new_n713), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n707), .A2(G330), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n705), .B1(new_n771), .B2(new_n648), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT96), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(G396));
  INV_X1    g0575(.A(new_n699), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(KEYINPUT98), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n640), .B1(new_n623), .B2(new_n630), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n493), .A2(new_n640), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n424), .A2(new_n426), .B1(new_n416), .B2(new_n640), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n780), .B1(new_n605), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n778), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n777), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n776), .A2(KEYINPUT98), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n705), .B(new_n785), .C1(new_n787), .C2(new_n777), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n782), .A2(new_n709), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n730), .A2(G132), .B1(G68), .B2(new_n733), .ZN(new_n790));
  INV_X1    g0590(.A(new_n754), .ZN(new_n791));
  AOI22_X1  g0591(.A1(G150), .A2(new_n739), .B1(new_n791), .B2(G143), .ZN(new_n792));
  INV_X1    g0592(.A(G137), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n792), .B1(new_n793), .B2(new_n737), .C1(new_n439), .C2(new_n756), .ZN(new_n794));
  INV_X1    g0594(.A(KEYINPUT34), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n790), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n339), .B1(new_n794), .B2(new_n795), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(new_n202), .B2(new_n751), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n796), .B(new_n798), .C1(G58), .C2(new_n748), .ZN(new_n799));
  XOR2_X1   g0599(.A(KEYINPUT97), .B(G283), .Z(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n339), .B1(new_n254), .B2(new_n754), .C1(new_n740), .C2(new_n801), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n751), .A2(new_n275), .B1(new_n732), .B2(new_n582), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(new_n748), .B2(G97), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n804), .B1(new_n552), .B2(new_n756), .C1(new_n757), .C2(new_n729), .ZN(new_n805));
  INV_X1    g0605(.A(new_n737), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n802), .B(new_n805), .C1(G303), .C2(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n722), .B1(new_n799), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n722), .A2(new_n708), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n218), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n789), .A2(new_n808), .A3(new_n706), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n788), .A2(new_n811), .ZN(G384));
  XOR2_X1   g0612(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n813));
  INV_X1    g0613(.A(new_n638), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n460), .B(new_n814), .C1(new_n477), .C2(new_n607), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n483), .A2(new_n433), .B1(new_n473), .B2(new_n638), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n432), .B(new_n486), .C1(new_n479), .C2(new_n482), .ZN(new_n817));
  OAI21_X1  g0617(.A(KEYINPUT37), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n460), .B1(new_n474), .B2(new_n814), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT37), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n819), .A2(new_n820), .A3(new_n488), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n813), .B1(new_n815), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n441), .A2(new_n444), .A3(new_n457), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n481), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n826), .A2(new_n317), .A3(new_n458), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n638), .B1(new_n827), .B2(new_n433), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n477), .B2(new_n607), .ZN(new_n829));
  NOR3_X1   g0629(.A1(new_n816), .A2(new_n817), .A3(KEYINPUT37), .ZN(new_n830));
  AND3_X1   g0630(.A1(new_n826), .A2(new_n317), .A3(new_n458), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n831), .A2(new_n432), .B1(new_n474), .B2(new_n814), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n820), .B1(new_n832), .B2(new_n488), .ZN(new_n833));
  OAI21_X1  g0633(.A(KEYINPUT100), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n827), .A2(new_n433), .B1(new_n473), .B2(new_n638), .ZN(new_n835));
  OAI21_X1  g0635(.A(KEYINPUT37), .B1(new_n817), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT100), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n821), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n829), .A2(new_n834), .A3(KEYINPUT38), .A4(new_n838), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n839), .A2(KEYINPUT102), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n839), .A2(KEYINPUT102), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n824), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(KEYINPUT104), .B1(new_n694), .B2(new_n695), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT104), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n844), .B(KEYINPUT31), .C1(new_n693), .C2(new_n640), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n680), .B(new_n697), .C1(new_n843), .C2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n404), .A2(new_n640), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n405), .A2(new_n408), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n392), .A2(new_n404), .A3(new_n640), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n782), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n846), .A2(new_n850), .A3(KEYINPUT40), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n842), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n853), .A2(new_n495), .A3(new_n846), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT40), .ZN(new_n855));
  AND3_X1   g0655(.A1(new_n821), .A2(new_n836), .A3(new_n837), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n837), .B1(new_n821), .B2(new_n836), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT38), .B1(new_n858), .B2(new_n829), .ZN(new_n859));
  AND4_X1   g0659(.A1(KEYINPUT38), .A2(new_n829), .A3(new_n834), .A4(new_n838), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n850), .B(new_n846), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n854), .B1(new_n855), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n495), .A2(G330), .A3(new_n846), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n647), .B1(new_n861), .B2(new_n855), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n864), .B1(new_n865), .B2(new_n853), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n405), .A2(new_n640), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n829), .A2(new_n834), .A3(new_n838), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT38), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n871), .A2(KEYINPUT39), .A3(new_n839), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n839), .A2(KEYINPUT102), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT102), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n858), .A2(new_n874), .A3(KEYINPUT38), .A4(new_n829), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n823), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n868), .B(new_n872), .C1(new_n876), .C2(KEYINPUT39), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n779), .B1(new_n778), .B2(new_n783), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n848), .A2(new_n849), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT99), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n871), .A2(new_n839), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT99), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n640), .B(new_n782), .C1(new_n623), .C2(new_n630), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n883), .B(new_n879), .C1(new_n884), .C2(new_n779), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n881), .A2(new_n882), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n477), .A2(new_n638), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n877), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n867), .B(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n495), .B1(new_n677), .B2(new_n678), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n610), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n891), .B(KEYINPUT103), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n889), .B(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n206), .B2(new_n634), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n552), .B1(new_n518), .B2(KEYINPUT35), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n895), .B(new_n227), .C1(KEYINPUT35), .C2(new_n518), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n896), .B(KEYINPUT36), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n230), .A2(G77), .A3(new_n437), .ZN(new_n898));
  INV_X1    g0698(.A(G68), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n898), .B1(G50), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n900), .A2(G1), .A3(new_n633), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n894), .A2(new_n897), .A3(new_n901), .ZN(G367));
  NOR3_X1   g0702(.A1(new_n526), .A2(new_n514), .A3(new_n523), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n536), .B1(new_n903), .B2(new_n641), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n627), .A2(new_n640), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n906), .A2(new_n653), .A3(new_n658), .ZN(new_n907));
  INV_X1    g0707(.A(new_n528), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n907), .A2(KEYINPUT42), .B1(new_n908), .B2(new_n641), .ZN(new_n909));
  INV_X1    g0709(.A(new_n659), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT42), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n910), .B1(new_n911), .B2(new_n655), .ZN(new_n912));
  INV_X1    g0712(.A(new_n906), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n909), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n590), .A2(new_n640), .ZN(new_n915));
  OR2_X1    g0715(.A1(new_n667), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n613), .A2(new_n915), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g0718(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT106), .ZN(new_n921));
  INV_X1    g0721(.A(new_n918), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT43), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n914), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n654), .A2(new_n913), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n921), .B1(new_n914), .B2(new_n923), .ZN(new_n928));
  OR3_X1    g0728(.A1(new_n925), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n927), .B1(new_n925), .B2(new_n928), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n661), .B(KEYINPUT41), .Z(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n910), .A2(KEYINPUT44), .A3(new_n913), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT44), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n659), .B2(new_n906), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n659), .A2(new_n906), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT45), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n659), .A2(KEYINPUT45), .A3(new_n906), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n936), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n654), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n653), .A2(new_n658), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n653), .A2(new_n658), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n648), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n947), .A2(KEYINPUT107), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(KEYINPUT107), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n950), .A2(new_n946), .A3(new_n945), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n952), .A2(new_n700), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n936), .A2(new_n941), .A3(new_n654), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n944), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n932), .B1(new_n955), .B2(new_n701), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n704), .A2(G1), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n929), .B(new_n930), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n748), .A2(G68), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n959), .B1(new_n202), .B2(new_n756), .C1(new_n439), .C2(new_n740), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n339), .B(new_n960), .C1(G150), .C2(new_n791), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n730), .A2(G137), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n732), .A2(new_n218), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(G143), .B2(new_n806), .ZN(new_n964));
  INV_X1    g0764(.A(new_n751), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(G58), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n961), .A2(new_n962), .A3(new_n964), .A4(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(G317), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n729), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n801), .A2(new_n756), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n751), .A2(new_n552), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n749), .A2(new_n275), .B1(KEYINPUT46), .B2(new_n971), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n970), .B(new_n972), .C1(G294), .C2(new_n739), .ZN(new_n973));
  AOI22_X1  g0773(.A1(KEYINPUT46), .A2(new_n971), .B1(new_n791), .B2(G303), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n806), .A2(G311), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n280), .B1(new_n733), .B2(G97), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n973), .A2(new_n974), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n967), .B1(new_n969), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT47), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n722), .ZN(new_n980));
  INV_X1    g0780(.A(new_n717), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n723), .B1(new_n208), .B2(new_n413), .C1(new_n981), .C2(new_n239), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n980), .A2(new_n706), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(new_n711), .B2(new_n918), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n958), .A2(new_n985), .ZN(G387));
  NOR2_X1   g0786(.A1(new_n749), .A2(new_n413), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n756), .A2(new_n899), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n740), .A2(new_n324), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n751), .A2(new_n218), .B1(new_n732), .B2(new_n522), .ZN(new_n990));
  NOR4_X1   g0790(.A1(new_n987), .A2(new_n988), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n730), .A2(G150), .ZN(new_n992));
  AOI22_X1  g0792(.A1(G50), .A2(new_n791), .B1(new_n806), .B2(G159), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n991), .A2(new_n280), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n754), .A2(new_n968), .B1(new_n756), .B2(new_n752), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT109), .Z(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n757), .B2(new_n740), .C1(new_n753), .C2(new_n737), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT48), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n254), .B2(new_n751), .C1(new_n749), .C2(new_n801), .ZN(new_n999));
  XNOR2_X1  g0799(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n339), .B1(new_n552), .B2(new_n732), .C1(new_n729), .C2(new_n735), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n994), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n722), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n258), .B1(new_n899), .B2(new_n218), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n662), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1005), .B1(new_n1006), .B2(KEYINPUT108), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(KEYINPUT108), .B2(new_n1006), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n410), .A2(new_n202), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT50), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n717), .B1(new_n1008), .B2(new_n1010), .C1(new_n236), .C2(new_n258), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(G107), .B2(new_n208), .C1(new_n662), .C2(new_n720), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n723), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n650), .A2(new_n652), .A3(new_n711), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1004), .A2(new_n706), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n957), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n952), .A2(new_n700), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(KEYINPUT112), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n947), .B(new_n950), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n701), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n661), .B(KEYINPUT111), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n1017), .B2(KEYINPUT112), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1015), .B1(new_n1016), .B2(new_n952), .C1(new_n1021), .C2(new_n1024), .ZN(G393));
  AOI21_X1  g0825(.A(new_n705), .B1(new_n913), .B2(new_n711), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n749), .A2(new_n552), .B1(new_n254), .B2(new_n756), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(G107), .B2(new_n733), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n739), .A2(G303), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n754), .A2(new_n757), .B1(new_n737), .B2(new_n968), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT52), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n339), .B1(new_n801), .B2(new_n751), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(new_n730), .B2(G322), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1028), .A2(new_n1029), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n280), .B1(new_n732), .B2(new_n582), .C1(new_n400), .C2(new_n751), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n730), .B2(G143), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT113), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n756), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n739), .A2(G50), .B1(new_n1038), .B2(new_n410), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n748), .A2(G77), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1037), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n754), .A2(new_n439), .B1(new_n737), .B2(new_n320), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT51), .Z(new_n1043));
  OAI21_X1  g0843(.A(new_n1034), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n722), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n723), .B1(new_n522), .B2(new_n208), .C1(new_n981), .C2(new_n246), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1026), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n944), .A2(new_n954), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1047), .B1(new_n1048), .B2(new_n1016), .ZN(new_n1049));
  AND2_X1   g0849(.A1(new_n955), .A2(new_n1023), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1048), .A2(new_n1020), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(G390));
  OAI21_X1  g0853(.A(new_n872), .B1(new_n876), .B2(KEYINPUT39), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n709), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n339), .B1(new_n756), .B2(new_n522), .C1(new_n552), .C2(new_n754), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n751), .A2(new_n582), .B1(new_n732), .B2(new_n899), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(new_n748), .B2(G77), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n275), .B2(new_n740), .C1(new_n254), .C2(new_n729), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1056), .B(new_n1059), .C1(G283), .C2(new_n806), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n730), .A2(G125), .B1(G128), .B2(new_n806), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n791), .A2(G132), .B1(new_n733), .B2(G50), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(new_n793), .C2(new_n740), .ZN(new_n1063));
  XOR2_X1   g0863(.A(KEYINPUT54), .B(G143), .Z(new_n1064));
  NAND2_X1  g0864(.A1(new_n1038), .A2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n280), .B(new_n1065), .C1(new_n749), .C2(new_n439), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n965), .A2(G150), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT53), .ZN(new_n1068));
  NOR3_X1   g0868(.A1(new_n1063), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n722), .B1(new_n1060), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n324), .A2(new_n809), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1055), .A2(new_n706), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n781), .A2(new_n605), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n676), .A2(new_n641), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n780), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n868), .B1(new_n1075), .B2(new_n879), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n842), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n776), .A2(new_n783), .A3(new_n879), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n872), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT39), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1079), .B1(new_n842), .B2(new_n1080), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n878), .A2(new_n880), .B1(new_n405), .B2(new_n640), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1077), .B(new_n1078), .C1(new_n1081), .C2(new_n1083), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n1054), .A2(new_n1082), .B1(new_n1076), .B2(new_n842), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n846), .A2(new_n850), .A3(G330), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1084), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1072), .B1(new_n1087), .B2(new_n1016), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n890), .A2(new_n863), .A3(new_n610), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n846), .A2(G330), .A3(new_n783), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n880), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1078), .A2(new_n1091), .A3(new_n780), .A4(new_n1074), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n880), .B1(new_n699), .B2(new_n782), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n1086), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n878), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1089), .B1(new_n1092), .B2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1084), .B(new_n1097), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1092), .A2(new_n1096), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1089), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1022), .B1(new_n1087), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1088), .B1(new_n1098), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(G378));
  NAND2_X1  g0904(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n330), .A2(new_n814), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n358), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n358), .A2(new_n1108), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1107), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1111), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1113), .A2(new_n1109), .A3(new_n1106), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n865), .A2(new_n853), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1115), .B1(new_n865), .B2(new_n853), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n888), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1115), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n846), .A2(new_n850), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n839), .B2(new_n871), .ZN(new_n1121));
  OAI21_X1  g0921(.A(G330), .B1(new_n1121), .B2(KEYINPUT40), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n876), .A2(new_n851), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1119), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n877), .A2(new_n886), .A3(new_n887), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n865), .A2(new_n853), .A3(new_n1115), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1118), .A2(KEYINPUT116), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT116), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1124), .A2(new_n1125), .A3(new_n1129), .A4(new_n1126), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1105), .A2(new_n1128), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT57), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1118), .A2(KEYINPUT118), .A3(new_n1127), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT118), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1124), .A2(new_n1125), .A3(new_n1135), .A4(new_n1126), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1105), .A2(new_n1134), .A3(KEYINPUT57), .A4(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1133), .A2(new_n1023), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT117), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1128), .A2(new_n957), .A3(new_n1130), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n739), .A2(G132), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n748), .A2(G150), .B1(G125), .B2(new_n806), .ZN(new_n1142));
  XOR2_X1   g0942(.A(new_n1142), .B(KEYINPUT115), .Z(new_n1143));
  AOI211_X1 g0943(.A(new_n1141), .B(new_n1143), .C1(new_n965), .C2(new_n1064), .ZN(new_n1144));
  INV_X1    g0944(.A(G128), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1144), .B1(new_n1145), .B2(new_n754), .C1(new_n793), .C2(new_n756), .ZN(new_n1146));
  OR2_X1    g0946(.A1(new_n1146), .A2(KEYINPUT59), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n733), .A2(G159), .ZN(new_n1148));
  AOI21_X1  g0948(.A(G41), .B1(new_n730), .B2(G124), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1147), .A2(new_n253), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1146), .A2(KEYINPUT59), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT58), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n751), .A2(new_n218), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n730), .A2(G283), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n739), .A2(G97), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n412), .A2(new_n1038), .B1(new_n733), .B2(G58), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1154), .A2(new_n959), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1153), .B(new_n1157), .C1(G107), .C2(new_n791), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n806), .A2(G116), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1158), .A2(new_n335), .A3(new_n339), .A4(new_n1159), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n1150), .A2(new_n1151), .B1(new_n1152), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(G50), .B1(new_n279), .B2(new_n335), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(new_n1160), .B2(new_n1152), .ZN(new_n1163));
  XOR2_X1   g0963(.A(new_n1163), .B(KEYINPUT114), .Z(new_n1164));
  OAI21_X1  g0964(.A(new_n722), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n705), .B1(new_n1115), .B2(new_n709), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n809), .A2(new_n202), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1139), .B1(new_n1140), .B2(new_n1168), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n1140), .A2(new_n1139), .A3(new_n1168), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1138), .B1(new_n1169), .B2(new_n1170), .ZN(G375));
  NAND3_X1  g0971(.A1(new_n1092), .A2(new_n1096), .A3(new_n1089), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n1101), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n931), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT119), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n880), .A2(new_n708), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n809), .A2(new_n899), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n749), .A2(new_n202), .B1(new_n793), .B2(new_n754), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(G132), .B2(new_n806), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n739), .A2(new_n1064), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n280), .B1(new_n732), .B2(new_n216), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT122), .Z(new_n1183));
  OAI22_X1  g0983(.A1(new_n729), .A2(new_n1145), .B1(new_n439), .B2(new_n751), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(G150), .B2(new_n1038), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1180), .A2(new_n1181), .A3(new_n1183), .A4(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n987), .B1(G283), .B2(new_n791), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT121), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n963), .B(new_n1188), .C1(G107), .C2(new_n1038), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n339), .B1(new_n729), .B2(new_n752), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(G294), .B2(new_n806), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1189), .B(new_n1191), .C1(new_n552), .C2(new_n740), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n751), .A2(new_n522), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1186), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n705), .B(new_n1178), .C1(new_n722), .C2(new_n1194), .ZN(new_n1195));
  XOR2_X1   g0995(.A(new_n957), .B(KEYINPUT120), .Z(new_n1196));
  AOI21_X1  g0996(.A(new_n1195), .B1(new_n1099), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1175), .A2(new_n1197), .ZN(G381));
  NOR2_X1   g0998(.A1(G375), .A2(G378), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(G381), .A2(G384), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n958), .A2(new_n1052), .A3(new_n985), .ZN(new_n1201));
  NOR3_X1   g1001(.A1(new_n1201), .A2(G396), .A3(G393), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1199), .A2(new_n1200), .A3(new_n1202), .ZN(G407));
  NAND2_X1  g1003(.A1(new_n1199), .A2(new_n639), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(G407), .A2(G213), .A3(new_n1204), .ZN(G409));
  INV_X1    g1005(.A(KEYINPUT60), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1022), .B1(new_n1172), .B2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n1173), .B2(new_n1206), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n1197), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1209), .A2(new_n788), .A3(new_n811), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1208), .A2(G384), .A3(new_n1197), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n639), .A2(G213), .A3(G2897), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1212), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1138), .B(G378), .C1(new_n1169), .C2(new_n1170), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1105), .A2(new_n1128), .A3(new_n931), .A4(new_n1130), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1134), .A2(new_n1136), .A3(new_n1196), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1217), .A2(new_n1168), .A3(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(KEYINPUT123), .B1(new_n1219), .B2(new_n1103), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1219), .A2(KEYINPUT123), .A3(new_n1103), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1216), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n639), .A2(G213), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1215), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(KEYINPUT127), .B1(new_n1225), .B2(KEYINPUT61), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT127), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT61), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1219), .A2(KEYINPUT123), .A3(new_n1103), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1229), .A2(new_n1220), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1230), .A2(new_n1216), .B1(G213), .B2(new_n639), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1227), .B(new_n1228), .C1(new_n1231), .C2(new_n1215), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1223), .A2(new_n1233), .A3(new_n1224), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(KEYINPUT62), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT62), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1231), .A2(new_n1236), .A3(new_n1233), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1226), .A2(new_n1232), .A3(new_n1235), .A4(new_n1237), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(G393), .B(G396), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1201), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1052), .B1(new_n958), .B2(new_n985), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1239), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(G387), .A2(G390), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(G393), .B(new_n774), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1243), .A2(new_n1244), .A3(new_n1201), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1242), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1238), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT126), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n1246), .B2(new_n1228), .ZN(new_n1250));
  AOI211_X1 g1050(.A(KEYINPUT126), .B(KEYINPUT61), .C1(new_n1242), .C2(new_n1245), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT63), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1234), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT124), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1252), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT125), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1231), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(KEYINPUT125), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1215), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1258), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1231), .A2(KEYINPUT63), .A3(new_n1233), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1234), .A2(KEYINPUT124), .A3(new_n1253), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1256), .A2(new_n1262), .A3(new_n1263), .A4(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1248), .A2(new_n1265), .ZN(G405));
  XNOR2_X1  g1066(.A(G375), .B(new_n1103), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1233), .ZN(new_n1268));
  OR2_X1    g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(new_n1271), .B(new_n1246), .ZN(G402));
endmodule


