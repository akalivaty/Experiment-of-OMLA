//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n820, new_n821,
    new_n822, new_n823, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  AND2_X1   g004(.A1(new_n205), .A2(G8gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(G8gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT85), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT14), .B(G29gat), .ZN(new_n211));
  INV_X1    g010(.A(G36gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G29gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G43gat), .B(G50gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT15), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n210), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n217), .A2(KEYINPUT15), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n220), .A2(KEYINPUT85), .A3(new_n213), .A4(new_n215), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n217), .A2(KEYINPUT15), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT86), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n222), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  AOI22_X1  g023(.A1(KEYINPUT86), .A2(new_n218), .B1(new_n213), .B2(new_n215), .ZN(new_n225));
  AOI22_X1  g024(.A1(new_n219), .A2(new_n221), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n209), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G229gat), .A2(G233gat), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n226), .A2(KEYINPUT17), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n208), .B1(new_n226), .B2(KEYINPUT17), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n228), .B(new_n229), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT18), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n208), .A2(new_n226), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n228), .A2(new_n235), .A3(KEYINPUT87), .ZN(new_n236));
  XOR2_X1   g035(.A(new_n229), .B(KEYINPUT13), .Z(new_n237));
  OR3_X1    g036(.A1(new_n208), .A2(new_n226), .A3(KEYINPUT87), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n232), .A2(new_n233), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n234), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G113gat), .B(G141gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT84), .B(G197gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g043(.A(KEYINPUT11), .B(G169gat), .Z(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(KEYINPUT12), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n241), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n234), .A2(new_n240), .A3(new_n239), .A4(new_n247), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AND2_X1   g050(.A1(G71gat), .A2(G78gat), .ZN(new_n252));
  NOR2_X1   g051(.A1(G71gat), .A2(G78gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G57gat), .B(G64gat), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G57gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(G64gat), .ZN(new_n259));
  INV_X1    g058(.A(G64gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G57gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G71gat), .B(G78gat), .ZN(new_n263));
  INV_X1    g062(.A(new_n256), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n257), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT21), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G231gat), .A2(G233gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(G127gat), .B(G155gat), .Z(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT20), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n270), .B(new_n272), .Z(new_n273));
  XNOR2_X1  g072(.A(G183gat), .B(G211gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT89), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n266), .B(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n208), .B1(new_n278), .B2(new_n267), .ZN(new_n279));
  XOR2_X1   g078(.A(new_n279), .B(KEYINPUT90), .Z(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n280), .B(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n276), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n280), .B(new_n281), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(new_n275), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G99gat), .A2(G106gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT8), .ZN(new_n290));
  NAND2_X1  g089(.A1(G85gat), .A2(G92gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT7), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G85gat), .ZN(new_n294));
  INV_X1    g093(.A(G92gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n290), .A2(new_n293), .A3(new_n296), .A4(new_n297), .ZN(new_n298));
  OR2_X1    g097(.A1(G99gat), .A2(G106gat), .ZN(new_n299));
  AND2_X1   g098(.A1(new_n299), .A2(new_n289), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n289), .ZN(new_n302));
  AND3_X1   g101(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI22_X1  g104(.A1(KEYINPUT8), .A2(new_n289), .B1(new_n294), .B2(new_n295), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n302), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  AND2_X1   g107(.A1(G232gat), .A2(G233gat), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n227), .A2(new_n308), .B1(KEYINPUT41), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n298), .A2(new_n300), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n305), .A2(new_n302), .A3(new_n306), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n313), .B1(new_n226), .B2(KEYINPUT17), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n310), .B1(new_n314), .B2(new_n230), .ZN(new_n315));
  XNOR2_X1  g114(.A(G190gat), .B(G218gat), .ZN(new_n316));
  XOR2_X1   g115(.A(new_n316), .B(KEYINPUT91), .Z(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n309), .A2(KEYINPUT41), .ZN(new_n319));
  XNOR2_X1  g118(.A(G134gat), .B(G162gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n319), .B(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n317), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n310), .B(new_n322), .C1(new_n314), .C2(new_n230), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n318), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n321), .B1(new_n318), .B2(new_n323), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n288), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT92), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n299), .A2(new_n329), .A3(new_n289), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n257), .A2(new_n265), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n308), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT10), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n257), .A2(new_n265), .A3(new_n330), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n313), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n332), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT93), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT93), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n332), .A2(new_n338), .A3(new_n333), .A4(new_n335), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n308), .A2(KEYINPUT10), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n278), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT94), .ZN(new_n345));
  NAND2_X1  g144(.A1(G230gat), .A2(G233gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n342), .B1(new_n337), .B2(new_n339), .ZN(new_n348));
  INV_X1    g147(.A(new_n346), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT94), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G120gat), .B(G148gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n351), .B(KEYINPUT96), .ZN(new_n352));
  XOR2_X1   g151(.A(G176gat), .B(G204gat), .Z(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n332), .A2(new_n335), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(new_n349), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n354), .B1(new_n356), .B2(KEYINPUT95), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n357), .B1(KEYINPUT95), .B2(new_n356), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n347), .A2(new_n350), .A3(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n354), .B(KEYINPUT97), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n348), .A2(new_n349), .ZN(new_n361));
  INV_X1    g160(.A(new_n356), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n328), .A2(new_n364), .ZN(new_n365));
  XOR2_X1   g164(.A(G197gat), .B(G204gat), .Z(new_n366));
  AOI21_X1  g165(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G211gat), .B(G218gat), .ZN(new_n369));
  OR2_X1    g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n369), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G169gat), .A2(G176gat), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT65), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G169gat), .ZN(new_n377));
  INV_X1    g176(.A(G176gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OR2_X1    g178(.A1(new_n379), .A2(KEYINPUT26), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(KEYINPUT26), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n376), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(G183gat), .A2(G190gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT66), .ZN(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT27), .B(G183gat), .ZN(new_n386));
  INV_X1    g185(.A(G190gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n388), .B(KEYINPUT28), .Z(new_n389));
  INV_X1    g188(.A(KEYINPUT66), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n382), .A2(new_n390), .A3(new_n383), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n385), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT23), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n379), .A2(new_n393), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n376), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n387), .A2(G183gat), .ZN(new_n396));
  INV_X1    g195(.A(G183gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n397), .A2(G190gat), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT24), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  OR2_X1    g198(.A1(new_n383), .A2(KEYINPUT24), .ZN(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT64), .B(G176gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n377), .A2(KEYINPUT23), .ZN(new_n402));
  OR2_X1    g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n395), .A2(new_n399), .A3(new_n400), .A4(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT25), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n377), .A2(new_n378), .A3(KEYINPUT23), .ZN(new_n406));
  AND4_X1   g205(.A1(KEYINPUT25), .A2(new_n399), .A3(new_n400), .A4(new_n406), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n404), .A2(new_n405), .B1(new_n395), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(KEYINPUT70), .B1(new_n392), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n404), .A2(new_n405), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n407), .A2(new_n395), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT70), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n385), .A2(new_n389), .A3(new_n391), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT29), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n409), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(G226gat), .A2(G233gat), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n417), .A2(KEYINPUT71), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n412), .A2(new_n414), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n420), .A2(G226gat), .A3(G233gat), .ZN(new_n421));
  AOI22_X1  g220(.A1(new_n417), .A2(new_n418), .B1(KEYINPUT71), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n373), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n420), .A2(new_n416), .A3(new_n418), .ZN(new_n424));
  AND2_X1   g223(.A1(new_n409), .A2(new_n415), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n424), .B1(new_n425), .B2(new_n418), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n372), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n423), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G8gat), .B(G36gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(G64gat), .B(G92gat), .ZN(new_n430));
  XOR2_X1   g229(.A(new_n429), .B(new_n430), .Z(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n423), .A2(new_n431), .A3(new_n427), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(KEYINPUT30), .A3(new_n434), .ZN(new_n435));
  OR3_X1    g234(.A1(new_n428), .A2(KEYINPUT30), .A3(new_n432), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  XOR2_X1   g236(.A(G141gat), .B(G148gat), .Z(new_n438));
  INV_X1    g237(.A(G155gat), .ZN(new_n439));
  INV_X1    g238(.A(G162gat), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT2), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(G155gat), .B(G162gat), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n438), .A2(new_n443), .A3(new_n441), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(G113gat), .ZN(new_n448));
  INV_X1    g247(.A(G120gat), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT1), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(G127gat), .B(G134gat), .ZN(new_n451));
  XOR2_X1   g250(.A(KEYINPUT67), .B(G120gat), .Z(new_n452));
  OAI211_X1 g251(.A(new_n450), .B(new_n451), .C1(new_n452), .C2(new_n448), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n450), .B1(new_n448), .B2(new_n449), .ZN(new_n454));
  INV_X1    g253(.A(new_n451), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n447), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n445), .A2(new_n446), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n453), .A2(new_n456), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(G225gat), .A2(G233gat), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(KEYINPUT74), .B(KEYINPUT5), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(KEYINPUT72), .B1(new_n459), .B2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n459), .A2(KEYINPUT72), .A3(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n460), .B1(new_n459), .B2(KEYINPUT3), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n464), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n459), .A2(new_n460), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT4), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT73), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n476), .A2(KEYINPUT73), .A3(new_n477), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n458), .A2(KEYINPUT4), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n468), .B1(new_n475), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G1gat), .B(G29gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(KEYINPUT0), .ZN(new_n487));
  XNOR2_X1  g286(.A(G57gat), .B(G85gat), .ZN(new_n488));
  XOR2_X1   g287(.A(new_n487), .B(new_n488), .Z(new_n489));
  AOI21_X1  g288(.A(new_n467), .B1(new_n482), .B2(new_n478), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n485), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT6), .ZN(new_n493));
  INV_X1    g292(.A(new_n489), .ZN(new_n494));
  INV_X1    g293(.A(new_n491), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n494), .B1(new_n495), .B2(new_n484), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n492), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  OAI211_X1 g296(.A(KEYINPUT6), .B(new_n494), .C1(new_n495), .C2(new_n484), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n437), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT75), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT3), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n373), .A2(KEYINPUT29), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n503), .B1(new_n504), .B2(KEYINPUT77), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n372), .A2(KEYINPUT77), .A3(new_n416), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n459), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n416), .B1(new_n459), .B2(KEYINPUT3), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n373), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n507), .A2(G228gat), .A3(G233gat), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(G228gat), .A2(G233gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT76), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n373), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n513), .B(new_n416), .C1(new_n512), .C2(new_n370), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n447), .B1(new_n514), .B2(new_n503), .ZN(new_n515));
  INV_X1    g314(.A(new_n509), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n511), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n510), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(G22gat), .ZN(new_n519));
  INV_X1    g318(.A(G22gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n510), .A2(new_n517), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n521), .A2(KEYINPUT78), .ZN(new_n523));
  XNOR2_X1  g322(.A(G78gat), .B(G106gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(KEYINPUT31), .B(G50gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n522), .B1(new_n523), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT78), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n519), .A2(new_n529), .A3(new_n521), .A4(new_n526), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n437), .A2(KEYINPUT75), .A3(new_n499), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n502), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n471), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n474), .B1(new_n534), .B2(new_n469), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n482), .A2(new_n478), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT79), .B1(new_n537), .B2(new_n464), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT79), .ZN(new_n539));
  AOI211_X1 g338(.A(new_n539), .B(new_n463), .C1(new_n535), .C2(new_n536), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n458), .A2(new_n463), .A3(new_n461), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT81), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n542), .A2(new_n543), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n541), .A2(KEYINPUT39), .A3(new_n544), .A4(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT39), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(new_n538), .B2(new_n540), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT80), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n548), .A2(new_n549), .A3(new_n489), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n549), .B1(new_n548), .B2(new_n489), .ZN(new_n551));
  OAI211_X1 g350(.A(KEYINPUT40), .B(new_n546), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n496), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n548), .A2(new_n489), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT80), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n548), .A2(new_n549), .A3(new_n489), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT40), .B1(new_n557), .B2(new_n546), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  AND2_X1   g358(.A1(new_n435), .A2(new_n436), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n531), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT83), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n372), .B1(new_n419), .B2(new_n422), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT37), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n564), .B1(new_n426), .B2(new_n373), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT82), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n563), .A2(new_n565), .A3(KEYINPUT82), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT38), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n431), .B1(new_n423), .B2(new_n427), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n431), .A2(new_n564), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n562), .B1(new_n570), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n574), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n568), .A2(new_n569), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n576), .A2(KEYINPUT83), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n434), .A2(new_n498), .A3(new_n497), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n428), .A2(KEYINPUT37), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n580), .B1(new_n572), .B2(new_n573), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n579), .B1(new_n581), .B2(KEYINPUT38), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n575), .A2(new_n578), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n561), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G15gat), .B(G43gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(G71gat), .B(G99gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n457), .B1(new_n392), .B2(new_n408), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n412), .A2(new_n460), .A3(new_n414), .ZN(new_n589));
  INV_X1    g388(.A(G227gat), .ZN(new_n590));
  INV_X1    g389(.A(G233gat), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n588), .A2(new_n589), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n587), .B1(new_n593), .B2(KEYINPUT32), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT33), .ZN(new_n595));
  AND3_X1   g394(.A1(new_n593), .A2(KEYINPUT68), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT68), .B1(new_n593), .B2(new_n595), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n594), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n592), .B1(new_n588), .B2(new_n589), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT34), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n593), .B(KEYINPUT32), .C1(new_n595), .C2(new_n587), .ZN(new_n601));
  AND3_X1   g400(.A1(new_n598), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n600), .B1(new_n598), .B2(new_n601), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT36), .ZN(new_n604));
  NOR3_X1   g403(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT69), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n606), .B1(new_n602), .B2(new_n603), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n598), .A2(new_n600), .A3(new_n601), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT69), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n605), .B1(new_n610), .B2(new_n604), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  AND3_X1   g411(.A1(new_n533), .A2(new_n584), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n528), .A2(new_n530), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT35), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n500), .A2(new_n616), .A3(new_n610), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n602), .A2(new_n603), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(KEYINPUT75), .B1(new_n437), .B2(new_n499), .ZN(new_n621));
  INV_X1    g420(.A(new_n499), .ZN(new_n622));
  AOI211_X1 g421(.A(new_n501), .B(new_n622), .C1(new_n435), .C2(new_n436), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n620), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n617), .B1(new_n624), .B2(KEYINPUT35), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n251), .B(new_n365), .C1(new_n613), .C2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT98), .ZN(new_n627));
  INV_X1    g426(.A(new_n251), .ZN(new_n628));
  INV_X1    g427(.A(new_n617), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n619), .B1(new_n502), .B2(new_n532), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n629), .B1(new_n630), .B2(new_n615), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n611), .B1(new_n561), .B2(new_n583), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n533), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n628), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT98), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n634), .A2(new_n635), .A3(new_n365), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n627), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n622), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g438(.A(KEYINPUT16), .B(G8gat), .Z(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  AOI211_X1 g440(.A(new_n437), .B(new_n641), .C1(new_n627), .C2(new_n636), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n637), .A2(new_n560), .ZN(new_n643));
  AOI22_X1  g442(.A1(new_n642), .A2(KEYINPUT42), .B1(new_n643), .B2(G8gat), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n626), .A2(KEYINPUT98), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n635), .B1(new_n634), .B2(new_n365), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n560), .B(new_n640), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT99), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT42), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n648), .B1(new_n647), .B2(new_n649), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n644), .B1(new_n650), .B2(new_n651), .ZN(G1325gat));
  INV_X1    g451(.A(new_n637), .ZN(new_n653));
  OAI21_X1  g452(.A(G15gat), .B1(new_n653), .B2(new_n612), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n610), .A2(G15gat), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n654), .B1(new_n653), .B2(new_n655), .ZN(G1326gat));
  NAND2_X1  g455(.A1(new_n637), .A2(new_n531), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT43), .B(G22gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(G1327gat));
  NAND2_X1  g458(.A1(new_n624), .A2(KEYINPUT35), .ZN(new_n660));
  AOI22_X1  g459(.A1(new_n660), .A2(new_n629), .B1(new_n632), .B2(new_n533), .ZN(new_n661));
  INV_X1    g460(.A(new_n364), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n287), .A2(new_n662), .ZN(new_n663));
  NOR4_X1   g462(.A1(new_n661), .A2(new_n628), .A3(new_n327), .A4(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT100), .B(KEYINPUT45), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n622), .A2(new_n214), .ZN(new_n667));
  OR3_X1    g466(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n666), .B1(new_n665), .B2(new_n667), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n670), .B1(new_n661), .B2(new_n327), .ZN(new_n671));
  OAI211_X1 g470(.A(KEYINPUT44), .B(new_n326), .C1(new_n613), .C2(new_n625), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n663), .A2(new_n628), .ZN(new_n674));
  AND3_X1   g473(.A1(new_n673), .A2(new_n622), .A3(new_n674), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n668), .B(new_n669), .C1(new_n675), .C2(new_n214), .ZN(G1328gat));
  NAND2_X1  g475(.A1(new_n560), .A2(new_n212), .ZN(new_n677));
  OR3_X1    g476(.A1(new_n665), .A2(KEYINPUT46), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(KEYINPUT46), .B1(new_n665), .B2(new_n677), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n673), .A2(new_n560), .A3(new_n674), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n678), .B(new_n679), .C1(new_n680), .C2(new_n212), .ZN(G1329gat));
  NOR2_X1   g480(.A1(new_n610), .A2(G43gat), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n664), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT47), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n671), .A2(new_n611), .A3(new_n672), .A4(new_n674), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(KEYINPUT102), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(G43gat), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n686), .A2(KEYINPUT102), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n685), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT101), .B(KEYINPUT47), .Z(new_n691));
  AND2_X1   g490(.A1(new_n686), .A2(G43gat), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n691), .B1(new_n692), .B2(new_n683), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n690), .A2(new_n693), .ZN(G1330gat));
  NAND4_X1  g493(.A1(new_n673), .A2(G50gat), .A3(new_n531), .A4(new_n674), .ZN(new_n695));
  INV_X1    g494(.A(G50gat), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n696), .B1(new_n665), .B2(new_n614), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(KEYINPUT48), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT48), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n695), .A2(new_n697), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(new_n701), .ZN(G1331gat));
  INV_X1    g501(.A(KEYINPUT103), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n328), .A2(new_n251), .A3(new_n662), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n703), .B1(new_n661), .B2(new_n705), .ZN(new_n706));
  OAI211_X1 g505(.A(KEYINPUT103), .B(new_n704), .C1(new_n613), .C2(new_n625), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n708), .A2(new_n499), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(new_n258), .ZN(G1332gat));
  AOI21_X1  g509(.A(new_n437), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT104), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(G1333gat));
  NAND3_X1  g514(.A1(new_n706), .A2(new_n707), .A3(new_n611), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G71gat), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n610), .A2(G71gat), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n706), .A2(new_n707), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT50), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1334gat));
  NOR2_X1   g521(.A1(new_n708), .A2(new_n614), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n723), .B(G78gat), .Z(G1335gat));
  NOR3_X1   g523(.A1(new_n288), .A2(new_n251), .A3(new_n662), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n671), .A2(new_n622), .A3(new_n672), .A4(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(G85gat), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n622), .A2(new_n294), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n288), .A2(new_n251), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n326), .B(new_n730), .C1(new_n613), .C2(new_n625), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT51), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n327), .B1(new_n631), .B2(new_n633), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n734), .A2(KEYINPUT51), .A3(new_n730), .ZN(new_n735));
  AOI211_X1 g534(.A(new_n662), .B(new_n729), .C1(new_n733), .C2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(KEYINPUT105), .B1(new_n728), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT105), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n733), .A2(new_n735), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n364), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n738), .B(new_n727), .C1(new_n740), .C2(new_n729), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n737), .A2(new_n741), .ZN(G1336gat));
  INV_X1    g541(.A(KEYINPUT52), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(KEYINPUT106), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n671), .A2(new_n560), .A3(new_n672), .A4(new_n725), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G92gat), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n560), .A2(new_n364), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n747), .A2(G92gat), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n731), .A2(new_n732), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT51), .B1(new_n734), .B2(new_n730), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n743), .A2(KEYINPUT106), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  AND4_X1   g552(.A1(new_n744), .A2(new_n746), .A3(new_n751), .A4(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n752), .B1(new_n739), .B2(new_n748), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n744), .B1(new_n755), .B2(new_n746), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n754), .A2(new_n756), .ZN(G1337gat));
  AND3_X1   g556(.A1(new_n673), .A2(new_n611), .A3(new_n725), .ZN(new_n758));
  INV_X1    g557(.A(G99gat), .ZN(new_n759));
  INV_X1    g558(.A(new_n610), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n759), .ZN(new_n761));
  OAI22_X1  g560(.A1(new_n758), .A2(new_n759), .B1(new_n740), .B2(new_n761), .ZN(G1338gat));
  NOR3_X1   g561(.A1(new_n614), .A2(G106gat), .A3(new_n662), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n739), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n671), .A2(new_n531), .A3(new_n672), .A4(new_n725), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G106gat), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n764), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n763), .B(KEYINPUT107), .ZN(new_n769));
  AOI22_X1  g568(.A1(new_n739), .A2(new_n769), .B1(new_n765), .B2(G106gat), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n768), .B1(new_n770), .B2(new_n767), .ZN(G1339gat));
  INV_X1    g570(.A(KEYINPUT54), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n772), .B1(new_n348), .B2(new_n349), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n347), .A2(new_n350), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n354), .B1(new_n361), .B2(new_n772), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n774), .A2(KEYINPUT55), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT108), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT108), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n774), .A2(new_n778), .A3(new_n775), .A4(KEYINPUT55), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n774), .A2(new_n775), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n780), .A2(new_n251), .A3(new_n359), .A4(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n228), .B1(new_n230), .B2(new_n231), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n785), .A2(G229gat), .A3(G233gat), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n237), .B1(new_n236), .B2(new_n238), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT109), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AOI211_X1 g588(.A(KEYINPUT109), .B(new_n237), .C1(new_n236), .C2(new_n238), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n246), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n791), .A2(new_n250), .A3(new_n364), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n326), .B1(new_n784), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n780), .A2(new_n359), .A3(new_n783), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n791), .A2(new_n326), .A3(new_n250), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n287), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n365), .A2(new_n628), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n499), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n620), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n800), .A2(KEYINPUT111), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n560), .B1(new_n800), .B2(KEYINPUT111), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(G113gat), .B1(new_n804), .B2(new_n251), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT110), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n797), .A2(new_n798), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n806), .B1(new_n807), .B2(new_n614), .ZN(new_n808));
  AOI211_X1 g607(.A(KEYINPUT110), .B(new_n531), .C1(new_n797), .C2(new_n798), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n560), .A2(new_n499), .A3(new_n610), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n628), .A2(new_n448), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n805), .B1(new_n813), .B2(new_n814), .ZN(G1340gat));
  OAI21_X1  g614(.A(G120gat), .B1(new_n812), .B2(new_n662), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n364), .A2(new_n452), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n816), .B1(new_n803), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(KEYINPUT112), .ZN(G1341gat));
  INV_X1    g618(.A(G127gat), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n804), .A2(new_n820), .A3(new_n288), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n813), .A2(new_n288), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n821), .B1(new_n823), .B2(new_n820), .ZN(G1342gat));
  OAI21_X1  g623(.A(G134gat), .B1(new_n812), .B2(new_n327), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n327), .A2(G134gat), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n804), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT113), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n828), .B1(new_n827), .B2(KEYINPUT56), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT56), .ZN(new_n830));
  AOI211_X1 g629(.A(KEYINPUT113), .B(new_n830), .C1(new_n804), .C2(new_n826), .ZN(new_n831));
  OAI221_X1 g630(.A(new_n825), .B1(KEYINPUT56), .B2(new_n827), .C1(new_n829), .C2(new_n831), .ZN(G1343gat));
  NOR3_X1   g631(.A1(new_n611), .A2(new_n499), .A3(new_n560), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT57), .B1(new_n807), .B2(new_n531), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n531), .A2(KEYINPUT57), .ZN(new_n835));
  XNOR2_X1  g634(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n781), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n780), .A2(new_n251), .A3(new_n359), .A4(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n326), .B1(new_n838), .B2(new_n792), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n287), .B1(new_n839), .B2(new_n796), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n835), .B1(new_n840), .B2(new_n798), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n251), .B(new_n833), .C1(new_n834), .C2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(G141gat), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n611), .A2(new_n614), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n799), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n628), .A2(G141gat), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n437), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n843), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT58), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT116), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT58), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT115), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n845), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n799), .A2(KEYINPUT115), .A3(new_n844), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n853), .A2(new_n437), .A3(new_n846), .A4(new_n854), .ZN(new_n855));
  AND4_X1   g654(.A1(new_n850), .A2(new_n843), .A3(new_n851), .A4(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT58), .B1(new_n842), .B2(G141gat), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n850), .B1(new_n857), .B2(new_n855), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n849), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n849), .B(KEYINPUT117), .C1(new_n856), .C2(new_n858), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(G1344gat));
  NAND3_X1  g662(.A1(new_n807), .A2(KEYINPUT57), .A3(new_n531), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n614), .B1(new_n840), .B2(new_n798), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n864), .B1(KEYINPUT57), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n364), .A3(new_n833), .ZN(new_n867));
  AND2_X1   g666(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n834), .A2(new_n841), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870));
  AND3_X1   g669(.A1(new_n833), .A2(new_n870), .A3(new_n364), .ZN(new_n871));
  AOI22_X1  g670(.A1(new_n867), .A2(new_n868), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n853), .A2(new_n437), .A3(new_n854), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n870), .B1(new_n874), .B2(new_n364), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n872), .B1(new_n875), .B2(G148gat), .ZN(G1345gat));
  NAND3_X1  g675(.A1(new_n874), .A2(new_n439), .A3(new_n288), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n869), .A2(new_n288), .A3(new_n833), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(G155gat), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(new_n879), .ZN(G1346gat));
  OAI21_X1  g679(.A(new_n440), .B1(new_n873), .B2(new_n327), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n869), .A2(G162gat), .A3(new_n326), .A4(new_n833), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT118), .ZN(G1347gat));
  NAND2_X1  g683(.A1(new_n807), .A2(new_n499), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT119), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n886), .A2(new_n620), .A3(new_n560), .ZN(new_n887));
  AOI21_X1  g686(.A(G169gat), .B1(new_n887), .B2(new_n251), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n760), .A2(new_n560), .A3(new_n499), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT120), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n890), .B1(new_n808), .B2(new_n809), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT121), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g692(.A(KEYINPUT121), .B(new_n890), .C1(new_n808), .C2(new_n809), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n628), .A2(new_n377), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n888), .B1(new_n895), .B2(new_n896), .ZN(G1348gat));
  AOI21_X1  g696(.A(G176gat), .B1(new_n887), .B2(new_n364), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n364), .A2(new_n401), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n895), .B2(new_n899), .ZN(G1349gat));
  INV_X1    g699(.A(KEYINPUT122), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n288), .A2(new_n386), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n901), .B1(new_n887), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n893), .A2(new_n288), .A3(new_n894), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(G183gat), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(KEYINPUT60), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT60), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n903), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(G1350gat));
  NAND3_X1  g709(.A1(new_n893), .A2(new_n326), .A3(new_n894), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(G190gat), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT61), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n911), .A2(KEYINPUT61), .A3(G190gat), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT123), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n327), .A2(G190gat), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n887), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n916), .B1(new_n887), .B2(new_n917), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n914), .B(new_n915), .C1(new_n918), .C2(new_n919), .ZN(G1351gat));
  NOR3_X1   g719(.A1(new_n611), .A2(new_n622), .A3(new_n437), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n866), .A2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(G197gat), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n922), .A2(new_n923), .A3(new_n628), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n886), .A2(new_n560), .A3(new_n844), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n251), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n924), .B1(new_n927), .B2(new_n923), .ZN(G1352gat));
  XOR2_X1   g727(.A(KEYINPUT124), .B(G204gat), .Z(new_n929));
  NOR2_X1   g728(.A1(new_n747), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n886), .A2(new_n844), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT62), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n929), .B1(new_n922), .B2(new_n662), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT62), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n886), .A2(new_n934), .A3(new_n844), .A4(new_n930), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n932), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n936), .B(new_n937), .ZN(G1353gat));
  NOR2_X1   g737(.A1(new_n287), .A2(G211gat), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n926), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n866), .A2(new_n288), .A3(new_n921), .ZN(new_n941));
  AND3_X1   g740(.A1(new_n941), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n942));
  AOI21_X1  g741(.A(KEYINPUT63), .B1(new_n941), .B2(G211gat), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(KEYINPUT126), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT126), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n940), .B(new_n946), .C1(new_n943), .C2(new_n942), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n947), .ZN(G1354gat));
  INV_X1    g747(.A(G218gat), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n922), .A2(new_n949), .A3(new_n327), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n949), .B1(new_n925), .B2(new_n327), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n952), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n950), .B1(new_n953), .B2(new_n954), .ZN(G1355gat));
endmodule


