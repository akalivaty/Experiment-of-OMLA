//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 1 0 1 0 0 1 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 0 1 0 0 0 0 0 0 1 1 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1006, new_n1007, new_n1008, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT88), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT67), .A2(G953), .ZN(new_n193));
  AND2_X1   g007(.A1(KEYINPUT66), .A2(G237), .ZN(new_n194));
  NOR2_X1   g008(.A1(KEYINPUT66), .A2(G237), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n192), .B(new_n193), .C1(new_n194), .C2(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(G214), .B1(KEYINPUT88), .B2(G143), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n189), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  XOR2_X1   g012(.A(KEYINPUT67), .B(G953), .Z(new_n199));
  XNOR2_X1  g013(.A(KEYINPUT66), .B(G237), .ZN(new_n200));
  INV_X1    g014(.A(new_n197), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n199), .A2(new_n200), .A3(new_n188), .A4(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G131), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT17), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n198), .A2(G131), .A3(new_n202), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G140), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G125), .ZN(new_n210));
  INV_X1    g024(.A(G125), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G140), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n210), .A2(new_n212), .A3(KEYINPUT16), .ZN(new_n213));
  OR3_X1    g027(.A1(new_n211), .A2(KEYINPUT16), .A3(G140), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(G146), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT74), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT74), .A4(G146), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n213), .A2(new_n214), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n217), .B(new_n218), .C1(G146), .C2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n198), .A2(new_n202), .A3(KEYINPUT17), .A4(G131), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n208), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(G113), .B(G122), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT91), .B(G104), .ZN(new_n225));
  XOR2_X1   g039(.A(new_n224), .B(new_n225), .Z(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT18), .A2(G131), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n198), .A2(new_n229), .A3(new_n202), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT89), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT89), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n198), .A2(new_n202), .A3(new_n232), .A4(new_n229), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(G125), .B(G140), .ZN(new_n235));
  INV_X1    g049(.A(G146), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n210), .A2(new_n212), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G146), .ZN(new_n239));
  AOI22_X1  g053(.A1(new_n203), .A2(new_n228), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n234), .A2(new_n240), .ZN(new_n241));
  AND3_X1   g055(.A1(new_n223), .A2(new_n227), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n227), .B1(new_n223), .B2(new_n241), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n187), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT92), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OAI211_X1 g060(.A(KEYINPUT92), .B(new_n187), .C1(new_n242), .C2(new_n243), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(G475), .A3(new_n247), .ZN(new_n248));
  XOR2_X1   g062(.A(G116), .B(G122), .Z(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G107), .ZN(new_n250));
  XNOR2_X1  g064(.A(G116), .B(G122), .ZN(new_n251));
  INV_X1    g065(.A(G107), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G128), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G143), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n255), .A2(G143), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n256), .B1(new_n257), .B2(KEYINPUT13), .ZN(new_n258));
  INV_X1    g072(.A(G143), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G128), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT13), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(G134), .B1(new_n258), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G134), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n260), .A2(new_n256), .A3(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n254), .A2(new_n263), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G116), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(KEYINPUT14), .A3(G122), .ZN(new_n268));
  OAI211_X1 g082(.A(G107), .B(new_n268), .C1(new_n249), .C2(KEYINPUT14), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT93), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n253), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n259), .A2(G128), .ZN(new_n272));
  OAI21_X1  g086(.A(G134), .B1(new_n257), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n265), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n251), .A2(KEYINPUT93), .A3(new_n252), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n269), .A2(new_n271), .A3(new_n274), .A4(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n266), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT94), .ZN(new_n278));
  XOR2_X1   g092(.A(KEYINPUT9), .B(G234), .Z(new_n279));
  NAND3_X1  g093(.A1(new_n279), .A2(G217), .A3(new_n191), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT94), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n266), .A2(new_n276), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n278), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n280), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n277), .A2(KEYINPUT94), .A3(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n283), .A2(new_n187), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G478), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n287), .A2(KEYINPUT15), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n286), .B(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G952), .ZN(new_n290));
  AOI211_X1 g104(.A(G953), .B(new_n290), .C1(G234), .C2(G237), .ZN(new_n291));
  INV_X1    g105(.A(new_n199), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n187), .B1(G234), .B2(G237), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT21), .B(G898), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n291), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n289), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n205), .A2(new_n207), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT19), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n235), .B(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n300), .A2(G146), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n215), .A2(new_n302), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT75), .A4(G146), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n298), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n241), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n227), .B1(new_n308), .B2(KEYINPUT90), .ZN(new_n309));
  AOI22_X1  g123(.A1(new_n234), .A2(new_n240), .B1(new_n298), .B2(new_n306), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT90), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n242), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(G475), .A2(G902), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  NOR3_X1   g129(.A1(new_n313), .A2(KEYINPUT20), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT20), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n223), .A2(new_n227), .A3(new_n241), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n226), .B1(new_n310), .B2(new_n311), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n308), .A2(KEYINPUT90), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n317), .B1(new_n321), .B2(new_n314), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n248), .B(new_n297), .C1(new_n316), .C2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT95), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT20), .B1(new_n313), .B2(new_n315), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n321), .A2(new_n317), .A3(new_n314), .ZN(new_n326));
  INV_X1    g140(.A(G475), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n234), .A2(new_n240), .ZN(new_n328));
  AOI21_X1  g142(.A(G146), .B1(new_n213), .B2(new_n214), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n329), .B1(new_n216), .B2(new_n215), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n222), .A2(new_n330), .A3(new_n218), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n198), .A2(G131), .A3(new_n202), .ZN(new_n332));
  AOI21_X1  g146(.A(G131), .B1(new_n198), .B2(new_n202), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n331), .B1(new_n334), .B2(new_n206), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n226), .B1(new_n328), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(G902), .B1(new_n336), .B2(new_n318), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n327), .B1(new_n337), .B2(KEYINPUT92), .ZN(new_n338));
  AOI22_X1  g152(.A1(new_n325), .A2(new_n326), .B1(new_n338), .B2(new_n246), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT95), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(new_n340), .A3(new_n297), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n324), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G217), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n343), .B1(G234), .B2(new_n187), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n255), .A2(KEYINPUT23), .A3(G119), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT23), .ZN(new_n346));
  INV_X1    g160(.A(G119), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n346), .B1(new_n347), .B2(G128), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n347), .A2(G128), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n345), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G110), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT72), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n352), .B1(new_n347), .B2(G128), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n255), .A2(KEYINPUT72), .A3(G119), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT73), .B1(new_n255), .B2(G119), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT73), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n357), .A2(new_n347), .A3(G128), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(KEYINPUT24), .B(G110), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n351), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n362), .B1(new_n218), .B2(new_n330), .ZN(new_n363));
  INV_X1    g177(.A(new_n361), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(new_n355), .B2(new_n359), .ZN(new_n365));
  INV_X1    g179(.A(G110), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n366), .B(new_n345), .C1(new_n348), .C2(new_n349), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n237), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(new_n305), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT78), .B1(new_n363), .B2(new_n370), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n355), .A2(new_n359), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n367), .B1(new_n372), .B2(new_n364), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n373), .A2(new_n303), .A3(new_n304), .A4(new_n237), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n364), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n220), .A2(new_n375), .A3(new_n351), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT78), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n374), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n199), .A2(G221), .A3(G234), .ZN(new_n379));
  XNOR2_X1  g193(.A(KEYINPUT22), .B(G137), .ZN(new_n380));
  OR2_X1    g194(.A1(new_n380), .A2(KEYINPUT76), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT77), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(KEYINPUT76), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n382), .B1(new_n381), .B2(new_n383), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n379), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n386), .ZN(new_n388));
  INV_X1    g202(.A(new_n379), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n389), .A3(new_n384), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n371), .A2(new_n378), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n374), .A2(new_n376), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n393), .A2(KEYINPUT78), .A3(new_n390), .A4(new_n387), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(KEYINPUT25), .B1(new_n395), .B2(new_n187), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT25), .ZN(new_n397));
  AOI211_X1 g211(.A(new_n397), .B(G902), .C1(new_n392), .C2(new_n394), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n344), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT80), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n344), .A2(G902), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n401), .B(KEYINPUT79), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n400), .B1(new_n395), .B2(new_n403), .ZN(new_n404));
  AOI211_X1 g218(.A(KEYINPUT80), .B(new_n402), .C1(new_n392), .C2(new_n394), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n399), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(G472), .A2(G902), .ZN(new_n408));
  INV_X1    g222(.A(G113), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT2), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT2), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G113), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(G116), .B(G119), .ZN(new_n414));
  OR2_X1    g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n414), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n236), .A2(G143), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n259), .A2(G146), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT1), .B1(new_n259), .B2(G146), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(G128), .A3(new_n421), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n418), .B(new_n419), .C1(KEYINPUT1), .C2(new_n255), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT65), .ZN(new_n426));
  INV_X1    g240(.A(G137), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n427), .A3(G134), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT65), .B1(new_n264), .B2(G137), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n427), .A2(G134), .ZN(new_n430));
  OAI211_X1 g244(.A(G131), .B(new_n428), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT11), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n432), .B1(new_n264), .B2(G137), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n427), .A2(KEYINPUT11), .A3(G134), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n264), .A2(G137), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n433), .A2(new_n434), .A3(new_n204), .A4(new_n435), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n431), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G131), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n436), .ZN(new_n440));
  AND2_X1   g254(.A1(KEYINPUT0), .A2(G128), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n418), .A2(new_n419), .A3(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(G143), .B(G146), .ZN(new_n443));
  XNOR2_X1  g257(.A(KEYINPUT0), .B(G128), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n425), .A2(new_n437), .B1(new_n440), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT30), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(KEYINPUT64), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT64), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n442), .B(new_n450), .C1(new_n443), .C2(new_n444), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(new_n440), .A3(new_n451), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n422), .A2(new_n431), .A3(new_n436), .A4(new_n423), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n417), .B(new_n448), .C1(new_n454), .C2(KEYINPUT30), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n440), .A2(new_n446), .ZN(new_n456));
  INV_X1    g270(.A(new_n417), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n457), .A3(new_n453), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n199), .A2(G210), .A3(new_n200), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT26), .B(G101), .ZN(new_n460));
  OR2_X1    g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n459), .A2(new_n460), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n462), .B1(new_n461), .B2(new_n463), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n455), .A2(new_n458), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT31), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT31), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n455), .A2(new_n469), .A3(new_n466), .A4(new_n458), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n452), .A2(new_n453), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT69), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n473), .A3(new_n417), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n458), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n457), .B1(new_n452), .B2(new_n453), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(new_n473), .ZN(new_n477));
  OAI21_X1  g291(.A(KEYINPUT28), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT28), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n458), .A2(KEYINPUT70), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT70), .B1(new_n458), .B2(new_n479), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n466), .B1(new_n478), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n408), .B1(new_n471), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT32), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT32), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n486), .B(new_n408), .C1(new_n471), .C2(new_n483), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n466), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT29), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n455), .A2(new_n489), .A3(new_n490), .A4(new_n458), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n187), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT71), .ZN(new_n494));
  INV_X1    g308(.A(new_n447), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n417), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n458), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n482), .A2(new_n494), .B1(KEYINPUT28), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n458), .A2(new_n479), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT70), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n458), .A2(KEYINPUT70), .A3(new_n479), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(KEYINPUT71), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n490), .B1(new_n498), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n478), .A2(new_n490), .A3(new_n482), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n466), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n493), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(G472), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n407), .B1(new_n488), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n252), .A2(G104), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT81), .ZN(new_n513));
  INV_X1    g327(.A(G104), .ZN(new_n514));
  OAI22_X1  g328(.A1(new_n513), .A2(KEYINPUT3), .B1(new_n514), .B2(G107), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n252), .A2(G104), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT3), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT81), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n513), .A2(KEYINPUT3), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR3_X1   g335(.A1(new_n516), .A2(new_n521), .A3(G101), .ZN(new_n522));
  INV_X1    g336(.A(G101), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n523), .B1(new_n512), .B2(new_n517), .ZN(new_n524));
  NOR3_X1   g338(.A1(new_n522), .A2(new_n424), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n517), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n513), .A2(KEYINPUT3), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n518), .A2(KEYINPUT81), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n511), .B1(new_n517), .B2(new_n519), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(new_n530), .A3(new_n523), .ZN(new_n531));
  INV_X1    g345(.A(new_n524), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n531), .A2(new_n532), .B1(new_n423), .B2(new_n422), .ZN(new_n533));
  OAI211_X1 g347(.A(KEYINPUT12), .B(new_n440), .C1(new_n525), .C2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT84), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n531), .A2(new_n532), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n424), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n425), .A2(new_n531), .A3(new_n532), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT84), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n539), .A2(new_n540), .A3(KEYINPUT12), .A4(new_n440), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n440), .B1(new_n525), .B2(new_n533), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT12), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n535), .A2(new_n541), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT83), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n440), .B(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n512), .B(new_n515), .C1(new_n548), .C2(new_n517), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT82), .B(KEYINPUT4), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(G101), .A3(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(KEYINPUT4), .B1(new_n549), .B2(G101), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n523), .B1(new_n529), .B2(new_n530), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n446), .B(new_n551), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT10), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n555), .B1(new_n536), .B2(new_n424), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n425), .A2(KEYINPUT10), .A3(new_n531), .A4(new_n532), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n547), .A2(new_n554), .A3(new_n556), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n199), .A2(G227), .ZN(new_n559));
  XOR2_X1   g373(.A(G110), .B(G140), .Z(new_n560));
  XOR2_X1   g374(.A(new_n559), .B(new_n560), .Z(new_n561));
  AND2_X1   g375(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n545), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n554), .A2(new_n556), .A3(new_n557), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n440), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n558), .ZN(new_n566));
  INV_X1    g380(.A(new_n561), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n563), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(G469), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(new_n570), .A3(new_n187), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n545), .A2(new_n558), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n567), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n562), .A2(new_n565), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(G469), .A3(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n570), .A2(new_n187), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n571), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(G221), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n579), .B1(new_n279), .B2(new_n187), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(G214), .B1(G237), .B2(G902), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n445), .A2(G125), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(G125), .B1(new_n422), .B2(new_n423), .ZN(new_n586));
  OAI21_X1  g400(.A(KEYINPUT87), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(G224), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(G953), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT87), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n584), .A2(new_n591), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n587), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n590), .B1(new_n587), .B2(new_n592), .ZN(new_n594));
  OR2_X1    g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n417), .B(new_n551), .C1(new_n552), .C2(new_n553), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n267), .A2(G119), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT5), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n409), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n347), .A2(G116), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n267), .A2(G119), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n601), .A3(KEYINPUT5), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n599), .A2(new_n602), .B1(new_n414), .B2(new_n413), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n531), .A2(new_n603), .A3(new_n532), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(KEYINPUT85), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT85), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n531), .A2(new_n603), .A3(new_n532), .A4(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(G110), .B(G122), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n596), .A2(new_n605), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n596), .A2(new_n605), .A3(new_n607), .ZN(new_n610));
  INV_X1    g424(.A(new_n608), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n611), .A2(KEYINPUT86), .ZN(new_n612));
  AOI22_X1  g426(.A1(KEYINPUT6), .A2(new_n609), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n610), .A2(KEYINPUT6), .A3(new_n612), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n595), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n587), .A2(KEYINPUT7), .A3(new_n590), .A4(new_n592), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n608), .B(KEYINPUT8), .ZN(new_n617));
  INV_X1    g431(.A(new_n604), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n603), .B1(new_n531), .B2(new_n532), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n590), .A2(KEYINPUT7), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n621), .B1(new_n585), .B2(new_n586), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n616), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(G902), .B1(new_n623), .B2(new_n609), .ZN(new_n624));
  OAI21_X1  g438(.A(G210), .B1(G237), .B2(G902), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n615), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n625), .B1(new_n615), .B2(new_n624), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n583), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n582), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n342), .A2(new_n510), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(G101), .ZN(G3));
  OAI21_X1  g446(.A(new_n187), .B1(new_n471), .B2(new_n483), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(G472), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n484), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(new_n407), .ZN(new_n636));
  INV_X1    g450(.A(new_n582), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n583), .ZN(new_n640));
  INV_X1    g454(.A(new_n625), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n593), .A2(new_n594), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n609), .A2(KEYINPUT6), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n610), .A2(new_n612), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n610), .A2(KEYINPUT6), .A3(new_n612), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n642), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n616), .A2(new_n620), .A3(new_n622), .ZN(new_n648));
  INV_X1    g462(.A(new_n609), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n187), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n641), .B1(new_n647), .B2(new_n650), .ZN(new_n651));
  AOI211_X1 g465(.A(new_n296), .B(new_n640), .C1(new_n651), .C2(new_n626), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n639), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n248), .B1(new_n316), .B2(new_n322), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n280), .A2(KEYINPUT96), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n277), .B(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT33), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(KEYINPUT33), .B1(new_n283), .B2(new_n285), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n287), .A2(G902), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(KEYINPUT97), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT97), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n664), .B(new_n661), .C1(new_n658), .C2(new_n659), .ZN(new_n665));
  INV_X1    g479(.A(new_n286), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n663), .B(new_n665), .C1(G478), .C2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n654), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n653), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT34), .B(G104), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G6));
  NAND2_X1  g485(.A1(new_n248), .A2(new_n289), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT98), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n673), .B1(new_n316), .B2(new_n322), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n325), .A2(KEYINPUT98), .A3(new_n326), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n672), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n639), .A2(new_n652), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n677), .B(KEYINPUT99), .Z(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT35), .B(G107), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G9));
  NOR2_X1   g494(.A1(new_n391), .A2(KEYINPUT36), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(new_n393), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n403), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n399), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n635), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n342), .A2(new_n630), .A3(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT37), .B(G110), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G12));
  AOI21_X1  g502(.A(new_n684), .B1(new_n488), .B2(new_n509), .ZN(new_n689));
  INV_X1    g503(.A(new_n291), .ZN(new_n690));
  INV_X1    g504(.A(new_n294), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n690), .B1(new_n691), .B2(G900), .ZN(new_n692));
  XOR2_X1   g506(.A(new_n692), .B(KEYINPUT100), .Z(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n689), .A2(new_n676), .A3(new_n630), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G128), .ZN(G30));
  XOR2_X1   g510(.A(new_n693), .B(KEYINPUT39), .Z(new_n697));
  NAND2_X1  g511(.A1(new_n637), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(new_n698), .B(KEYINPUT101), .Z(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT40), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n698), .B(KEYINPUT101), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT40), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n627), .A2(new_n628), .ZN(new_n704));
  XOR2_X1   g518(.A(new_n704), .B(KEYINPUT38), .Z(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n654), .A3(new_n289), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n399), .A2(new_n683), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n455), .A2(new_n458), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n708), .A2(new_n489), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n187), .B1(new_n497), .B2(new_n466), .ZN(new_n710));
  OAI21_X1  g524(.A(G472), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n488), .A2(new_n711), .ZN(new_n712));
  NOR4_X1   g526(.A1(new_n706), .A2(new_n640), .A3(new_n707), .A4(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n700), .A2(new_n703), .A3(new_n713), .ZN(new_n714));
  XOR2_X1   g528(.A(KEYINPUT102), .B(G143), .Z(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G45));
  OAI21_X1  g530(.A(new_n665), .B1(new_n666), .B2(G478), .ZN(new_n717));
  OR2_X1    g531(.A1(new_n656), .A2(new_n657), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n283), .A2(new_n285), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n657), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n664), .B1(new_n721), .B2(new_n661), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n717), .A2(new_n722), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n339), .A2(new_n723), .A3(new_n693), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n689), .A2(new_n630), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G146), .ZN(G48));
  INV_X1    g540(.A(new_n668), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n652), .ZN(new_n728));
  INV_X1    g542(.A(new_n487), .ZN(new_n729));
  AOI22_X1  g543(.A1(new_n476), .A2(new_n473), .B1(new_n457), .B2(new_n447), .ZN(new_n730));
  OAI21_X1  g544(.A(KEYINPUT69), .B1(new_n454), .B2(new_n457), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n503), .B1(new_n732), .B2(KEYINPUT28), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n468), .B(new_n470), .C1(new_n733), .C2(new_n466), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n486), .B1(new_n734), .B2(new_n408), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n482), .A2(new_n494), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n497), .A2(KEYINPUT28), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n736), .A2(new_n504), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT29), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n489), .B1(new_n733), .B2(new_n490), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n492), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(G472), .ZN(new_n742));
  OAI22_X1  g556(.A1(new_n729), .A2(new_n735), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n407), .ZN(new_n744));
  AOI22_X1  g558(.A1(new_n545), .A2(new_n562), .B1(new_n566), .B2(new_n567), .ZN(new_n745));
  OAI21_X1  g559(.A(G469), .B1(new_n745), .B2(G902), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n571), .A3(new_n581), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n743), .A2(new_n744), .A3(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n728), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(KEYINPUT41), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(new_n409), .ZN(G15));
  INV_X1    g566(.A(new_n289), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n753), .B1(new_n246), .B2(new_n338), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n325), .A2(KEYINPUT98), .A3(new_n326), .ZN(new_n755));
  AOI21_X1  g569(.A(KEYINPUT98), .B1(new_n325), .B2(new_n326), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n754), .B(new_n652), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n749), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(new_n267), .ZN(G18));
  NOR2_X1   g573(.A1(new_n629), .A2(new_n747), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n342), .A2(new_n689), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT103), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n743), .A2(new_n760), .A3(new_n707), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT103), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n764), .A3(new_n342), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G119), .ZN(G21));
  INV_X1    g581(.A(new_n408), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n738), .A2(new_n489), .ZN(new_n769));
  INV_X1    g583(.A(new_n471), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  XOR2_X1   g585(.A(KEYINPUT104), .B(G472), .Z(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n773), .B1(new_n734), .B2(new_n187), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n407), .A2(new_n771), .A3(new_n774), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n629), .A2(new_n747), .A3(new_n296), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT105), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n777), .B1(new_n339), .B2(new_n753), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n654), .A2(KEYINPUT105), .A3(new_n289), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n775), .A2(new_n776), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  XOR2_X1   g594(.A(KEYINPUT106), .B(G122), .Z(new_n781));
  XNOR2_X1  g595(.A(new_n780), .B(new_n781), .ZN(G24));
  NAND2_X1  g596(.A1(new_n769), .A2(new_n770), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n408), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n633), .A2(new_n772), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n784), .A2(new_n707), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(new_n724), .A3(new_n760), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G125), .ZN(G27));
  AND3_X1   g602(.A1(new_n651), .A2(new_n583), .A3(new_n626), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n789), .A2(new_n581), .A3(new_n578), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n724), .A2(new_n790), .A3(new_n743), .A4(new_n744), .ZN(new_n791));
  XNOR2_X1  g605(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT108), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n510), .A2(KEYINPUT42), .A3(new_n724), .A4(new_n790), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n794), .B1(new_n793), .B2(new_n795), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XOR2_X1   g612(.A(KEYINPUT109), .B(G131), .Z(new_n799));
  XNOR2_X1  g613(.A(new_n798), .B(new_n799), .ZN(G33));
  AOI211_X1 g614(.A(new_n693), .B(new_n672), .C1(new_n674), .C2(new_n675), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n801), .A2(new_n510), .A3(new_n790), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G134), .ZN(G36));
  AOI22_X1  g617(.A1(new_n572), .A2(new_n567), .B1(new_n565), .B2(new_n562), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n804), .A2(KEYINPUT45), .ZN(new_n805));
  OAI21_X1  g619(.A(G469), .B1(new_n804), .B2(KEYINPUT45), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n577), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT46), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n807), .A2(KEYINPUT46), .A3(new_n577), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(new_n571), .A3(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n812), .A2(new_n581), .A3(new_n697), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n339), .B(KEYINPUT110), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT43), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n723), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n815), .B1(new_n654), .B2(new_n723), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(new_n635), .A3(new_n707), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT44), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n813), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n822), .B(new_n789), .C1(new_n821), .C2(new_n820), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(G137), .ZN(G39));
  INV_X1    g638(.A(new_n789), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n743), .A2(new_n825), .A3(new_n744), .ZN(new_n826));
  XNOR2_X1  g640(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n812), .A2(new_n581), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n827), .B1(new_n812), .B2(new_n581), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n724), .B(new_n826), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(G140), .ZN(G42));
  NAND2_X1  g645(.A1(new_n290), .A2(new_n191), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n690), .B1(new_n817), .B2(new_n818), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n835), .A2(new_n775), .A3(new_n789), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n828), .A2(new_n829), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n746), .A2(new_n571), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n580), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n705), .A2(new_n583), .A3(new_n747), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n835), .A2(KEYINPUT50), .A3(new_n775), .A4(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n834), .B1(new_n819), .B2(new_n291), .ZN(new_n844));
  AOI211_X1 g658(.A(KEYINPUT116), .B(new_n690), .C1(new_n817), .C2(new_n818), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n775), .B(new_n842), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT50), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n825), .A2(new_n747), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n835), .A2(KEYINPUT117), .A3(new_n786), .A4(new_n850), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n786), .B(new_n850), .C1(new_n844), .C2(new_n845), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT117), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n712), .A2(new_n850), .A3(new_n744), .A4(new_n291), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(new_n339), .A3(new_n723), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n849), .A2(new_n855), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n841), .B1(new_n859), .B2(KEYINPUT118), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n849), .A2(new_n855), .A3(new_n858), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT51), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n835), .A2(new_n510), .A3(new_n850), .ZN(new_n865));
  XNOR2_X1  g679(.A(KEYINPUT120), .B(KEYINPUT48), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT48), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(KEYINPUT120), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n835), .A2(new_n510), .A3(new_n850), .A4(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n835), .A2(new_n760), .A3(new_n775), .ZN(new_n871));
  AOI211_X1 g685(.A(new_n290), .B(G953), .C1(new_n857), .C2(new_n727), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n867), .A2(new_n870), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT51), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n875), .B1(new_n837), .B2(new_n839), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n836), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n840), .A2(new_n875), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n874), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n873), .B1(new_n859), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n399), .A2(new_n683), .A3(new_n694), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n881), .B1(new_n488), .B2(new_n711), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n882), .A2(new_n630), .A3(new_n778), .A4(new_n779), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n695), .A2(new_n883), .A3(new_n725), .A4(new_n787), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT114), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n630), .B(new_n689), .C1(new_n801), .C2(new_n724), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT114), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n886), .A2(new_n887), .A3(new_n787), .A4(new_n883), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT52), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n761), .A2(KEYINPUT103), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n764), .B1(new_n763), .B2(new_n342), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI211_X1 g708(.A(new_n407), .B(new_n747), .C1(new_n488), .C2(new_n509), .ZN(new_n895));
  INV_X1    g709(.A(new_n757), .ZN(new_n896));
  INV_X1    g710(.A(new_n652), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n668), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n895), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n342), .B(new_n630), .C1(new_n510), .C2(new_n685), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n339), .A2(new_n289), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n636), .A2(new_n902), .A3(new_n637), .A4(new_n652), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n899), .A2(new_n900), .A3(new_n780), .A4(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT113), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT112), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n906), .B1(new_n339), .B2(new_n723), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n654), .A2(new_n667), .A3(KEYINPUT112), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n905), .B1(new_n909), .B2(new_n897), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n907), .A2(new_n908), .A3(KEYINPUT113), .A4(new_n652), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n638), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n894), .A2(new_n904), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n248), .A2(new_n753), .A3(new_n694), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n914), .B1(new_n674), .B2(new_n675), .ZN(new_n915));
  AOI22_X1  g729(.A1(new_n689), .A2(new_n915), .B1(new_n786), .B2(new_n724), .ZN(new_n916));
  INV_X1    g730(.A(new_n790), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n802), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n796), .A2(new_n797), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n885), .A2(KEYINPUT52), .A3(new_n888), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n891), .A2(new_n913), .A3(new_n919), .A4(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT53), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n913), .A2(new_n919), .A3(new_n922), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n884), .A2(KEYINPUT52), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n889), .B2(new_n890), .ZN(new_n925));
  AOI22_X1  g739(.A1(KEYINPUT53), .A2(new_n921), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(KEYINPUT54), .ZN(new_n927));
  XNOR2_X1  g741(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n910), .A2(new_n911), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n639), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n903), .A2(new_n780), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n749), .B1(new_n728), .B2(new_n757), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n931), .A2(new_n934), .A3(new_n766), .A4(new_n900), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n922), .B1(new_n793), .B2(new_n795), .ZN(new_n936));
  OR2_X1    g750(.A1(new_n916), .A2(new_n917), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n936), .A2(new_n937), .A3(new_n802), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  AOI221_X4 g753(.A(new_n929), .B1(new_n925), .B2(new_n939), .C1(new_n921), .C2(new_n922), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n880), .A2(new_n927), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n832), .B1(new_n864), .B2(new_n942), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n838), .B(KEYINPUT49), .Z(new_n944));
  NAND3_X1  g758(.A1(new_n667), .A2(new_n583), .A3(new_n581), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n944), .A2(new_n407), .A3(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n705), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n946), .A2(new_n712), .A3(new_n947), .A4(new_n814), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n943), .A2(new_n948), .ZN(G75));
  NAND2_X1  g763(.A1(new_n292), .A2(new_n290), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT122), .Z(new_n951));
  NAND3_X1  g765(.A1(new_n913), .A2(new_n919), .A3(new_n920), .ZN(new_n952));
  AOI21_X1  g766(.A(KEYINPUT52), .B1(new_n885), .B2(new_n888), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n922), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n925), .A2(new_n939), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(G902), .ZN(new_n957));
  INV_X1    g771(.A(G210), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n645), .A2(new_n646), .A3(new_n642), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n615), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT55), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n962), .A2(KEYINPUT56), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n951), .B1(new_n959), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n959), .A2(KEYINPUT121), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT56), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT121), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(new_n957), .B2(new_n958), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n965), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n964), .B1(new_n969), .B2(new_n962), .ZN(G51));
  INV_X1    g784(.A(new_n951), .ZN(new_n971));
  XNOR2_X1  g785(.A(KEYINPUT123), .B(KEYINPUT57), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(new_n576), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n928), .B1(new_n954), .B2(new_n955), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n973), .B1(new_n940), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(KEYINPUT124), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT124), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n977), .B(new_n973), .C1(new_n940), .C2(new_n974), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n976), .A2(new_n569), .A3(new_n978), .ZN(new_n979));
  OR2_X1    g793(.A1(new_n957), .A2(new_n807), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n971), .B1(new_n979), .B2(new_n980), .ZN(G54));
  INV_X1    g795(.A(KEYINPUT58), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n957), .A2(new_n982), .A3(new_n327), .ZN(new_n983));
  OR2_X1    g797(.A1(new_n983), .A2(new_n313), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n313), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n971), .B1(new_n984), .B2(new_n985), .ZN(G60));
  NAND2_X1  g800(.A1(G478), .A2(G902), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT59), .Z(new_n988));
  AOI21_X1  g802(.A(new_n988), .B1(new_n941), .B2(new_n927), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n989), .A2(new_n721), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n940), .A2(new_n974), .ZN(new_n991));
  OR2_X1    g805(.A1(new_n660), .A2(new_n988), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n951), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n990), .A2(new_n993), .ZN(G63));
  NAND2_X1  g808(.A1(G217), .A2(G902), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(KEYINPUT60), .Z(new_n996));
  NAND2_X1  g810(.A1(new_n956), .A2(new_n996), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n395), .B(KEYINPUT126), .Z(new_n998));
  AOI21_X1  g812(.A(new_n971), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(KEYINPUT61), .B1(new_n999), .B2(KEYINPUT125), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n956), .A2(new_n682), .A3(new_n996), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g817(.A(new_n999), .B(new_n1001), .C1(KEYINPUT125), .C2(KEYINPUT61), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(new_n1004), .ZN(G66));
  OAI21_X1  g819(.A(G953), .B1(new_n295), .B2(new_n588), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1006), .B1(new_n913), .B2(new_n292), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n645), .B(new_n646), .C1(G898), .C2(new_n199), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1007), .B(new_n1008), .ZN(G69));
  NAND3_X1  g823(.A1(new_n714), .A2(new_n787), .A3(new_n886), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1010), .B(KEYINPUT62), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n909), .A2(new_n901), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n1012), .A2(KEYINPUT127), .ZN(new_n1013));
  AND3_X1   g827(.A1(new_n701), .A2(new_n510), .A3(new_n789), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1012), .A2(KEYINPUT127), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n823), .B(new_n830), .C1(new_n1013), .C2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n199), .B1(new_n1011), .B2(new_n1017), .ZN(new_n1018));
  MUX2_X1   g832(.A(new_n454), .B(new_n495), .S(KEYINPUT30), .Z(new_n1019));
  XOR2_X1   g833(.A(new_n1019), .B(new_n300), .Z(new_n1020));
  INV_X1    g834(.A(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n292), .A2(G900), .ZN(new_n1023));
  INV_X1    g837(.A(new_n510), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n778), .A2(new_n779), .ZN(new_n1025));
  NOR4_X1   g839(.A1(new_n813), .A2(new_n1024), .A3(new_n629), .A4(new_n1025), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n886), .A2(new_n787), .A3(new_n802), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g842(.A1(new_n823), .A2(new_n1028), .A3(new_n798), .A4(new_n830), .ZN(new_n1029));
  OAI211_X1 g843(.A(new_n1020), .B(new_n1023), .C1(new_n1029), .C2(new_n292), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1022), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n199), .B1(G227), .B2(G900), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g847(.A(new_n1032), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n1022), .A2(new_n1034), .A3(new_n1030), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1033), .A2(new_n1035), .ZN(G72));
  NOR3_X1   g850(.A1(new_n1011), .A2(new_n935), .A3(new_n1017), .ZN(new_n1037));
  NAND2_X1  g851(.A1(G472), .A2(G902), .ZN(new_n1038));
  XOR2_X1   g852(.A(new_n1038), .B(KEYINPUT63), .Z(new_n1039));
  INV_X1    g853(.A(new_n1039), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n709), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n1039), .B1(new_n1029), .B2(new_n935), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n708), .A2(new_n489), .ZN(new_n1043));
  INV_X1    g857(.A(new_n1043), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n971), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1041), .A2(new_n1045), .ZN(new_n1046));
  NOR3_X1   g860(.A1(new_n1044), .A2(new_n709), .A3(new_n1040), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n1046), .B1(new_n926), .B2(new_n1047), .ZN(G57));
endmodule


