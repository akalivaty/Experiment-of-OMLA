//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 1 1 0 0 1 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n981, new_n982, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(new_n187), .B(KEYINPUT84), .Z(new_n188));
  OAI21_X1  g002(.A(G210), .B1(G237), .B2(G902), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT88), .ZN(new_n190));
  XNOR2_X1  g004(.A(G110), .B(G122), .ZN(new_n191));
  XOR2_X1   g005(.A(new_n191), .B(KEYINPUT85), .Z(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT68), .ZN(new_n194));
  INV_X1    g008(.A(G116), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT68), .A2(G116), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(G119), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G113), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT2), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G113), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n195), .A2(G119), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n198), .A2(new_n203), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT69), .ZN(new_n208));
  AND2_X1   g022(.A1(KEYINPUT68), .A2(G116), .ZN(new_n209));
  NOR2_X1   g023(.A1(KEYINPUT68), .A2(G116), .ZN(new_n210));
  INV_X1    g024(.A(G119), .ZN(new_n211));
  NOR3_X1   g025(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n208), .B1(new_n212), .B2(new_n204), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n198), .A2(KEYINPUT69), .A3(new_n205), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n203), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT70), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n207), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n203), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n198), .A2(KEYINPUT69), .A3(new_n205), .ZN(new_n219));
  AOI21_X1  g033(.A(KEYINPUT69), .B1(new_n198), .B2(new_n205), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT70), .ZN(new_n222));
  INV_X1    g036(.A(G101), .ZN(new_n223));
  INV_X1    g037(.A(G104), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT3), .B1(new_n224), .B2(G107), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n226));
  INV_X1    g040(.A(G107), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n226), .A2(new_n227), .A3(G104), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n224), .A2(G107), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n225), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT80), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n223), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n225), .A2(new_n228), .A3(KEYINPUT80), .A4(new_n229), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n225), .A2(new_n228), .A3(new_n223), .A4(new_n229), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n232), .A2(new_n233), .B1(KEYINPUT4), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n232), .A2(KEYINPUT4), .A3(new_n233), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n217), .A2(new_n222), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n213), .A2(KEYINPUT5), .A3(new_n214), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT5), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n199), .B1(new_n204), .B2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n207), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n224), .A2(G107), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n227), .A2(G104), .ZN(new_n244));
  OAI21_X1  g058(.A(G101), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT81), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n234), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n246), .B1(new_n234), .B2(new_n245), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n242), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n193), .B1(new_n238), .B2(new_n251), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n216), .B(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n222), .A2(new_n206), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n236), .A2(new_n237), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(new_n250), .A3(new_n192), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n252), .A2(new_n257), .A3(KEYINPUT6), .ZN(new_n258));
  INV_X1    g072(.A(G128), .ZN(new_n259));
  INV_X1    g073(.A(G146), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G143), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n259), .B1(new_n261), .B2(KEYINPUT1), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G143), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT65), .B1(new_n264), .B2(G146), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT65), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(new_n260), .A3(G143), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(KEYINPUT66), .B1(new_n260), .B2(G143), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT66), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(new_n264), .A3(G146), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n263), .B1(new_n268), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT1), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n264), .A2(G146), .ZN(new_n275));
  AND4_X1   g089(.A1(new_n274), .A2(new_n275), .A3(new_n261), .A4(G128), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(KEYINPUT78), .B(G125), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AND4_X1   g094(.A1(KEYINPUT0), .A2(new_n275), .A3(new_n261), .A4(G128), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n269), .A2(new_n271), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n265), .A2(new_n267), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(KEYINPUT0), .B(G128), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n281), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n279), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n280), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G953), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(G224), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n290), .B(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT6), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n294), .B(new_n193), .C1(new_n238), .C2(new_n251), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n258), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G902), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT87), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n192), .B(KEYINPUT8), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n234), .A2(new_n245), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n239), .A2(new_n241), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n300), .B1(new_n301), .B2(new_n206), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n198), .A2(KEYINPUT5), .A3(new_n205), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n303), .A2(new_n241), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n206), .A2(new_n234), .A3(new_n245), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT86), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n303), .A2(new_n241), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT86), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n300), .A2(new_n307), .A3(new_n308), .A4(new_n206), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n298), .B(new_n299), .C1(new_n302), .C2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n309), .B(new_n306), .C1(new_n242), .C2(new_n300), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n298), .B1(new_n313), .B2(new_n299), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n292), .A2(KEYINPUT7), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n290), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n280), .A2(new_n289), .A3(new_n316), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n257), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n297), .B1(new_n315), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n190), .B1(new_n296), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n313), .A2(new_n299), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT87), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n311), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n318), .A2(new_n319), .ZN(new_n326));
  AOI22_X1  g140(.A1(new_n254), .A2(new_n255), .B1(new_n249), .B2(new_n242), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n326), .B1(new_n327), .B2(new_n192), .ZN(new_n328));
  AOI21_X1  g142(.A(G902), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n258), .A2(new_n293), .A3(new_n295), .ZN(new_n330));
  INV_X1    g144(.A(new_n190), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n188), .B1(new_n322), .B2(new_n332), .ZN(new_n333));
  XOR2_X1   g147(.A(KEYINPUT77), .B(G902), .Z(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT9), .B(G234), .ZN(new_n335));
  INV_X1    g149(.A(G217), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n335), .A2(new_n336), .A3(G953), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n264), .A2(G128), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n259), .A2(G143), .ZN(new_n339));
  INV_X1    g153(.A(G134), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n195), .A2(G122), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n209), .A2(new_n210), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n343), .B1(new_n344), .B2(G122), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n227), .ZN(new_n346));
  AND3_X1   g160(.A1(new_n196), .A2(G122), .A3(new_n197), .ZN(new_n347));
  OAI21_X1  g161(.A(G107), .B1(new_n347), .B2(new_n343), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n342), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT90), .B(KEYINPUT13), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n339), .B1(new_n350), .B2(new_n338), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n338), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT91), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT91), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n350), .A2(new_n354), .A3(new_n338), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n351), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n349), .B1(new_n340), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT92), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT14), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n345), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n196), .A2(KEYINPUT14), .A3(G122), .A4(new_n197), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(G107), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n338), .A2(new_n339), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G134), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n341), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n362), .A2(KEYINPUT93), .A3(new_n346), .A4(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT93), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n346), .A2(new_n365), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n361), .A2(G107), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n369), .B1(new_n359), .B2(new_n345), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n367), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n357), .A2(new_n358), .B1(new_n366), .B2(new_n371), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n349), .B(KEYINPUT92), .C1(new_n340), .C2(new_n356), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n337), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n357), .A2(new_n358), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n366), .A2(new_n371), .ZN(new_n376));
  AND4_X1   g190(.A1(new_n373), .A2(new_n375), .A3(new_n376), .A4(new_n337), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n334), .B1(new_n374), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G478), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n379), .A2(KEYINPUT15), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n375), .A2(new_n376), .A3(new_n373), .ZN(new_n382));
  INV_X1    g196(.A(new_n337), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n372), .A2(new_n373), .A3(new_n337), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n380), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n334), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n381), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT16), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT78), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(G125), .ZN(new_n392));
  INV_X1    g206(.A(G125), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n393), .A2(KEYINPUT78), .ZN(new_n394));
  OAI21_X1  g208(.A(G140), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(G125), .A2(G140), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n390), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G140), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n390), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n393), .A2(KEYINPUT78), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n391), .A2(G125), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n260), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n399), .B1(new_n401), .B2(new_n402), .ZN(new_n405));
  OAI21_X1  g219(.A(KEYINPUT16), .B1(new_n405), .B2(new_n396), .ZN(new_n406));
  INV_X1    g220(.A(new_n403), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(G146), .A3(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(G237), .A2(G953), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(G143), .A3(G214), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(G143), .B1(new_n409), .B2(G214), .ZN(new_n412));
  OAI21_X1  g226(.A(G131), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n412), .ZN(new_n414));
  INV_X1    g228(.A(G131), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n415), .A3(new_n410), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT17), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n413), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n414), .A2(new_n410), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(KEYINPUT17), .A3(G131), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n404), .A2(new_n408), .A3(new_n418), .A4(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(G113), .B(G122), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n422), .B(new_n224), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT89), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n419), .A2(new_n424), .A3(KEYINPUT18), .A4(G131), .ZN(new_n425));
  XNOR2_X1  g239(.A(G125), .B(G140), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n260), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n397), .B1(new_n279), .B2(new_n399), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n427), .B1(new_n428), .B2(new_n260), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n424), .A2(KEYINPUT18), .A3(G131), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n414), .A2(new_n410), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n425), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n421), .A2(new_n423), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n413), .A2(new_n416), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n426), .A2(KEYINPUT19), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n435), .B1(new_n428), .B2(KEYINPUT19), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n408), .B(new_n434), .C1(G146), .C2(new_n436), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n437), .A2(new_n432), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n433), .B1(new_n438), .B2(new_n423), .ZN(new_n439));
  NOR2_X1   g253(.A1(G475), .A2(G902), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT20), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT20), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n439), .A2(new_n443), .A3(new_n440), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n421), .A2(new_n423), .A3(new_n432), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n423), .B1(new_n421), .B2(new_n432), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n297), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(G475), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(G952), .ZN(new_n451));
  AOI211_X1 g265(.A(G953), .B(new_n451), .C1(G234), .C2(G237), .ZN(new_n452));
  AOI211_X1 g266(.A(new_n291), .B(new_n334), .C1(G234), .C2(G237), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(G898), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n389), .A2(new_n450), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT83), .ZN(new_n457));
  INV_X1    g271(.A(G221), .ZN(new_n458));
  INV_X1    g272(.A(new_n335), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n458), .B1(new_n459), .B2(new_n297), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT71), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n285), .B1(new_n282), .B2(new_n283), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n462), .B1(new_n463), .B2(new_n281), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n286), .B1(new_n268), .B2(new_n272), .ZN(new_n465));
  INV_X1    g279(.A(new_n281), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(KEYINPUT71), .A3(new_n466), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n232), .A2(KEYINPUT4), .A3(new_n233), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n464), .B(new_n467), .C1(new_n468), .C2(new_n235), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT10), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n470), .B1(new_n273), .B2(new_n277), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n275), .A2(new_n261), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n472), .A2(new_n262), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n234), .B(new_n245), .C1(new_n473), .C2(new_n276), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n249), .A2(new_n471), .B1(new_n474), .B2(new_n470), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT67), .B1(new_n340), .B2(G137), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT11), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT11), .ZN(new_n478));
  OAI211_X1 g292(.A(KEYINPUT67), .B(new_n478), .C1(new_n340), .C2(G137), .ZN(new_n479));
  INV_X1    g293(.A(G137), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n480), .A2(G134), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n477), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(G131), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n477), .A2(new_n415), .A3(new_n479), .A4(new_n482), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n469), .A2(new_n475), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n474), .B1(new_n278), .B2(new_n300), .ZN(new_n489));
  AOI21_X1  g303(.A(KEYINPUT82), .B1(new_n484), .B2(new_n485), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(KEYINPUT12), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT12), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n489), .A2(new_n493), .A3(new_n490), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n488), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(G110), .B(G140), .ZN(new_n496));
  INV_X1    g310(.A(G227), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n497), .A2(G953), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n496), .B(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n469), .A2(new_n475), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n486), .ZN(new_n502));
  INV_X1    g316(.A(new_n499), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n488), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n500), .A2(G469), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(G469), .A2(G902), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n334), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n469), .A2(new_n475), .A3(new_n487), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n487), .B1(new_n469), .B2(new_n475), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n499), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n488), .A2(new_n492), .A3(new_n503), .A4(new_n494), .ZN(new_n512));
  AOI211_X1 g326(.A(G469), .B(new_n508), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n457), .B(new_n461), .C1(new_n507), .C2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(G469), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n503), .B1(new_n502), .B2(new_n488), .ZN(new_n517));
  AND4_X1   g331(.A1(new_n488), .A2(new_n492), .A3(new_n503), .A4(new_n494), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n516), .B(new_n334), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(new_n506), .A3(new_n505), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n457), .B1(new_n520), .B2(new_n461), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n333), .B(new_n456), .C1(new_n515), .C2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT94), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n461), .B1(new_n507), .B2(new_n513), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT83), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n514), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n527), .A2(KEYINPUT94), .A3(new_n333), .A4(new_n456), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n464), .A2(new_n486), .A3(new_n467), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n340), .A2(G137), .ZN(new_n530));
  OAI21_X1  g344(.A(G131), .B1(new_n530), .B2(new_n481), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n262), .B1(new_n282), .B2(new_n283), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n485), .B(new_n531), .C1(new_n532), .C2(new_n276), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT72), .B1(new_n534), .B2(new_n254), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n253), .A2(new_n206), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n213), .A2(new_n214), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n216), .B1(new_n537), .B2(new_n218), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT72), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n539), .A2(new_n540), .A3(new_n529), .A4(new_n533), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n534), .A2(new_n254), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n535), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT28), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT28), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(new_n534), .B2(new_n254), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n409), .A2(G210), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n547), .B(KEYINPUT27), .ZN(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT26), .B(G101), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n548), .B(new_n549), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n550), .A2(KEYINPUT29), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n544), .A2(new_n546), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT76), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT76), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n544), .A2(new_n554), .A3(new_n546), .A4(new_n551), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n535), .A2(new_n541), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT75), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n485), .A2(new_n531), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n287), .A2(new_n486), .B1(new_n278), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n558), .B1(new_n539), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n485), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n481), .B1(new_n476), .B2(KEYINPUT11), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n415), .B1(new_n563), .B2(new_n479), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n465), .B(new_n466), .C1(new_n562), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n533), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n254), .A2(KEYINPUT75), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n561), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(KEYINPUT28), .B1(new_n557), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(new_n546), .A3(new_n550), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n529), .A2(KEYINPUT30), .A3(new_n533), .ZN(new_n571));
  XOR2_X1   g385(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n572));
  NAND2_X1  g386(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n571), .A2(new_n573), .A3(new_n254), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n574), .A2(new_n535), .A3(new_n541), .ZN(new_n575));
  INV_X1    g389(.A(new_n550), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT29), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n508), .B1(new_n570), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n556), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(G472), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT32), .ZN(new_n581));
  AND4_X1   g395(.A1(new_n535), .A2(new_n574), .A3(new_n541), .A4(new_n550), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT74), .ZN(new_n583));
  XOR2_X1   g397(.A(KEYINPUT73), .B(KEYINPUT31), .Z(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n582), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n574), .A2(new_n535), .A3(new_n541), .A4(new_n550), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n587), .A2(KEYINPUT31), .ZN(new_n588));
  OAI21_X1  g402(.A(KEYINPUT74), .B1(new_n587), .B2(new_n584), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n586), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n569), .A2(new_n546), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n576), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(G472), .A2(G902), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n581), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n594), .ZN(new_n596));
  AOI211_X1 g410(.A(KEYINPUT32), .B(new_n596), .C1(new_n590), .C2(new_n592), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n580), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n336), .B1(new_n334), .B2(G234), .ZN(new_n599));
  XNOR2_X1  g413(.A(KEYINPUT22), .B(G137), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n291), .A2(G221), .A3(G234), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT79), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n259), .A2(G119), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT23), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n211), .A2(G128), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n259), .A2(KEYINPUT23), .A3(G119), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(G110), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n608), .A2(new_n605), .ZN(new_n612));
  XNOR2_X1  g426(.A(KEYINPUT24), .B(G110), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n404), .B2(new_n408), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n612), .A2(new_n613), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n616), .B1(G110), .B2(new_n610), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n408), .A2(new_n427), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n604), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n612), .A2(new_n613), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(G110), .B2(new_n610), .ZN(new_n621));
  AOI211_X1 g435(.A(new_n260), .B(new_n403), .C1(new_n428), .C2(KEYINPUT16), .ZN(new_n622));
  AOI21_X1  g436(.A(G146), .B1(new_n406), .B2(new_n407), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n408), .A2(new_n427), .A3(new_n617), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(KEYINPUT79), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n603), .B1(new_n619), .B2(new_n626), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n626), .A2(new_n603), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(KEYINPUT25), .B1(new_n629), .B2(new_n334), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT25), .ZN(new_n631));
  NOR4_X1   g445(.A1(new_n627), .A2(new_n628), .A3(new_n631), .A4(new_n508), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n599), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n599), .A2(G902), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n629), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n524), .A2(new_n528), .A3(new_n598), .A4(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G101), .ZN(G3));
  AOI21_X1  g453(.A(new_n508), .B1(new_n590), .B2(new_n592), .ZN(new_n640));
  INV_X1    g454(.A(G472), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n550), .B1(new_n569), .B2(new_n546), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n587), .A2(KEYINPUT31), .ZN(new_n643));
  OAI211_X1 g457(.A(new_n643), .B(KEYINPUT74), .C1(new_n587), .C2(new_n584), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n642), .B1(new_n644), .B2(new_n586), .ZN(new_n645));
  OAI22_X1  g459(.A1(new_n640), .A2(new_n641), .B1(new_n645), .B2(new_n596), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n322), .A2(new_n332), .ZN(new_n648));
  INV_X1    g462(.A(new_n188), .ZN(new_n649));
  INV_X1    g463(.A(new_n455), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n508), .A2(new_n379), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT33), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n384), .A2(new_n385), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n653), .B1(new_n384), .B2(new_n385), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n652), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(G478), .B1(new_n386), .B2(new_n334), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n450), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n651), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n636), .B1(new_n526), .B2(new_n514), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n647), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT34), .B(G104), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT95), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n663), .B(new_n665), .ZN(G6));
  NAND2_X1  g480(.A1(new_n449), .A2(KEYINPUT96), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT96), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n448), .A2(new_n668), .A3(G475), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n445), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n389), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n651), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n647), .A2(new_n674), .A3(new_n662), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G107), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT97), .B(KEYINPUT35), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G9));
  INV_X1    g492(.A(KEYINPUT98), .ZN(new_n679));
  INV_X1    g493(.A(new_n599), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n615), .A2(new_n618), .A3(new_n604), .ZN(new_n681));
  AOI21_X1  g495(.A(KEYINPUT79), .B1(new_n624), .B2(new_n625), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n602), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n626), .A2(new_n603), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n683), .A2(new_n334), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n631), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n629), .A2(KEYINPUT25), .A3(new_n334), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n680), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n624), .A2(new_n625), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n603), .A2(KEYINPUT36), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n634), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n679), .B1(new_n688), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n633), .A2(KEYINPUT98), .A3(new_n692), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g510(.A(KEYINPUT99), .B1(new_n646), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g511(.A(G472), .B1(new_n645), .B2(new_n508), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n694), .A2(new_n695), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n593), .A2(new_n594), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT99), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n698), .A2(new_n699), .A3(new_n700), .A4(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n697), .A2(new_n524), .A3(new_n528), .A4(new_n702), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT37), .B(G110), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G12));
  NAND2_X1  g519(.A1(new_n648), .A2(new_n649), .ZN(new_n706));
  INV_X1    g520(.A(G900), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n452), .B1(new_n453), .B2(new_n707), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n706), .A2(new_n673), .A3(new_n708), .ZN(new_n709));
  AOI22_X1  g523(.A1(new_n526), .A2(new_n514), .B1(new_n694), .B2(new_n695), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n598), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(KEYINPUT100), .B(G128), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G30));
  XOR2_X1   g527(.A(new_n708), .B(KEYINPUT39), .Z(new_n714));
  AND2_X1   g528(.A1(new_n527), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT40), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n543), .A2(new_n576), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(G472), .A3(new_n587), .ZN(new_n718));
  NAND2_X1  g532(.A1(G472), .A2(G902), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g534(.A(new_n720), .B(KEYINPUT101), .Z(new_n721));
  OAI21_X1  g535(.A(new_n721), .B1(new_n595), .B2(new_n597), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n331), .B1(new_n329), .B2(new_n330), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(KEYINPUT38), .ZN(new_n726));
  AOI22_X1  g540(.A1(new_n381), .A2(new_n388), .B1(new_n445), .B2(new_n449), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n649), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n726), .A2(new_n699), .A3(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n716), .A2(new_n722), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G143), .ZN(G45));
  INV_X1    g545(.A(new_n708), .ZN(new_n732));
  INV_X1    g546(.A(new_n652), .ZN(new_n733));
  OAI21_X1  g547(.A(KEYINPUT33), .B1(new_n374), .B2(new_n377), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n384), .A2(new_n385), .A3(new_n653), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n450), .B(new_n732), .C1(new_n736), .C2(new_n657), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n706), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n598), .A2(new_n738), .A3(new_n710), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G146), .ZN(G48));
  NAND2_X1  g554(.A1(new_n511), .A2(new_n512), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n516), .B1(new_n741), .B2(new_n334), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n742), .A2(new_n513), .A3(new_n460), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n598), .A2(new_n661), .A3(new_n637), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT41), .B(G113), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G15));
  NAND4_X1  g560(.A1(new_n598), .A2(new_n637), .A3(new_n674), .A4(new_n743), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G116), .ZN(G18));
  AND2_X1   g562(.A1(new_n699), .A2(new_n456), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n333), .A2(new_n743), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n598), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G119), .ZN(G21));
  OAI211_X1 g566(.A(new_n727), .B(new_n649), .C1(new_n723), .C2(new_n724), .ZN(new_n753));
  INV_X1    g567(.A(new_n743), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n753), .A2(new_n455), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n544), .A2(new_n546), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n576), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n596), .B1(new_n590), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n593), .A2(new_n334), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n758), .B1(new_n759), .B2(G472), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n755), .A2(new_n637), .A3(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G122), .ZN(G24));
  INV_X1    g576(.A(new_n758), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n698), .A2(new_n699), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n737), .A2(KEYINPUT102), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT102), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n659), .A2(new_n766), .A3(new_n450), .A4(new_n732), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n765), .A2(new_n767), .A3(new_n333), .A4(new_n743), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(new_n393), .ZN(G27));
  OAI21_X1  g584(.A(KEYINPUT32), .B1(new_n645), .B2(new_n596), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n593), .A2(new_n581), .A3(new_n594), .ZN(new_n772));
  AOI22_X1  g586(.A1(new_n771), .A2(new_n772), .B1(G472), .B2(new_n579), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT104), .B1(new_n773), .B2(new_n636), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT104), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n598), .A2(new_n775), .A3(new_n637), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n765), .A2(new_n767), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT103), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n520), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n519), .A2(KEYINPUT103), .A3(new_n506), .A4(new_n505), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n779), .A2(new_n461), .A3(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n322), .A2(new_n649), .A3(new_n332), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n777), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n774), .A2(new_n776), .A3(new_n784), .A4(KEYINPUT42), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n598), .A2(new_n637), .A3(new_n777), .A4(new_n783), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT42), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G131), .ZN(G33));
  NOR2_X1   g604(.A1(new_n673), .A2(new_n708), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n598), .A2(new_n637), .A3(new_n791), .A4(new_n783), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G134), .ZN(G36));
  NAND2_X1  g607(.A1(new_n500), .A2(new_n504), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT45), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n516), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n796), .B1(new_n795), .B2(new_n794), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n797), .A2(new_n506), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(KEYINPUT46), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT105), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT105), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n798), .A2(new_n801), .A3(KEYINPUT46), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n519), .B1(new_n798), .B2(KEYINPUT46), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n461), .A3(new_n714), .ZN(new_n807));
  XOR2_X1   g621(.A(new_n807), .B(KEYINPUT106), .Z(new_n808));
  OAI211_X1 g622(.A(new_n449), .B(new_n445), .C1(new_n736), .C2(new_n657), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(KEYINPUT107), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT43), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n809), .A2(KEYINPUT107), .A3(KEYINPUT43), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n646), .A2(new_n812), .A3(new_n699), .A4(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT44), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n782), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n816), .B1(new_n815), .B2(new_n814), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n808), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(new_n480), .ZN(G39));
  NAND3_X1  g633(.A1(new_n806), .A2(KEYINPUT47), .A3(new_n461), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT47), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n804), .B1(new_n800), .B2(new_n802), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n821), .B1(new_n822), .B2(new_n460), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n637), .A2(new_n782), .A3(new_n737), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n824), .A2(new_n773), .A3(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(G140), .ZN(G42));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n828));
  INV_X1    g642(.A(new_n782), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n760), .A2(new_n637), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n812), .A2(new_n452), .A3(new_n813), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n742), .A2(new_n513), .A3(new_n461), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n829), .B(new_n832), .C1(new_n824), .C2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n829), .A2(new_n743), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n831), .A2(new_n764), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT50), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n726), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n743), .A2(new_n188), .ZN(new_n841));
  XOR2_X1   g655(.A(new_n841), .B(KEYINPUT115), .Z(new_n842));
  NAND3_X1  g656(.A1(new_n832), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n843), .B1(new_n837), .B2(new_n838), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n837), .A2(new_n838), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n832), .A2(new_n840), .A3(new_n845), .A4(new_n842), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n836), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n637), .A2(new_n452), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n722), .A2(new_n835), .A3(new_n848), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n849), .A2(KEYINPUT117), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(KEYINPUT117), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n659), .A2(new_n450), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n834), .A2(new_n847), .A3(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT51), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n854), .A2(KEYINPUT118), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT118), .B1(new_n854), .B2(new_n855), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n774), .A2(new_n776), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n859), .A2(new_n831), .A3(new_n835), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT48), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n860), .B(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n832), .A2(new_n750), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n863), .A2(G952), .A3(new_n291), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n850), .A2(new_n851), .ZN(new_n865));
  INV_X1    g679(.A(new_n660), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n862), .A2(KEYINPUT119), .A3(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT119), .B1(new_n862), .B2(new_n867), .ZN(new_n870));
  OAI22_X1  g684(.A1(new_n869), .A2(new_n870), .B1(new_n855), .B2(new_n854), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n828), .B1(new_n858), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n857), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n854), .A2(KEYINPUT118), .A3(new_n855), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n854), .A2(new_n855), .ZN(new_n876));
  INV_X1    g690(.A(new_n870), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n876), .B1(new_n877), .B2(new_n868), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n875), .A2(new_n878), .A3(KEYINPUT120), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n872), .A2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT114), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n638), .A2(new_n663), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT108), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(new_n389), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n885), .A2(new_n450), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n333), .A2(new_n886), .A3(new_n650), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT109), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n333), .A2(new_n886), .A3(KEYINPUT109), .A4(new_n650), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n889), .A2(new_n647), .A3(new_n662), .A4(new_n890), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n703), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n638), .A2(KEYINPUT108), .A3(new_n663), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n884), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n777), .A2(new_n760), .A3(new_n783), .A4(new_n699), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n792), .A2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT110), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n381), .A2(new_n388), .A3(new_n732), .ZN(new_n898));
  OR2_X1    g712(.A1(new_n671), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n897), .B1(new_n899), .B2(new_n782), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n671), .A2(new_n898), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n725), .A2(new_n901), .A3(KEYINPUT110), .A4(new_n649), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n903), .A2(new_n598), .A3(new_n710), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT111), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n527), .A2(new_n699), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n773), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT111), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n907), .A2(new_n908), .A3(new_n903), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n896), .B1(new_n905), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n881), .B1(new_n894), .B2(new_n911), .ZN(new_n912));
  AND4_X1   g726(.A1(new_n744), .A2(new_n747), .A3(new_n751), .A4(new_n761), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n789), .A2(KEYINPUT53), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n769), .B1(new_n907), .B2(new_n709), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT52), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n633), .A2(new_n692), .A3(new_n732), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n781), .A2(new_n753), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n722), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n915), .A2(new_n916), .A3(new_n739), .A4(new_n919), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n777), .A2(new_n760), .A3(new_n750), .A4(new_n699), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n711), .A2(new_n739), .A3(new_n919), .A4(new_n921), .ZN(new_n922));
  XOR2_X1   g736(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n920), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n914), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(KEYINPUT108), .B1(new_n638), .B2(new_n663), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n703), .A2(new_n891), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n930), .A2(new_n910), .A3(KEYINPUT114), .A4(new_n893), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n912), .A2(new_n927), .A3(new_n931), .ZN(new_n932));
  XNOR2_X1  g746(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n744), .A2(new_n747), .A3(new_n751), .A4(new_n761), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n934), .B1(new_n785), .B2(new_n788), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n935), .A2(new_n893), .A3(new_n930), .A4(new_n910), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n922), .A2(KEYINPUT52), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n920), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n933), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT54), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n932), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n936), .A2(new_n926), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n942), .A2(KEYINPUT53), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n936), .A2(new_n938), .A3(new_n933), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n941), .B1(new_n945), .B2(new_n940), .ZN(new_n946));
  OAI22_X1  g760(.A1(new_n880), .A2(new_n946), .B1(G952), .B2(G953), .ZN(new_n947));
  INV_X1    g761(.A(new_n722), .ZN(new_n948));
  NOR4_X1   g762(.A1(new_n636), .A2(new_n809), .A3(new_n188), .A4(new_n460), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n742), .A2(new_n513), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT49), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n948), .A2(new_n726), .A3(new_n949), .A4(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n947), .A2(new_n952), .ZN(G75));
  NAND2_X1  g767(.A1(new_n932), .A2(new_n939), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n508), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n955), .A2(new_n331), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n956), .A2(KEYINPUT56), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n258), .A2(new_n295), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(new_n293), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT55), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n291), .A2(G952), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  XOR2_X1   g777(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n964));
  NAND2_X1  g778(.A1(new_n960), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n963), .B1(new_n956), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n961), .A2(new_n966), .ZN(G51));
  NAND2_X1  g781(.A1(new_n954), .A2(KEYINPUT54), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n941), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n506), .B(KEYINPUT57), .Z(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n741), .ZN(new_n972));
  OR2_X1    g786(.A1(new_n955), .A2(new_n797), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n962), .B1(new_n972), .B2(new_n973), .ZN(G54));
  AND4_X1   g788(.A1(KEYINPUT58), .A2(new_n954), .A3(G475), .A4(new_n508), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n963), .B1(new_n975), .B2(new_n439), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(new_n439), .B2(new_n975), .ZN(G60));
  NAND2_X1  g791(.A1(new_n734), .A2(new_n735), .ZN(new_n978));
  NAND2_X1  g792(.A1(G478), .A2(G902), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT59), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n978), .B1(new_n946), .B2(new_n980), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n969), .A2(new_n978), .A3(new_n980), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n981), .A2(new_n982), .A3(new_n962), .ZN(G63));
  INV_X1    g797(.A(KEYINPUT61), .ZN(new_n984));
  NAND2_X1  g798(.A1(G217), .A2(G902), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT60), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n986), .B1(new_n932), .B2(new_n939), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n691), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n963), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n987), .A2(new_n629), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n984), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n986), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n954), .A2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n629), .ZN(new_n994));
  AOI21_X1  g808(.A(KEYINPUT122), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT122), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n987), .A2(new_n996), .A3(new_n629), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n988), .A2(KEYINPUT61), .A3(new_n963), .ZN(new_n999));
  INV_X1    g813(.A(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(KEYINPUT123), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n993), .A2(KEYINPUT122), .A3(new_n994), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n996), .B1(new_n987), .B2(new_n629), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT123), .ZN(new_n1005));
  NOR3_X1   g819(.A1(new_n1004), .A2(new_n999), .A3(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n991), .B1(new_n1001), .B2(new_n1006), .ZN(G66));
  INV_X1    g821(.A(new_n454), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n291), .B1(new_n1008), .B2(G224), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n894), .A2(new_n934), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1009), .B1(new_n1011), .B2(new_n291), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n958), .B1(G898), .B2(new_n291), .ZN(new_n1013));
  XOR2_X1   g827(.A(new_n1012), .B(new_n1013), .Z(G69));
  NOR2_X1   g828(.A1(new_n773), .A2(new_n636), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n660), .B1(new_n885), .B2(new_n450), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n1015), .A2(new_n715), .A3(new_n829), .A4(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n826), .A2(new_n1017), .ZN(new_n1018));
  AND2_X1   g832(.A1(new_n915), .A2(new_n739), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(new_n730), .ZN(new_n1020));
  AOI211_X1 g834(.A(new_n1018), .B(new_n818), .C1(KEYINPUT62), .C2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1020), .A2(KEYINPUT62), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1022), .B(KEYINPUT124), .Z(new_n1023));
  NAND2_X1  g837(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n571), .A2(new_n573), .ZN(new_n1025));
  XOR2_X1   g839(.A(new_n1025), .B(new_n436), .Z(new_n1026));
  AOI21_X1  g840(.A(G953), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n826), .A2(new_n792), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n818), .A2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n859), .A2(new_n753), .ZN(new_n1030));
  INV_X1    g844(.A(new_n1030), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n789), .B1(new_n808), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g846(.A(new_n1032), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1029), .A2(new_n1033), .A3(new_n1019), .ZN(new_n1034));
  INV_X1    g848(.A(KEYINPUT125), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g850(.A(new_n1026), .ZN(new_n1037));
  NAND4_X1  g851(.A1(new_n1029), .A2(new_n1033), .A3(KEYINPUT125), .A4(new_n1019), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1037), .A2(G227), .ZN(new_n1040));
  AOI211_X1 g854(.A(new_n707), .B(new_n291), .C1(new_n1026), .C2(new_n497), .ZN(new_n1041));
  AOI22_X1  g855(.A1(new_n1027), .A2(new_n1039), .B1(new_n1040), .B2(new_n1041), .ZN(G72));
  XNOR2_X1  g856(.A(new_n575), .B(KEYINPUT126), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1043), .A2(new_n576), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n1036), .A2(new_n1038), .A3(new_n1010), .ZN(new_n1045));
  XOR2_X1   g859(.A(new_n719), .B(KEYINPUT63), .Z(new_n1046));
  AOI21_X1  g860(.A(new_n1044), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AND2_X1   g861(.A1(new_n575), .A2(new_n576), .ZN(new_n1048));
  OAI21_X1  g862(.A(new_n1046), .B1(new_n1048), .B2(new_n582), .ZN(new_n1049));
  XNOR2_X1  g863(.A(new_n1049), .B(KEYINPUT127), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n963), .B1(new_n945), .B2(new_n1050), .ZN(new_n1051));
  OR2_X1    g865(.A1(new_n1043), .A2(new_n576), .ZN(new_n1052));
  NAND3_X1  g866(.A1(new_n1021), .A2(new_n1023), .A3(new_n1010), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n1052), .B1(new_n1053), .B2(new_n1046), .ZN(new_n1054));
  NOR3_X1   g868(.A1(new_n1047), .A2(new_n1051), .A3(new_n1054), .ZN(G57));
endmodule


