//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1 1 0 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G125), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT78), .B1(new_n190), .B2(KEYINPUT77), .ZN(new_n191));
  INV_X1    g005(.A(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  OAI211_X1 g007(.A(KEYINPUT78), .B(G140), .C1(new_n190), .C2(KEYINPUT77), .ZN(new_n194));
  AND2_X1   g008(.A1(G125), .A2(G140), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT78), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n193), .A2(KEYINPUT16), .A3(new_n194), .A4(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT79), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  AOI22_X1  g014(.A1(new_n191), .A2(new_n192), .B1(new_n196), .B2(new_n195), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n201), .A2(KEYINPUT79), .A3(KEYINPUT16), .A4(new_n194), .ZN(new_n202));
  NOR3_X1   g016(.A1(new_n190), .A2(KEYINPUT16), .A3(G140), .ZN(new_n203));
  XNOR2_X1  g017(.A(new_n203), .B(KEYINPUT80), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n200), .A2(new_n202), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n200), .A2(G146), .A3(new_n202), .A4(new_n204), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  XOR2_X1   g023(.A(KEYINPUT24), .B(G110), .Z(new_n210));
  OR2_X1    g024(.A1(KEYINPUT69), .A2(G119), .ZN(new_n211));
  NAND2_X1  g025(.A1(KEYINPUT69), .A2(G119), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(G128), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G128), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G119), .ZN(new_n215));
  AND3_X1   g029(.A1(new_n210), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  AND2_X1   g030(.A1(KEYINPUT69), .A2(G119), .ZN(new_n217));
  NOR2_X1   g031(.A1(KEYINPUT69), .A2(G119), .ZN(new_n218));
  NOR3_X1   g032(.A1(new_n217), .A2(new_n218), .A3(new_n214), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT23), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT75), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT75), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n213), .A2(new_n222), .A3(KEYINPUT23), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n214), .B1(new_n217), .B2(new_n218), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT76), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI211_X1 g040(.A(KEYINPUT76), .B(new_n214), .C1(new_n217), .C2(new_n218), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n221), .A2(new_n223), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n214), .A2(KEYINPUT23), .A3(G119), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n216), .B1(new_n230), .B2(G110), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n209), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(G125), .A2(G140), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n195), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n234), .A2(G146), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n208), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G110), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n228), .A2(new_n238), .A3(new_n229), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n210), .B1(new_n215), .B2(new_n213), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT81), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n240), .B(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n237), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT22), .B(G137), .ZN(new_n245));
  INV_X1    g059(.A(G221), .ZN(new_n246));
  INV_X1    g060(.A(G234), .ZN(new_n247));
  NOR3_X1   g061(.A1(new_n246), .A2(new_n247), .A3(G953), .ZN(new_n248));
  XOR2_X1   g062(.A(new_n245), .B(new_n248), .Z(new_n249));
  AND3_X1   g063(.A1(new_n232), .A2(new_n244), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n249), .B1(new_n232), .B2(new_n244), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT25), .B1(new_n252), .B2(new_n188), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n232), .A2(new_n244), .ZN(new_n254));
  INV_X1    g068(.A(new_n249), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n232), .A2(new_n244), .A3(new_n249), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n256), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n189), .B1(new_n253), .B2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n189), .A2(G902), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n252), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(G472), .A2(G902), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT32), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT65), .ZN(new_n266));
  INV_X1    g080(.A(G143), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n266), .B1(new_n267), .B2(G146), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n206), .A2(KEYINPUT65), .A3(G143), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n267), .A2(G146), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  AND2_X1   g085(.A1(KEYINPUT0), .A2(G128), .ZN(new_n272));
  OR3_X1    g086(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n206), .A2(G143), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n272), .B1(new_n276), .B2(new_n270), .ZN(new_n277));
  AOI22_X1  g091(.A1(new_n271), .A2(new_n272), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G131), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT67), .ZN(new_n280));
  INV_X1    g094(.A(G137), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n280), .B1(new_n281), .B2(G134), .ZN(new_n282));
  INV_X1    g096(.A(G134), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(KEYINPUT67), .A3(G137), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n281), .A2(KEYINPUT66), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT66), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G137), .ZN(new_n288));
  AND2_X1   g102(.A1(KEYINPUT11), .A2(G134), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n286), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n281), .A2(G134), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT11), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AND4_X1   g107(.A1(new_n279), .A2(new_n285), .A3(new_n290), .A4(new_n293), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n282), .A2(new_n284), .B1(new_n291), .B2(new_n292), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n279), .B1(new_n295), .B2(new_n290), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n278), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n211), .A2(G116), .A3(new_n212), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT70), .ZN(new_n299));
  INV_X1    g113(.A(G116), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(KEYINPUT70), .A2(G116), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(G119), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G113), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT2), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT2), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G113), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n298), .A2(new_n303), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n308), .B1(new_n298), .B2(new_n303), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT66), .B(G137), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n291), .B1(new_n312), .B2(G134), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G131), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n276), .A2(new_n270), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT1), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n316), .B1(G143), .B2(new_n206), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n315), .B1(new_n317), .B2(new_n214), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n214), .A2(KEYINPUT1), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n268), .A2(new_n269), .A3(new_n319), .A4(new_n270), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n295), .A2(new_n279), .A3(new_n290), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n314), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n297), .A2(new_n311), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT71), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n297), .A2(new_n311), .A3(KEYINPUT71), .A4(new_n323), .ZN(new_n327));
  NOR2_X1   g141(.A1(G237), .A2(G953), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G210), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n329), .B(KEYINPUT27), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT26), .B(G101), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n330), .B(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n326), .A2(new_n327), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT72), .ZN(new_n334));
  OR2_X1    g148(.A1(new_n309), .A2(new_n310), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n285), .A2(new_n290), .A3(new_n293), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G131), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n322), .ZN(new_n338));
  AOI22_X1  g152(.A1(G131), .A2(new_n313), .B1(new_n318), .B2(new_n320), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n338), .A2(new_n278), .B1(new_n339), .B2(new_n322), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT30), .ZN(new_n341));
  INV_X1    g155(.A(new_n323), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT68), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n297), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n338), .A2(KEYINPUT68), .A3(new_n278), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n342), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n335), .B(new_n341), .C1(new_n346), .C2(KEYINPUT30), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT72), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n326), .A2(new_n348), .A3(new_n327), .A4(new_n332), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n334), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT31), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n334), .A2(new_n347), .A3(KEYINPUT31), .A4(new_n349), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  XOR2_X1   g168(.A(new_n332), .B(KEYINPUT73), .Z(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n344), .A2(new_n345), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n311), .B1(new_n357), .B2(new_n323), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n326), .A2(new_n327), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT28), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT28), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n324), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n356), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n265), .B1(new_n354), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G472), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n360), .A2(new_n362), .A3(new_n356), .ZN(new_n367));
  INV_X1    g181(.A(new_n359), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n347), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n332), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n367), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n326), .A2(KEYINPUT74), .A3(new_n327), .ZN(new_n374));
  OR2_X1    g188(.A1(new_n340), .A2(new_n311), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(KEYINPUT74), .B1(new_n326), .B2(new_n327), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT28), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n362), .A2(KEYINPUT29), .A3(new_n332), .ZN(new_n379));
  AOI21_X1  g193(.A(G902), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n366), .B1(new_n373), .B2(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n365), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT32), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n363), .B1(new_n352), .B2(new_n353), .ZN(new_n384));
  INV_X1    g198(.A(new_n264), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n263), .B1(new_n382), .B2(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(KEYINPUT9), .B(G234), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n246), .B1(new_n389), .B2(new_n188), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n267), .A2(G146), .ZN(new_n393));
  OAI21_X1  g207(.A(G128), .B1(new_n393), .B2(new_n316), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n320), .ZN(new_n396));
  INV_X1    g210(.A(G104), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT3), .B1(new_n397), .B2(G107), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT3), .ZN(new_n399));
  INV_X1    g213(.A(G107), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n400), .A3(G104), .ZN(new_n401));
  INV_X1    g215(.A(G101), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n397), .A2(G107), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n398), .A2(new_n401), .A3(new_n402), .A4(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n397), .A2(G107), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n400), .A2(G104), .ZN(new_n406));
  OAI21_X1  g220(.A(G101), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n396), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT10), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n410), .B1(new_n318), .B2(new_n320), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n409), .A2(new_n410), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n398), .A2(new_n401), .A3(new_n403), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(KEYINPUT82), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT82), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n398), .A2(new_n401), .A3(new_n415), .A4(new_n403), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(G101), .A3(new_n416), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n404), .A2(KEYINPUT4), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n402), .A2(KEYINPUT4), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n414), .A2(new_n416), .A3(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n419), .A2(new_n278), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n338), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n412), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n318), .A2(new_n320), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n404), .A2(new_n407), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n409), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n428), .A2(KEYINPUT12), .A3(new_n338), .ZN(new_n429));
  AOI21_X1  g243(.A(KEYINPUT12), .B1(new_n428), .B2(new_n338), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n424), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(G110), .B(G140), .ZN(new_n432));
  INV_X1    g246(.A(G953), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n433), .A2(G227), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n432), .B(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT83), .ZN(new_n437));
  INV_X1    g251(.A(new_n435), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n424), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n421), .A2(new_n278), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n440), .B1(new_n417), .B2(new_n418), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n411), .A2(new_n408), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n426), .B1(new_n320), .B2(new_n395), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n442), .B1(new_n443), .B2(KEYINPUT10), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n338), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n439), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n437), .B1(new_n424), .B2(new_n438), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n436), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT84), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT84), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n436), .B(new_n450), .C1(new_n446), .C2(new_n447), .ZN(new_n451));
  AOI21_X1  g265(.A(G902), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G469), .ZN(new_n453));
  OAI21_X1  g267(.A(KEYINPUT85), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n451), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n424), .A2(new_n438), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT83), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(new_n445), .A3(new_n439), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n450), .B1(new_n458), .B2(new_n436), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n188), .B1(new_n455), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT85), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n461), .A3(G469), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n412), .A2(new_n422), .A3(new_n423), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n423), .B1(new_n412), .B2(new_n422), .ZN(new_n464));
  OAI211_X1 g278(.A(KEYINPUT86), .B(new_n435), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n424), .B(new_n438), .C1(new_n429), .C2(new_n430), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n445), .A2(new_n424), .ZN(new_n468));
  AOI21_X1  g282(.A(KEYINPUT86), .B1(new_n468), .B2(new_n435), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n453), .B(new_n188), .C1(new_n467), .C2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT87), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n435), .B1(new_n463), .B2(new_n464), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT86), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(new_n466), .A3(new_n465), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n476), .A2(KEYINPUT87), .A3(new_n453), .A4(new_n188), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n454), .A2(new_n462), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(G214), .B1(G237), .B2(G902), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n328), .A2(G143), .A3(G214), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(G143), .B1(new_n328), .B2(G214), .ZN(new_n483));
  OAI21_X1  g297(.A(G131), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT17), .ZN(new_n485));
  INV_X1    g299(.A(G237), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(new_n433), .A3(G214), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n267), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(new_n279), .A3(new_n481), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n484), .A2(new_n485), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n481), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(KEYINPUT17), .A3(G131), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n207), .A2(new_n208), .A3(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(G113), .B(G122), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(G104), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT94), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n491), .A2(KEYINPUT18), .A3(G131), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT18), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n488), .B(new_n481), .C1(new_n500), .C2(new_n279), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n201), .A2(new_n194), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n235), .B1(new_n503), .B2(G146), .ZN(new_n504));
  OR2_X1    g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n494), .A2(new_n498), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n188), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n498), .B1(new_n494), .B2(new_n505), .ZN(new_n508));
  OAI21_X1  g322(.A(G475), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT20), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n496), .B1(new_n502), .B2(new_n504), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n201), .A2(KEYINPUT19), .A3(new_n194), .ZN(new_n512));
  INV_X1    g326(.A(new_n234), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n512), .B1(KEYINPUT19), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g328(.A1(new_n514), .A2(new_n206), .B1(new_n484), .B2(new_n489), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n511), .B1(new_n515), .B2(new_n208), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n494), .A2(new_n505), .ZN(new_n517));
  INV_X1    g331(.A(new_n496), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(G475), .A2(G902), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n510), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n496), .B1(new_n494), .B2(new_n505), .ZN(new_n522));
  INV_X1    g336(.A(new_n520), .ZN(new_n523));
  NOR4_X1   g337(.A1(new_n522), .A2(KEYINPUT20), .A3(new_n516), .A4(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n509), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n301), .A2(G122), .A3(new_n302), .ZN(new_n526));
  OR2_X1    g340(.A1(new_n300), .A2(G122), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n526), .A2(new_n400), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n267), .A2(G128), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n214), .A2(G143), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n529), .A2(new_n530), .A3(G134), .ZN(new_n531));
  AOI21_X1  g345(.A(G134), .B1(new_n529), .B2(new_n530), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT14), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n526), .A2(new_n534), .A3(new_n527), .ZN(new_n535));
  OAI21_X1  g349(.A(G107), .B1(new_n526), .B2(new_n534), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n528), .B(new_n533), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n529), .A2(new_n530), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT13), .B1(new_n214), .B2(G143), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n538), .B1(new_n283), .B2(new_n539), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT13), .A4(G134), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n528), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n400), .B1(new_n526), .B2(new_n527), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n388), .A2(new_n187), .A3(G953), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n537), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n546), .B1(new_n537), .B2(new_n545), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n188), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT95), .ZN(new_n551));
  INV_X1    g365(.A(G478), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(KEYINPUT15), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT95), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n554), .B(new_n188), .C1(new_n548), .C2(new_n549), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n551), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  OAI211_X1 g370(.A(G902), .B(G953), .C1(new_n247), .C2(new_n486), .ZN(new_n557));
  XOR2_X1   g371(.A(new_n557), .B(KEYINPUT96), .Z(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT21), .B(G898), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n433), .A2(G952), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n562), .B1(new_n247), .B2(new_n486), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  OR2_X1    g378(.A1(new_n550), .A2(new_n553), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n556), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n525), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT6), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT88), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n298), .A2(new_n303), .A3(KEYINPUT5), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT5), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n211), .A2(new_n571), .A3(G116), .A4(new_n212), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G113), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n569), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n309), .A2(new_n426), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n298), .A2(new_n303), .A3(KEYINPUT5), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n576), .A2(KEYINPUT88), .A3(G113), .A4(new_n572), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n574), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT89), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n574), .A2(new_n575), .A3(KEYINPUT89), .A4(new_n577), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n335), .A2(new_n421), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n580), .A2(new_n581), .B1(new_n582), .B2(new_n419), .ZN(new_n583));
  XNOR2_X1  g397(.A(G110), .B(G122), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n568), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n580), .A2(new_n581), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n582), .A2(new_n419), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n584), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  OR3_X1    g405(.A1(new_n278), .A2(KEYINPUT90), .A3(new_n190), .ZN(new_n592));
  OAI21_X1  g406(.A(KEYINPUT90), .B1(new_n278), .B2(new_n190), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n425), .A2(KEYINPUT91), .A3(new_n190), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT91), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n596), .B1(new_n321), .B2(G125), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n433), .A2(G224), .ZN(new_n600));
  XOR2_X1   g414(.A(new_n600), .B(KEYINPUT92), .Z(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n594), .A2(new_n598), .A3(new_n601), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n588), .A2(new_n568), .A3(new_n589), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n591), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(G210), .B1(G237), .B2(G902), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(KEYINPUT93), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n600), .A2(KEYINPUT7), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n598), .A2(new_n592), .A3(new_n593), .A4(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n278), .A2(new_n190), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n613), .B1(new_n595), .B2(new_n597), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n612), .B1(new_n611), .B2(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(new_n584), .B(KEYINPUT8), .Z(new_n616));
  NAND2_X1  g430(.A1(new_n574), .A2(new_n577), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n426), .B1(new_n617), .B2(new_n309), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n575), .B1(new_n570), .B2(new_n573), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n616), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n583), .A2(new_n584), .ZN(new_n622));
  AOI21_X1  g436(.A(G902), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n607), .A2(new_n610), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n610), .B1(new_n607), .B2(new_n623), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n480), .B(new_n567), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n387), .A2(new_n391), .A3(new_n479), .A4(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G101), .ZN(G3));
  AND2_X1   g443(.A1(new_n479), .A2(new_n391), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n354), .A2(new_n364), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n264), .ZN(new_n632));
  OAI21_X1  g446(.A(G472), .B1(new_n384), .B2(G902), .ZN(new_n633));
  INV_X1    g447(.A(new_n262), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n256), .A2(new_n188), .A3(new_n257), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT25), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n258), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n634), .B1(new_n638), .B2(new_n189), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n632), .A2(new_n633), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT97), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n547), .A2(new_n641), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n642), .B(KEYINPUT33), .C1(new_n548), .C2(new_n549), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n537), .A2(new_n545), .ZN(new_n644));
  INV_X1    g458(.A(new_n546), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT33), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n646), .B(new_n547), .C1(new_n641), .C2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n643), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n552), .A2(G902), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(KEYINPUT98), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n551), .A2(new_n552), .A3(new_n555), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT98), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n649), .A2(new_n654), .A3(new_n650), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n652), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  AND3_X1   g470(.A1(new_n656), .A2(new_n525), .A3(new_n564), .ZN(new_n657));
  INV_X1    g471(.A(new_n480), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n607), .A2(new_n623), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n658), .B1(new_n659), .B2(new_n608), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n607), .A2(new_n609), .A3(new_n623), .ZN(new_n661));
  AND3_X1   g475(.A1(new_n657), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n630), .A2(new_n640), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT34), .B(G104), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G6));
  NAND2_X1  g479(.A1(new_n556), .A2(new_n565), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n666), .B(new_n509), .C1(new_n521), .C2(new_n524), .ZN(new_n667));
  XOR2_X1   g481(.A(new_n564), .B(KEYINPUT99), .Z(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n660), .A2(new_n661), .A3(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n630), .A2(new_n640), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(new_n672), .B(KEYINPUT100), .Z(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT35), .B(G107), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G9));
  NOR2_X1   g489(.A1(new_n255), .A2(KEYINPUT36), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n254), .B(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n261), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n260), .A2(new_n678), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n679), .A2(new_n632), .A3(new_n633), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n680), .A2(new_n479), .A3(new_n391), .A4(new_n627), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT37), .B(G110), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G12));
  NAND2_X1  g497(.A1(new_n519), .A2(new_n520), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT20), .ZN(new_n685));
  INV_X1    g499(.A(new_n524), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n507), .A2(new_n508), .ZN(new_n687));
  AOI22_X1  g501(.A1(new_n685), .A2(new_n686), .B1(new_n687), .B2(G475), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT102), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n558), .A2(G900), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT101), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n563), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n690), .A2(KEYINPUT101), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n688), .A2(new_n689), .A3(new_n666), .A4(new_n695), .ZN(new_n696));
  OAI21_X1  g510(.A(KEYINPUT102), .B1(new_n667), .B2(new_n694), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n479), .A2(new_n698), .A3(new_n391), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n384), .A2(new_n265), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n373), .A2(new_n380), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(G472), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n700), .A2(new_n386), .A3(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n661), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n609), .B1(new_n607), .B2(new_n623), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n704), .A2(new_n705), .A3(new_n658), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n703), .A2(new_n706), .A3(new_n679), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n699), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(new_n214), .ZN(G30));
  XOR2_X1   g523(.A(new_n694), .B(KEYINPUT39), .Z(new_n710));
  NAND2_X1  g524(.A1(new_n630), .A2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT104), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT40), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n711), .B(KEYINPUT104), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(KEYINPUT40), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n624), .A2(new_n625), .ZN(new_n718));
  XOR2_X1   g532(.A(new_n718), .B(KEYINPUT38), .Z(new_n719));
  OAI21_X1  g533(.A(new_n355), .B1(new_n376), .B2(new_n377), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n720), .A2(new_n350), .ZN(new_n721));
  OAI21_X1  g535(.A(G472), .B1(new_n721), .B2(G902), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n700), .A2(new_n386), .A3(new_n722), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n525), .A2(new_n666), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n189), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n727), .B1(new_n637), .B2(new_n258), .ZN(new_n728));
  INV_X1    g542(.A(new_n678), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n719), .A2(new_n726), .A3(new_n480), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(KEYINPUT103), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n715), .A2(new_n717), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G143), .ZN(G45));
  NAND2_X1  g548(.A1(new_n656), .A2(new_n525), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n694), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n479), .A2(new_n391), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n707), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n206), .ZN(G48));
  AOI21_X1  g553(.A(new_n453), .B1(new_n476), .B2(new_n188), .ZN(new_n740));
  AOI211_X1 g554(.A(new_n390), .B(new_n740), .C1(new_n472), .C2(new_n477), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n662), .A2(new_n703), .A3(new_n639), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(KEYINPUT41), .B(G113), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G15));
  NAND4_X1  g558(.A1(new_n671), .A2(new_n703), .A3(new_n741), .A4(new_n639), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT105), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n387), .A2(KEYINPUT105), .A3(new_n671), .A4(new_n741), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G116), .ZN(G18));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n751));
  INV_X1    g565(.A(new_n567), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n730), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n703), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n740), .B1(new_n472), .B2(new_n477), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n755), .A2(new_n391), .A3(new_n661), .A4(new_n660), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n751), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n756), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n758), .A2(KEYINPUT106), .A3(new_n703), .A4(new_n753), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G119), .ZN(G21));
  XNOR2_X1  g575(.A(new_n264), .B(KEYINPUT107), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n352), .A2(new_n353), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n356), .B1(new_n378), .B2(new_n362), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n765), .A2(new_n633), .A3(new_n639), .ZN(new_n766));
  INV_X1    g580(.A(new_n740), .ZN(new_n767));
  AND4_X1   g581(.A1(new_n391), .A2(new_n478), .A3(new_n668), .A4(new_n767), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n660), .A2(new_n724), .A3(new_n661), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n766), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G122), .ZN(G24));
  NAND4_X1  g585(.A1(new_n736), .A2(new_n679), .A3(new_n765), .A4(new_n633), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n756), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(new_n190), .ZN(G27));
  INV_X1    g588(.A(KEYINPUT109), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT32), .B1(new_n631), .B2(new_n264), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n775), .B1(new_n776), .B2(new_n365), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n700), .A2(KEYINPUT109), .A3(new_n386), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n702), .A3(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n610), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n659), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n607), .A2(new_n610), .A3(new_n623), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n781), .A2(new_n480), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n453), .B1(new_n448), .B2(new_n188), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n784), .B1(new_n472), .B2(new_n477), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n656), .A2(new_n525), .A3(KEYINPUT42), .A4(new_n695), .ZN(new_n786));
  NOR4_X1   g600(.A1(new_n783), .A2(new_n785), .A3(new_n390), .A4(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n779), .A2(new_n639), .A3(new_n787), .ZN(new_n788));
  XOR2_X1   g602(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n789));
  INV_X1    g603(.A(new_n784), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n390), .B1(new_n478), .B2(new_n790), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n624), .A2(new_n625), .A3(new_n658), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n703), .A2(new_n639), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n736), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n789), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n788), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G131), .ZN(G33));
  NOR3_X1   g611(.A1(new_n783), .A2(new_n785), .A3(new_n390), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n696), .A2(new_n697), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT110), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n696), .A2(new_n697), .A3(KEYINPUT110), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n387), .A2(new_n798), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  XOR2_X1   g617(.A(KEYINPUT111), .B(G134), .Z(new_n804));
  XNOR2_X1  g618(.A(new_n803), .B(new_n804), .ZN(G36));
  INV_X1    g619(.A(KEYINPUT45), .ZN(new_n806));
  OAI21_X1  g620(.A(G469), .B1(new_n448), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n449), .A2(new_n451), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n807), .B1(new_n808), .B2(new_n806), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n453), .A2(new_n188), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT46), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n478), .B1(new_n811), .B2(KEYINPUT46), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n390), .ZN(new_n816));
  INV_X1    g630(.A(new_n656), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(new_n525), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT43), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n819), .B1(new_n525), .B2(KEYINPUT112), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n818), .B(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n730), .B1(new_n632), .B2(new_n633), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT44), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n823), .A2(new_n783), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n821), .A2(KEYINPUT44), .A3(new_n822), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n816), .A2(new_n824), .A3(new_n710), .A4(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(KEYINPUT113), .B(G137), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n826), .B(new_n827), .ZN(G39));
  NAND2_X1  g642(.A1(KEYINPUT114), .A2(KEYINPUT47), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n816), .A2(new_n829), .ZN(new_n830));
  NOR4_X1   g644(.A1(new_n703), .A2(new_n794), .A3(new_n783), .A4(new_n639), .ZN(new_n831));
  XOR2_X1   g645(.A(KEYINPUT114), .B(KEYINPUT47), .Z(new_n832));
  OAI211_X1 g646(.A(new_n830), .B(new_n831), .C1(new_n816), .C2(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(G140), .ZN(G42));
  AND2_X1   g648(.A1(new_n779), .A2(new_n639), .ZN(new_n835));
  INV_X1    g649(.A(new_n563), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n755), .A2(new_n391), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n837), .A2(new_n783), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n821), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n835), .A2(new_n839), .ZN(new_n840));
  XOR2_X1   g654(.A(new_n840), .B(KEYINPUT48), .Z(new_n841));
  AND3_X1   g655(.A1(new_n821), .A2(new_n836), .A3(new_n766), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n758), .ZN(new_n843));
  INV_X1    g657(.A(new_n723), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n639), .A2(new_n838), .A3(new_n844), .A4(new_n836), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n843), .B(new_n562), .C1(new_n735), .C2(new_n846), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n847), .A2(KEYINPUT121), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(KEYINPUT121), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n841), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n839), .A2(new_n633), .A3(new_n679), .A4(new_n765), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n845), .A2(new_n688), .A3(new_n817), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n719), .A2(new_n480), .A3(new_n837), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(new_n842), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT50), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT50), .B1(new_n853), .B2(new_n842), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n851), .B(new_n852), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n816), .A2(new_n832), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(new_n816), .B2(new_n829), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n755), .A2(new_n390), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n792), .B(new_n842), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT51), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT120), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n858), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n858), .A2(new_n864), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n865), .A2(new_n862), .A3(new_n866), .ZN(new_n867));
  OAI221_X1 g681(.A(new_n850), .B1(new_n858), .B2(new_n863), .C1(new_n867), .C2(KEYINPUT51), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n770), .A2(new_n742), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n796), .A2(new_n749), .A3(new_n760), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT119), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n688), .A2(new_n565), .A3(new_n556), .A4(new_n695), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n783), .A2(new_n873), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n874), .A2(new_n703), .A3(new_n679), .ZN(new_n875));
  AND4_X1   g689(.A1(new_n633), .A2(new_n736), .A3(new_n679), .A4(new_n765), .ZN(new_n876));
  AOI22_X1  g690(.A1(new_n875), .A2(new_n630), .B1(new_n876), .B2(new_n798), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n630), .B(new_n627), .C1(new_n387), .C2(new_n680), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n480), .B(new_n668), .C1(new_n624), .C2(new_n625), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n735), .A2(new_n667), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n881), .A2(new_n640), .A3(new_n479), .A4(new_n391), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n877), .A2(new_n878), .A3(new_n803), .A4(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n479), .A2(new_n391), .A3(new_n736), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n703), .A2(new_n706), .A3(new_n679), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n728), .A2(new_n729), .A3(new_n694), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n791), .A2(new_n706), .A3(new_n888), .ZN(new_n889));
  AOI22_X1  g703(.A1(new_n886), .A2(new_n887), .B1(new_n726), .B2(new_n889), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n479), .A2(new_n391), .A3(new_n698), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n773), .B1(new_n891), .B2(new_n887), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n890), .A2(new_n892), .A3(KEYINPUT52), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT52), .ZN(new_n894));
  OAI22_X1  g708(.A1(new_n699), .A2(new_n707), .B1(new_n756), .B2(new_n772), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n791), .A2(new_n706), .A3(new_n888), .ZN(new_n896));
  OAI22_X1  g710(.A1(new_n737), .A2(new_n707), .B1(new_n725), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n894), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n770), .A2(new_n742), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n900), .B1(new_n757), .B2(new_n759), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT119), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n901), .A2(new_n902), .A3(new_n749), .A4(new_n796), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n872), .A2(new_n885), .A3(new_n899), .A4(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT118), .ZN(new_n905));
  XOR2_X1   g719(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n871), .A2(new_n883), .ZN(new_n908));
  AOI211_X1 g722(.A(new_n905), .B(new_n907), .C1(new_n908), .C2(new_n899), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n749), .A2(new_n760), .A3(new_n870), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n788), .A2(new_n795), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n730), .B1(new_n382), .B2(new_n386), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n913), .A2(new_n391), .A3(new_n479), .A4(new_n874), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n876), .A2(new_n798), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n803), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n628), .A2(new_n882), .A3(new_n681), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n912), .A2(new_n899), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT118), .B1(new_n919), .B2(new_n906), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n869), .B(new_n904), .C1(new_n909), .C2(new_n920), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n893), .A2(new_n898), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n918), .A2(new_n749), .A3(new_n796), .A4(new_n901), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n884), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n912), .A2(new_n899), .A3(new_n918), .A4(new_n907), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT117), .B1(new_n926), .B2(KEYINPUT54), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT117), .ZN(new_n928));
  AOI211_X1 g742(.A(new_n928), .B(new_n869), .C1(new_n924), .C2(new_n925), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n921), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  OAI22_X1  g744(.A1(new_n868), .A2(new_n930), .B1(G952), .B2(G953), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n719), .A2(new_n525), .A3(new_n817), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n755), .B(KEYINPUT49), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n639), .A2(new_n391), .A3(new_n480), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT115), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n932), .A2(new_n844), .A3(new_n933), .A4(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n931), .A2(new_n936), .ZN(G75));
  AND4_X1   g751(.A1(new_n899), .A2(new_n872), .A3(new_n885), .A4(new_n903), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n906), .B1(new_n922), .B2(new_n923), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n905), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n919), .A2(KEYINPUT118), .A3(new_n906), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n938), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(KEYINPUT122), .B1(new_n942), .B2(new_n188), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n904), .B1(new_n909), .B2(new_n920), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT122), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n944), .A2(new_n945), .A3(G902), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n943), .A2(new_n609), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n591), .A2(new_n606), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(new_n605), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT55), .Z(new_n950));
  NOR2_X1   g764(.A1(new_n950), .A2(KEYINPUT56), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n433), .A2(G952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n944), .A2(G210), .A3(G902), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT56), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n953), .B1(new_n956), .B2(new_n950), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n952), .A2(new_n957), .ZN(G51));
  NOR2_X1   g772(.A1(new_n942), .A2(new_n869), .ZN(new_n959));
  INV_X1    g773(.A(new_n921), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n810), .B(KEYINPUT57), .Z(new_n962));
  OAI21_X1  g776(.A(new_n476), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n943), .A2(new_n809), .A3(new_n946), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n953), .B1(new_n963), .B2(new_n964), .ZN(G54));
  AND2_X1   g779(.A1(KEYINPUT58), .A2(G475), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n943), .A2(new_n946), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(new_n522), .B2(new_n516), .ZN(new_n968));
  INV_X1    g782(.A(new_n953), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n943), .A2(new_n946), .A3(new_n519), .A4(new_n966), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(G60));
  NAND2_X1  g785(.A1(G478), .A2(G902), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT59), .Z(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n930), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n649), .ZN(new_n976));
  AOI21_X1  g790(.A(KEYINPUT123), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT123), .ZN(new_n978));
  AOI211_X1 g792(.A(new_n978), .B(new_n649), .C1(new_n930), .C2(new_n974), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n976), .A2(new_n973), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n959), .B2(new_n960), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n969), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n977), .A2(new_n979), .A3(new_n982), .ZN(G63));
  NAND2_X1  g797(.A1(G217), .A2(G902), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT60), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n942), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(new_n677), .ZN(new_n987));
  OAI22_X1  g801(.A1(new_n942), .A2(new_n985), .B1(new_n250), .B2(new_n251), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n987), .A2(new_n969), .A3(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT61), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n987), .A2(KEYINPUT61), .A3(new_n969), .A4(new_n988), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(G66));
  INV_X1    g807(.A(G224), .ZN(new_n994));
  OAI21_X1  g808(.A(G953), .B1(new_n560), .B2(new_n994), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n910), .A2(new_n917), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n995), .B1(new_n996), .B2(G953), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n948), .B1(G898), .B2(new_n433), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n997), .B(new_n998), .ZN(G69));
  AOI21_X1  g813(.A(new_n433), .B1(G227), .B2(G900), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT126), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n895), .A2(new_n738), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n733), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g819(.A(KEYINPUT124), .B1(new_n1005), .B2(KEYINPUT62), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1005), .A2(KEYINPUT62), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT124), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT62), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n733), .A2(new_n1008), .A3(new_n1009), .A4(new_n1004), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n833), .A2(new_n826), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n880), .A2(new_n783), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n387), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1011), .B1(new_n713), .B2(new_n1013), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1006), .A2(new_n1007), .A3(new_n1010), .A4(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(new_n433), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n341), .B1(new_n346), .B2(KEYINPUT30), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1017), .B(new_n514), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n796), .A2(new_n803), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT125), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1020), .B(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n816), .A2(new_n710), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n835), .A2(new_n769), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1004), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NOR3_X1   g839(.A1(new_n1022), .A2(new_n1011), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1026), .A2(new_n433), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1018), .B1(G900), .B2(G953), .ZN(new_n1028));
  AOI22_X1  g842(.A1(new_n1027), .A2(new_n1028), .B1(new_n1001), .B2(new_n1000), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1003), .B1(new_n1019), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g844(.A(new_n1018), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1031), .B1(new_n1015), .B2(new_n433), .ZN(new_n1032));
  INV_X1    g846(.A(new_n1029), .ZN(new_n1033));
  NOR3_X1   g847(.A1(new_n1032), .A2(new_n1033), .A3(new_n1002), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n1030), .A2(new_n1034), .ZN(G72));
  NAND2_X1  g849(.A1(G472), .A2(G902), .ZN(new_n1036));
  XOR2_X1   g850(.A(new_n1036), .B(KEYINPUT63), .Z(new_n1037));
  INV_X1    g851(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1038), .B1(new_n1026), .B2(new_n996), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n347), .A2(new_n368), .A3(new_n370), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n969), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g855(.A(KEYINPUT127), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g857(.A(KEYINPUT127), .B(new_n969), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g859(.A(new_n996), .ZN(new_n1046));
  OAI21_X1  g860(.A(new_n1037), .B1(new_n1015), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n1047), .A2(new_n332), .A3(new_n369), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n1038), .B1(new_n371), .B2(new_n350), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n926), .A2(new_n1049), .ZN(new_n1050));
  AND3_X1   g864(.A1(new_n1045), .A2(new_n1048), .A3(new_n1050), .ZN(G57));
endmodule


