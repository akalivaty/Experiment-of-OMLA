//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 1 0 0 0 1 1 0 1 1 1 0 1 0 0 0 1 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1272,
    new_n1273, new_n1274, new_n1276, new_n1277, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n217), .B1(new_n202), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n222));
  INV_X1    g0022(.A(G58), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  INV_X1    g0024(.A(G68), .ZN(new_n225));
  INV_X1    g0025(.A(G238), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n208), .B1(new_n221), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(new_n224), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XOR2_X1   g0039(.A(G50), .B(G58), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  NAND3_X1  g0045(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(new_n214), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT65), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  OAI21_X1  g0049(.A(new_n248), .B1(new_n249), .B2(G20), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n206), .A2(KEYINPUT65), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT8), .B(G58), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G150), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  OAI22_X1  g0057(.A1(new_n255), .A2(new_n257), .B1(new_n201), .B2(new_n206), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n247), .B1(new_n254), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(new_n247), .ZN(new_n262));
  INV_X1    g0062(.A(G50), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n263), .B1(new_n205), .B2(G20), .ZN(new_n264));
  AOI22_X1  g0064(.A1(new_n262), .A2(new_n264), .B1(new_n263), .B2(new_n261), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n259), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n266), .B(KEYINPUT9), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G1), .A3(G13), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT3), .B(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(G222), .A2(G1698), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G223), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n270), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n274), .B1(G77), .B2(new_n270), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n269), .B1(new_n275), .B2(KEYINPUT64), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n276), .B1(KEYINPUT64), .B2(new_n275), .ZN(new_n277));
  INV_X1    g0077(.A(G41), .ZN(new_n278));
  INV_X1    g0078(.A(G45), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(G1), .A2(G13), .ZN(new_n281));
  AOI22_X1  g0081(.A1(new_n205), .A2(new_n280), .B1(new_n281), .B2(new_n268), .ZN(new_n282));
  INV_X1    g0082(.A(G274), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n283), .B1(new_n281), .B2(new_n268), .ZN(new_n284));
  AOI21_X1  g0084(.A(G1), .B1(new_n278), .B2(new_n279), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n282), .A2(G226), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n277), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G200), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n267), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AND3_X1   g0089(.A1(new_n277), .A2(G190), .A3(new_n286), .ZN(new_n290));
  OR3_X1    g0090(.A1(new_n289), .A2(new_n290), .A3(KEYINPUT10), .ZN(new_n291));
  OAI21_X1  g0091(.A(KEYINPUT10), .B1(new_n289), .B2(new_n290), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT66), .B(G179), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n287), .A2(new_n294), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n295), .B(new_n266), .C1(G169), .C2(new_n287), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n219), .A2(KEYINPUT15), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n219), .A2(KEYINPUT15), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n250), .B(new_n251), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  OAI22_X1  g0100(.A1(new_n253), .A2(new_n257), .B1(new_n206), .B2(new_n202), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n247), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT67), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n223), .A2(KEYINPUT8), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT8), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G58), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n308), .A2(new_n256), .B1(G20), .B2(G77), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n299), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n310), .A2(KEYINPUT67), .A3(new_n247), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n304), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n272), .A2(G232), .ZN(new_n313));
  NAND2_X1  g0113(.A1(G238), .A2(G1698), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n270), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT3), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G33), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G107), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AND2_X1   g0121(.A1(G33), .A2(G41), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(new_n214), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n315), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n282), .A2(G244), .B1(new_n284), .B2(new_n285), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G200), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n202), .B1(new_n205), .B2(G20), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n262), .A2(new_n328), .B1(new_n202), .B2(new_n261), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n324), .A2(new_n325), .A3(G190), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n312), .A2(new_n327), .A3(new_n329), .A4(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT67), .B1(new_n310), .B2(new_n247), .ZN(new_n332));
  INV_X1    g0132(.A(new_n247), .ZN(new_n333));
  AOI211_X1 g0133(.A(new_n303), .B(new_n333), .C1(new_n309), .C2(new_n299), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n329), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n324), .A2(new_n325), .A3(new_n294), .ZN(new_n336));
  AOI21_X1  g0136(.A(G169), .B1(new_n324), .B2(new_n325), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  AND2_X1   g0139(.A1(new_n331), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n293), .A2(new_n296), .A3(new_n340), .ZN(new_n341));
  OR2_X1    g0141(.A1(new_n341), .A2(KEYINPUT68), .ZN(new_n342));
  INV_X1    g0142(.A(G226), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n272), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n224), .A2(G1698), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n316), .A2(new_n344), .A3(new_n318), .A4(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(G33), .A2(G97), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n323), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT13), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n285), .A2(new_n269), .A3(G274), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n269), .A2(G238), .A3(new_n352), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n349), .A2(new_n350), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n269), .B1(new_n346), .B2(new_n347), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n351), .A2(new_n353), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT13), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G169), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT14), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n359), .A2(KEYINPUT14), .A3(G169), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n355), .A2(KEYINPUT69), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT69), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n349), .A2(new_n354), .A3(new_n366), .A4(new_n350), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  AND2_X1   g0168(.A1(new_n358), .A2(G179), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n364), .A2(new_n370), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n256), .A2(G50), .B1(G20), .B2(new_n225), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(new_n252), .B2(new_n202), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n247), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT70), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(KEYINPUT70), .B1(new_n373), .B2(new_n247), .ZN(new_n377));
  OR3_X1    g0177(.A1(new_n376), .A2(KEYINPUT11), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n225), .B1(new_n205), .B2(G20), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n262), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT71), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT12), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n261), .A2(new_n225), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n381), .A2(new_n382), .ZN(new_n384));
  AND2_X1   g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n383), .A2(new_n384), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n380), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(KEYINPUT11), .B1(new_n376), .B2(new_n377), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n378), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n371), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g0191(.A(new_n374), .B(new_n375), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n387), .B1(new_n392), .B2(KEYINPUT11), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n365), .A2(new_n367), .A3(G190), .A4(new_n358), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n359), .A2(G200), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n393), .A2(new_n378), .A3(new_n394), .A4(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n391), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n397), .B1(new_n341), .B2(KEYINPUT68), .ZN(new_n398));
  INV_X1    g0198(.A(G169), .ZN(new_n399));
  OR2_X1    g0199(.A1(G223), .A2(G1698), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n343), .A2(G1698), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n316), .A2(new_n400), .A3(new_n318), .A4(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G33), .A2(G87), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n323), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n269), .A2(G232), .A3(new_n352), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n351), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n399), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n269), .B1(new_n402), .B2(new_n403), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n351), .A2(new_n406), .ZN(new_n410));
  NOR3_X1   g0210(.A1(new_n409), .A2(new_n410), .A3(new_n294), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT16), .ZN(new_n413));
  OAI21_X1  g0213(.A(KEYINPUT72), .B1(new_n317), .B2(G33), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT72), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n415), .A2(new_n249), .A3(KEYINPUT3), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(new_n416), .A3(new_n318), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT7), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n418), .A2(G20), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n418), .B1(new_n270), .B2(G20), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n225), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n223), .A2(new_n225), .ZN(new_n423));
  NOR2_X1   g0223(.A1(G58), .A2(G68), .ZN(new_n424));
  OAI21_X1  g0224(.A(G20), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n256), .A2(G159), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n413), .B1(new_n422), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT7), .B1(new_n319), .B2(new_n206), .ZN(new_n429));
  AOI211_X1 g0229(.A(new_n418), .B(G20), .C1(new_n316), .C2(new_n318), .ZN(new_n430));
  OAI21_X1  g0230(.A(G68), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n427), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n431), .A2(KEYINPUT16), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n428), .A2(new_n247), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n205), .A2(G20), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n308), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n437), .A2(new_n262), .B1(new_n261), .B2(new_n253), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n412), .B1(new_n434), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT18), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n438), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n319), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n421), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n427), .B1(new_n444), .B2(G68), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n333), .B1(new_n445), .B2(KEYINPUT16), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n442), .B1(new_n446), .B2(new_n428), .ZN(new_n447));
  OAI21_X1  g0247(.A(KEYINPUT18), .B1(new_n447), .B2(new_n412), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n441), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT73), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT17), .ZN(new_n451));
  INV_X1    g0251(.A(G190), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n405), .A2(new_n452), .A3(new_n407), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n288), .B1(new_n409), .B2(new_n410), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n451), .B1(new_n447), .B2(new_n455), .ZN(new_n456));
  AND4_X1   g0256(.A1(new_n451), .A2(new_n434), .A3(new_n438), .A4(new_n455), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n450), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n434), .A2(new_n438), .A3(new_n455), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT17), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n447), .A2(new_n451), .A3(new_n455), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT73), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n449), .B1(new_n458), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n342), .A2(new_n398), .A3(new_n463), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n205), .B(G45), .C1(new_n278), .C2(KEYINPUT5), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT75), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n279), .A2(G1), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT5), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G41), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n468), .A2(KEYINPUT75), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n278), .A2(KEYINPUT5), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n473), .B(G274), .C1(new_n322), .C2(new_n214), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n468), .A2(new_n470), .A3(new_n473), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n477), .A2(G257), .A3(new_n269), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n218), .A2(G1698), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n480), .A2(new_n316), .A3(new_n318), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT74), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT4), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n480), .A2(new_n316), .A3(new_n318), .A4(KEYINPUT4), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n316), .A2(new_n318), .A3(G250), .A4(G1698), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n482), .B1(new_n481), .B2(new_n483), .ZN(new_n490));
  NOR3_X1   g0290(.A1(new_n485), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n479), .B1(new_n491), .B2(new_n269), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n399), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n476), .A2(new_n478), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n481), .A2(new_n483), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT74), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(new_n497), .A3(new_n484), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n494), .B1(new_n498), .B2(new_n323), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n294), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT6), .ZN(new_n501));
  INV_X1    g0301(.A(G97), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n501), .A2(new_n502), .A3(G107), .ZN(new_n503));
  XNOR2_X1  g0303(.A(G97), .B(G107), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n503), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  OAI22_X1  g0305(.A1(new_n505), .A2(new_n206), .B1(new_n202), .B2(new_n257), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n320), .B1(new_n420), .B2(new_n421), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n247), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n260), .A2(G97), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n205), .A2(G33), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n262), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n509), .B1(new_n512), .B2(G97), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n508), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n493), .A2(new_n500), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n498), .A2(new_n323), .ZN(new_n516));
  AND4_X1   g0316(.A1(KEYINPUT76), .A2(new_n516), .A3(G190), .A4(new_n479), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT76), .B1(new_n499), .B2(G190), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n508), .B(new_n513), .C1(new_n499), .C2(new_n288), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n515), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n469), .A2(G41), .ZN(new_n522));
  OAI211_X1 g0322(.A(G270), .B(new_n269), .C1(new_n465), .C2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n272), .A2(G257), .ZN(new_n524));
  NAND2_X1  g0324(.A1(G264), .A2(G1698), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n316), .A2(new_n318), .A3(new_n524), .A4(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n526), .B(new_n323), .C1(G303), .C2(new_n270), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n476), .A2(new_n523), .A3(new_n527), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n488), .B(new_n206), .C1(G33), .C2(new_n502), .ZN(new_n529));
  INV_X1    g0329(.A(G116), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G20), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n529), .A2(new_n247), .A3(new_n531), .ZN(new_n532));
  XNOR2_X1  g0332(.A(KEYINPUT77), .B(KEYINPUT20), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n261), .A2(new_n530), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n333), .A2(G116), .A3(new_n260), .A4(new_n510), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT77), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n537), .A2(KEYINPUT20), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n529), .A2(new_n247), .A3(new_n538), .A4(new_n531), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n534), .A2(new_n535), .A3(new_n536), .A4(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n528), .A2(new_n540), .A3(KEYINPUT21), .A4(G169), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n540), .B1(new_n528), .B2(G200), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n323), .B1(new_n270), .B2(G303), .ZN(new_n543));
  AND4_X1   g0343(.A1(new_n316), .A2(new_n318), .A3(new_n524), .A4(new_n525), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n474), .B1(new_n467), .B2(new_n471), .ZN(new_n546));
  INV_X1    g0346(.A(new_n523), .ZN(new_n547));
  NOR3_X1   g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G190), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n542), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n528), .A2(new_n540), .A3(G169), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT21), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(G179), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n528), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n540), .ZN(new_n556));
  AND4_X1   g0356(.A1(new_n541), .A2(new_n550), .A3(new_n553), .A4(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT19), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n252), .B2(new_n502), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n270), .A2(new_n206), .A3(G68), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n206), .B1(new_n347), .B2(new_n558), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n219), .A2(new_n502), .A3(new_n320), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n559), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  XNOR2_X1  g0364(.A(KEYINPUT15), .B(G87), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n564), .A2(new_n247), .B1(new_n261), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n565), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n512), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n220), .B1(new_n279), .B2(G1), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n205), .A2(new_n283), .A3(G45), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n269), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n218), .A2(G1698), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(G238), .B2(G1698), .ZN(new_n574));
  OAI22_X1  g0374(.A1(new_n574), .A2(new_n319), .B1(new_n249), .B2(new_n530), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n572), .B1(new_n575), .B2(new_n323), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n566), .A2(new_n568), .B1(new_n294), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(G238), .A2(G1698), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n578), .B1(new_n218), .B2(G1698), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n579), .A2(new_n270), .B1(G33), .B2(G116), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n571), .B1(new_n580), .B2(new_n269), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n399), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n512), .A2(G87), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n566), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n581), .A2(G200), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n576), .A2(G190), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n577), .A2(new_n582), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  OAI211_X1 g0388(.A(G264), .B(new_n269), .C1(new_n465), .C2(new_n522), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT78), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n477), .A2(KEYINPUT78), .A3(G264), .A4(new_n269), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n316), .A2(new_n318), .A3(G250), .A4(new_n272), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n316), .A2(new_n318), .A3(G257), .A4(G1698), .ZN(new_n595));
  NAND2_X1  g0395(.A1(G33), .A2(G294), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n323), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n593), .A2(new_n476), .A3(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n599), .A2(new_n452), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n591), .A2(new_n592), .B1(new_n597), .B2(new_n323), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n288), .B1(new_n601), .B2(new_n476), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT25), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(new_n260), .B2(G107), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n261), .A2(KEYINPUT25), .A3(new_n320), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n512), .A2(G107), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n316), .A2(new_n318), .A3(new_n206), .A4(G87), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT22), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT22), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n270), .A2(new_n611), .A3(new_n206), .A4(G87), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NOR3_X1   g0413(.A1(new_n249), .A2(new_n530), .A3(G20), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT23), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n206), .B2(G107), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n320), .A2(KEYINPUT23), .A3(G20), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n614), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(KEYINPUT24), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT24), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n613), .A2(new_n621), .A3(new_n618), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n608), .B1(new_n623), .B2(new_n247), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n603), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n599), .A2(G179), .ZN(new_n626));
  AOI21_X1  g0426(.A(G169), .B1(new_n601), .B2(new_n476), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n613), .A2(new_n621), .A3(new_n618), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n621), .B1(new_n613), .B2(new_n618), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n247), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n607), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n557), .A2(new_n588), .A3(new_n625), .A4(new_n633), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n464), .A2(new_n521), .A3(new_n634), .ZN(G372));
  NAND3_X1  g0435(.A1(new_n291), .A2(KEYINPUT81), .A3(new_n292), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(KEYINPUT81), .B1(new_n291), .B2(new_n292), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n396), .A2(new_n335), .A3(new_n338), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n391), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n458), .A2(new_n462), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n639), .B1(new_n449), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n571), .A2(KEYINPUT79), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT79), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n269), .A2(new_n569), .A3(new_n570), .A4(new_n646), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n645), .B(new_n647), .C1(new_n580), .C2(new_n269), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n399), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n577), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n553), .A2(new_n556), .A3(new_n541), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n599), .A2(new_n399), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n601), .A2(new_n554), .A3(new_n476), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT80), .B1(new_n624), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT80), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n628), .A2(new_n657), .A3(new_n632), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n652), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n625), .B1(new_n519), .B2(new_n520), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n515), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n648), .A2(G200), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n584), .A2(new_n586), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n515), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n667), .A2(new_n588), .A3(KEYINPUT26), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n651), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n296), .B(new_n644), .C1(new_n464), .C2(new_n669), .ZN(G369));
  INV_X1    g0470(.A(G13), .ZN(new_n671));
  NOR3_X1   g0471(.A1(new_n671), .A2(G1), .A3(G20), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT82), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT27), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n674), .A2(new_n205), .A3(new_n206), .A4(G13), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(KEYINPUT82), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G213), .ZN(new_n679));
  INV_X1    g0479(.A(new_n672), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n679), .B1(new_n680), .B2(KEYINPUT27), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n678), .A2(KEYINPUT83), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(KEYINPUT83), .B1(new_n678), .B2(new_n681), .ZN(new_n683));
  INV_X1    g0483(.A(G343), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n540), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n557), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n652), .A2(new_n540), .A3(new_n685), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G330), .ZN(new_n690));
  XOR2_X1   g0490(.A(new_n690), .B(KEYINPUT84), .Z(new_n691));
  INV_X1    g0491(.A(new_n685), .ZN(new_n692));
  OAI21_X1  g0492(.A(KEYINPUT85), .B1(new_n624), .B2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT85), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n632), .A2(new_n694), .A3(new_n685), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n693), .A2(new_n633), .A3(new_n625), .A4(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n633), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n685), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n691), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n652), .A2(new_n692), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n656), .A2(new_n658), .A3(new_n692), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n700), .A2(new_n705), .ZN(G399));
  INV_X1    g0506(.A(new_n209), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G41), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n562), .A2(G116), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(G1), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n212), .B2(new_n709), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT28), .ZN(new_n713));
  OR3_X1    g0513(.A1(new_n669), .A2(KEYINPUT29), .A3(new_n685), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n634), .A2(new_n521), .A3(new_n685), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT30), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n548), .A2(G179), .A3(new_n601), .A4(new_n576), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n717), .B1(new_n718), .B2(new_n492), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n601), .A2(new_n576), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n720), .A2(new_n499), .A3(KEYINPUT30), .A4(new_n555), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n528), .A2(new_n648), .A3(new_n294), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(new_n492), .A3(new_n599), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n719), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n685), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT31), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n724), .A2(KEYINPUT31), .A3(new_n685), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n716), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G330), .ZN(new_n732));
  INV_X1    g0532(.A(new_n663), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT26), .B1(new_n733), .B2(new_n515), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n667), .A2(new_n588), .A3(new_n665), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n734), .A2(new_n735), .A3(new_n650), .ZN(new_n736));
  INV_X1    g0536(.A(new_n521), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n625), .A2(new_n650), .A3(new_n663), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n737), .B(new_n738), .C1(new_n652), .C2(new_n697), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n739), .A2(KEYINPUT86), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(KEYINPUT86), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n736), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(KEYINPUT29), .B1(new_n742), .B2(new_n685), .ZN(new_n743));
  AND3_X1   g0543(.A1(new_n714), .A2(new_n732), .A3(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n713), .B1(new_n744), .B2(G1), .ZN(G364));
  INV_X1    g0545(.A(new_n691), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n671), .A2(G20), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G45), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n709), .A2(G1), .A3(new_n748), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n746), .B(new_n749), .C1(G330), .C2(new_n689), .ZN(new_n750));
  INV_X1    g0550(.A(new_n749), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n209), .A2(new_n270), .ZN(new_n752));
  INV_X1    g0552(.A(G355), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n752), .A2(new_n753), .B1(G116), .B2(new_n209), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n707), .A2(new_n270), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n756), .B1(new_n279), .B2(new_n213), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n241), .A2(G45), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n754), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G13), .A2(G33), .ZN(new_n760));
  XOR2_X1   g0560(.A(new_n760), .B(KEYINPUT87), .Z(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n214), .B1(G20), .B2(new_n399), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n751), .B1(new_n759), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n294), .A2(new_n206), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G200), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n452), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT88), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n206), .A2(G179), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n771), .A2(G190), .A3(G200), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n319), .B1(new_n773), .B2(G87), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n769), .A2(G50), .B1(new_n770), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n768), .A2(G190), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n775), .B1(new_n770), .B2(new_n774), .C1(new_n225), .C2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n452), .A2(G200), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n767), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G190), .A2(G200), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n767), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI22_X1  g0584(.A1(G58), .A2(new_n781), .B1(new_n784), .B2(G77), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT32), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n771), .A2(new_n782), .ZN(new_n787));
  INV_X1    g0587(.A(G159), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n779), .A2(new_n554), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G20), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n786), .A2(new_n789), .B1(new_n791), .B2(G97), .ZN(new_n792));
  INV_X1    g0592(.A(new_n789), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n771), .A2(new_n452), .A3(G200), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n793), .A2(KEYINPUT32), .B1(G107), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n785), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G311), .A2(new_n784), .B1(new_n781), .B2(G322), .ZN(new_n798));
  INV_X1    g0598(.A(G283), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n794), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n787), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n270), .B(new_n800), .C1(G329), .C2(new_n801), .ZN(new_n802));
  AOI22_X1  g0602(.A1(G303), .A2(new_n773), .B1(new_n791), .B2(G294), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n798), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n769), .A2(G326), .ZN(new_n805));
  XOR2_X1   g0605(.A(KEYINPUT33), .B(G317), .Z(new_n806));
  OAI21_X1  g0606(.A(new_n805), .B1(new_n777), .B2(new_n806), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n778), .A2(new_n797), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n766), .B1(new_n808), .B2(new_n763), .ZN(new_n809));
  INV_X1    g0609(.A(new_n762), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n809), .B1(new_n689), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n750), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(G396));
  NAND2_X1  g0613(.A1(new_n335), .A2(new_n685), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT91), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n339), .B2(new_n692), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n335), .A2(new_n338), .A3(new_n685), .A4(KEYINPUT91), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n340), .A2(new_n814), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n669), .B2(new_n685), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n818), .A2(new_n685), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n819), .B1(new_n669), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n751), .B1(new_n822), .B2(new_n732), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n732), .B2(new_n822), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n763), .A2(new_n760), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n749), .B1(new_n202), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n818), .ZN(new_n827));
  INV_X1    g0627(.A(G311), .ZN(new_n828));
  INV_X1    g0628(.A(new_n791), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n319), .B1(new_n787), .B2(new_n828), .C1(new_n829), .C2(new_n502), .ZN(new_n830));
  INV_X1    g0630(.A(G294), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n530), .A2(new_n783), .B1(new_n780), .B2(new_n831), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n219), .A2(new_n794), .B1(new_n772), .B2(new_n320), .ZN(new_n833));
  NOR3_X1   g0633(.A1(new_n830), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(G303), .ZN(new_n835));
  INV_X1    g0635(.A(new_n769), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n777), .A2(KEYINPUT89), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n777), .A2(KEYINPUT89), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n834), .B1(new_n835), .B2(new_n836), .C1(new_n839), .C2(new_n799), .ZN(new_n840));
  AOI22_X1  g0640(.A1(G143), .A2(new_n781), .B1(new_n784), .B2(G159), .ZN(new_n841));
  INV_X1    g0641(.A(G137), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n841), .B1(new_n836), .B2(new_n842), .C1(new_n255), .C2(new_n777), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT34), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(G132), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n270), .B1(new_n787), .B2(new_n846), .C1(new_n263), .C2(new_n772), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n829), .A2(new_n223), .B1(new_n794), .B2(new_n225), .ZN(new_n848));
  OR3_X1    g0648(.A1(new_n845), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n843), .A2(new_n844), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n840), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(KEYINPUT90), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n763), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n851), .A2(KEYINPUT90), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n826), .B1(new_n761), .B2(new_n827), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n824), .A2(new_n855), .ZN(G384));
  INV_X1    g0656(.A(new_n505), .ZN(new_n857));
  OR2_X1    g0657(.A1(new_n857), .A2(KEYINPUT35), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(KEYINPUT35), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n858), .A2(G116), .A3(new_n215), .A4(new_n859), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT36), .Z(new_n861));
  OAI211_X1 g0661(.A(new_n213), .B(G77), .C1(new_n223), .C2(new_n225), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n263), .A2(G68), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n205), .B(G13), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n339), .A2(new_n685), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT26), .B1(new_n661), .B2(new_n663), .ZN(new_n867));
  INV_X1    g0667(.A(new_n668), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n650), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n866), .B1(new_n869), .B2(new_n820), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n434), .A2(new_n438), .ZN(new_n872));
  INV_X1    g0672(.A(new_n412), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n682), .A2(new_n683), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT37), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n874), .A2(new_n876), .A3(new_n877), .A4(new_n459), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n433), .A2(new_n247), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n445), .A2(KEYINPUT16), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n438), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n873), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n875), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n882), .A2(new_n883), .A3(new_n459), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n878), .B1(new_n884), .B2(new_n877), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n463), .B2(new_n883), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI211_X1 g0688(.A(KEYINPUT38), .B(new_n885), .C1(new_n463), .C2(new_n883), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n390), .A2(new_n685), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n362), .A2(new_n363), .B1(new_n368), .B2(new_n369), .ZN(new_n892));
  INV_X1    g0692(.A(new_n390), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n396), .B(new_n891), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n371), .A2(new_n390), .A3(new_n685), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n871), .A2(new_n890), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n440), .B1(new_n872), .B2(new_n873), .ZN(new_n898));
  AOI211_X1 g0698(.A(KEYINPUT18), .B(new_n412), .C1(new_n434), .C2(new_n438), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n897), .B1(new_n900), .B2(new_n875), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n890), .A2(KEYINPUT39), .ZN(new_n902));
  XOR2_X1   g0702(.A(KEYINPUT92), .B(KEYINPUT38), .Z(new_n903));
  AND3_X1   g0703(.A1(new_n434), .A2(new_n438), .A3(new_n455), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n904), .A2(new_n439), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n905), .A2(KEYINPUT93), .A3(KEYINPUT37), .A4(new_n876), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n874), .A2(new_n876), .A3(new_n459), .ZN(new_n907));
  INV_X1    g0707(.A(new_n875), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(new_n434), .B2(new_n438), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT37), .B1(new_n909), .B2(KEYINPUT93), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n906), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n460), .A2(new_n461), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n876), .B1(new_n900), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n903), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n889), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT94), .B1(new_n916), .B2(KEYINPUT39), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n902), .A2(new_n917), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n916), .A2(KEYINPUT94), .A3(KEYINPUT39), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n391), .A2(new_n685), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n901), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n464), .B1(new_n714), .B2(new_n743), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n644), .A2(new_n296), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n924), .B(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(G330), .ZN(new_n929));
  INV_X1    g0729(.A(new_n464), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n731), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n818), .B1(new_n894), .B2(new_n895), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n715), .B2(new_n729), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n890), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT40), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n934), .A2(KEYINPUT95), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT95), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n933), .B(new_n940), .C1(new_n715), .C2(new_n729), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n939), .A2(new_n916), .A3(KEYINPUT40), .A4(new_n941), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n938), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n929), .B1(new_n932), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n932), .B2(new_n943), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n928), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n205), .B2(new_n747), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n928), .A2(new_n945), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n865), .B1(new_n947), .B2(new_n948), .ZN(G367));
  AND2_X1   g0749(.A1(new_n755), .A2(new_n237), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n764), .B1(new_n209), .B2(new_n565), .ZN(new_n951));
  OR3_X1    g0751(.A1(new_n650), .A2(new_n584), .A3(new_n692), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n663), .B(new_n650), .C1(new_n584), .C2(new_n692), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n751), .B1(new_n950), .B2(new_n951), .C1(new_n954), .C2(new_n810), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n772), .A2(new_n530), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT46), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n270), .B1(new_n801), .B2(G317), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n958), .B1(new_n502), .B2(new_n794), .C1(new_n780), .C2(new_n835), .ZN(new_n959));
  AOI211_X1 g0759(.A(new_n957), .B(new_n959), .C1(G311), .C2(new_n769), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n783), .A2(new_n799), .B1(new_n829), .B2(new_n320), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT100), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n960), .B(new_n962), .C1(new_n831), .C2(new_n839), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n270), .B1(new_n787), .B2(new_n842), .C1(new_n202), .C2(new_n794), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n829), .A2(new_n225), .B1(new_n772), .B2(new_n223), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n964), .B(new_n965), .C1(G150), .C2(new_n781), .ZN(new_n966));
  INV_X1    g0766(.A(G143), .ZN(new_n967));
  INV_X1    g0767(.A(new_n839), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n968), .A2(G159), .B1(G50), .B2(new_n784), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n966), .B1(new_n967), .B2(new_n836), .C1(new_n969), .C2(KEYINPUT101), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n969), .A2(KEYINPUT101), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n963), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT47), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n763), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(new_n972), .B2(new_n973), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n955), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n514), .A2(new_n685), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n737), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n667), .A2(new_n685), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n982), .A2(new_n702), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT42), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n982), .B(KEYINPUT96), .Z(new_n985));
  AOI21_X1  g0785(.A(new_n667), .B1(new_n985), .B2(new_n697), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n984), .B1(new_n986), .B2(new_n685), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n700), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n990), .A2(new_n985), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT97), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n992), .A2(new_n994), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n989), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n992), .A2(new_n994), .ZN(new_n999));
  INV_X1    g0799(.A(new_n989), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n999), .A2(new_n1000), .A3(new_n995), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n748), .A2(G1), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT98), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n982), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1004), .B(KEYINPUT44), .C1(new_n1005), .C2(new_n705), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(KEYINPUT44), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1004), .A2(KEYINPUT44), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n982), .A2(new_n704), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n982), .A2(new_n704), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT45), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1013), .A2(new_n990), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1013), .A2(new_n990), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n696), .A2(new_n698), .A3(new_n701), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1018), .B(new_n702), .C1(new_n691), .C2(KEYINPUT99), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n691), .A2(KEYINPUT99), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1019), .B(new_n1020), .Z(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n744), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n744), .B1(new_n1017), .B2(new_n1022), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n708), .B(KEYINPUT41), .Z(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1003), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n978), .B1(new_n1002), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(KEYINPUT102), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT102), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1029), .B(new_n978), .C1(new_n1002), .C2(new_n1026), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(G387));
  INV_X1    g0832(.A(new_n1022), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1033), .A2(new_n709), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n744), .B2(new_n1021), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1021), .A2(new_n1003), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G303), .A2(new_n784), .B1(new_n781), .B2(G317), .ZN(new_n1037));
  INV_X1    g0837(.A(G322), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1037), .B1(new_n1038), .B2(new_n836), .C1(new_n839), .C2(new_n828), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT48), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G294), .A2(new_n773), .B1(new_n791), .B2(G283), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT49), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1046), .A2(KEYINPUT104), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(KEYINPUT104), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n794), .A2(new_n530), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n270), .B(new_n1049), .C1(G326), .C2(new_n801), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1047), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n263), .A2(new_n780), .B1(new_n783), .B2(new_n225), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n270), .B1(new_n787), .B2(new_n255), .C1(new_n502), .C2(new_n794), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n829), .A2(new_n565), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n772), .A2(new_n202), .ZN(new_n1055));
  NOR4_X1   g0855(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1056), .B1(new_n788), .B2(new_n836), .C1(new_n253), .C2(new_n777), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n975), .B1(new_n1051), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n710), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n279), .B1(new_n225), .B2(new_n202), .C1(new_n1059), .C2(KEYINPUT103), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(KEYINPUT103), .B2(new_n1059), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n253), .A2(G50), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT50), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n756), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n234), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1064), .B1(new_n1065), .B2(new_n279), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1066), .B1(G107), .B2(new_n209), .C1(new_n710), .C2(new_n752), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n749), .B1(new_n1067), .B2(new_n764), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n699), .B2(new_n810), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1035), .B(new_n1036), .C1(new_n1058), .C2(new_n1069), .ZN(G393));
  INV_X1    g0870(.A(new_n1017), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n709), .B1(new_n1071), .B2(new_n1033), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n1033), .B2(new_n1071), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1017), .A2(KEYINPUT105), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT105), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1015), .A2(new_n1016), .A3(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1074), .A2(new_n1003), .A3(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n764), .B1(new_n502), .B2(new_n209), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n756), .A2(new_n244), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n751), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n769), .A2(G317), .B1(new_n781), .B2(G311), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT52), .Z(new_n1082));
  OAI221_X1 g0882(.A(new_n319), .B1(new_n787), .B2(new_n1038), .C1(new_n320), .C2(new_n794), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n829), .A2(new_n530), .B1(new_n772), .B2(new_n799), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n1083), .B(new_n1084), .C1(G294), .C2(new_n784), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1082), .B(new_n1085), .C1(new_n835), .C2(new_n839), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT106), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n769), .A2(G150), .B1(new_n781), .B2(G159), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT51), .Z(new_n1090));
  OAI221_X1 g0890(.A(new_n270), .B1(new_n787), .B2(new_n967), .C1(new_n219), .C2(new_n794), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n829), .A2(new_n202), .B1(new_n772), .B2(new_n225), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1091), .B(new_n1092), .C1(new_n308), .C2(new_n784), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1090), .B(new_n1093), .C1(new_n263), .C2(new_n839), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1088), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1080), .B1(new_n1096), .B2(new_n763), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n985), .B2(new_n810), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n1077), .A2(KEYINPUT107), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(KEYINPUT107), .B1(new_n1077), .B2(new_n1098), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1073), .B1(new_n1099), .B2(new_n1100), .ZN(G390));
  INV_X1    g0901(.A(new_n896), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n922), .B1(new_n870), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT108), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g0905(.A(KEYINPUT108), .B(new_n922), .C1(new_n870), .C2(new_n1102), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1105), .A2(new_n920), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n740), .A2(new_n741), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n736), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n685), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n866), .B1(new_n1110), .B2(new_n827), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n922), .B(new_n916), .C1(new_n1111), .C2(new_n1102), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n934), .A2(new_n929), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n1107), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1114), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n1003), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n769), .A2(G283), .B1(new_n784), .B2(G97), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n839), .B2(new_n320), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n1120), .B(KEYINPUT113), .Z(new_n1121));
  OAI22_X1  g0921(.A1(new_n780), .A2(new_n530), .B1(new_n829), .B2(new_n202), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT115), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n319), .B1(new_n772), .B2(new_n219), .ZN(new_n1124));
  XOR2_X1   g0924(.A(new_n1124), .B(KEYINPUT114), .Z(new_n1125));
  OAI22_X1  g0925(.A1(new_n794), .A2(new_n225), .B1(new_n787), .B2(new_n831), .ZN(new_n1126));
  NOR4_X1   g0926(.A1(new_n1121), .A2(new_n1123), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT54), .B(G143), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n783), .A2(new_n1128), .B1(new_n829), .B2(new_n788), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(new_n968), .B2(G137), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT112), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n773), .A2(G150), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT53), .ZN(new_n1133));
  INV_X1    g0933(.A(G128), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n836), .A2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n780), .A2(new_n846), .ZN(new_n1136));
  INV_X1    g0936(.A(G125), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n270), .B1(new_n787), .B2(new_n1137), .C1(new_n263), .C2(new_n794), .ZN(new_n1138));
  OR3_X1    g0938(.A1(new_n1135), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1139));
  NOR3_X1   g0939(.A1(new_n1131), .A2(new_n1133), .A3(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n763), .B1(new_n1127), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n825), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1141), .B(new_n751), .C1(new_n308), .C2(new_n1142), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT116), .Z(new_n1144));
  NOR3_X1   g0944(.A1(new_n918), .A2(new_n761), .A3(new_n919), .ZN(new_n1145));
  OR2_X1    g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1118), .A2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n464), .A2(new_n732), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n927), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT109), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NOR4_X1   g0952(.A1(new_n925), .A2(new_n1151), .A3(new_n926), .A4(new_n1148), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT110), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n818), .B1(new_n732), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n1156), .B2(new_n732), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n1102), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1155), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1102), .B1(new_n732), .B2(new_n818), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n1114), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n871), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1152), .A2(new_n1154), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT111), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n709), .B1(new_n1167), .B2(new_n1117), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1165), .B(new_n1166), .C1(new_n1116), .C2(new_n1115), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1147), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(G378));
  INV_X1    g0971(.A(new_n924), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n875), .A2(new_n266), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT118), .Z(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n639), .B2(new_n296), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n638), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1179), .A2(new_n296), .A3(new_n636), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1180), .A2(new_n1176), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1174), .B1(new_n1178), .B2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n639), .A2(new_n296), .A3(new_n1177), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1180), .A2(new_n1176), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1183), .A2(new_n1184), .A3(new_n1173), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1182), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n943), .A2(new_n1186), .A3(G330), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n934), .B1(new_n888), .B2(new_n889), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n942), .B(G330), .C1(KEYINPUT40), .C2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(KEYINPUT119), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT119), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n938), .A2(new_n1191), .A3(G330), .A4(new_n942), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1186), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT120), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1187), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  AOI211_X1 g0995(.A(KEYINPUT120), .B(new_n1186), .C1(new_n1190), .C2(new_n1192), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1172), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1186), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(KEYINPUT120), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1201), .A2(new_n924), .A3(new_n1202), .A4(new_n1187), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1197), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1107), .A2(new_n1112), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n1113), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1107), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1206), .A2(new_n1207), .A3(new_n1164), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT121), .ZN(new_n1209));
  AOI21_X1  g1009(.A(KEYINPUT109), .B1(new_n927), .B2(new_n1149), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1210), .A2(new_n1153), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n1208), .A2(new_n1209), .A3(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1209), .B1(new_n1208), .B2(new_n1211), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1204), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT57), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n709), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  OAI211_X1 g1016(.A(KEYINPUT57), .B(new_n1204), .C1(new_n1212), .C2(new_n1213), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n751), .B1(G50), .B2(new_n1142), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT117), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n263), .B1(G33), .B2(G41), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(new_n319), .B2(new_n278), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G97), .A2(new_n776), .B1(new_n769), .B2(G116), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n829), .A2(new_n225), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n278), .B(new_n319), .C1(new_n787), .C2(new_n799), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n794), .A2(new_n223), .ZN(new_n1226));
  NOR4_X1   g1026(.A1(new_n1224), .A2(new_n1225), .A3(new_n1055), .A4(new_n1226), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(G107), .A2(new_n781), .B1(new_n784), .B2(new_n567), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1223), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT58), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1222), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n791), .A2(G150), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1232), .B1(new_n772), .B2(new_n1128), .C1(new_n780), .C2(new_n1134), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n1137), .A2(new_n836), .B1(new_n777), .B2(new_n846), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n1233), .B(new_n1234), .C1(G137), .C2(new_n784), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(KEYINPUT59), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n795), .A2(G159), .ZN(new_n1238));
  AOI211_X1 g1038(.A(G33), .B(G41), .C1(new_n801), .C2(G124), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1236), .A2(KEYINPUT59), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1231), .B1(new_n1230), .B2(new_n1229), .C1(new_n1240), .C2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1220), .B1(new_n1242), .B2(new_n763), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n1186), .B2(new_n761), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(new_n1204), .B2(new_n1003), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1218), .A2(new_n1246), .ZN(G375));
  AOI22_X1  g1047(.A1(new_n1155), .A2(new_n1159), .B1(new_n871), .B2(new_n1162), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n1210), .B2(new_n1153), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1165), .A2(new_n1025), .A3(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n751), .B1(G68), .B2(new_n1142), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n829), .A2(new_n263), .B1(new_n1134), .B2(new_n787), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n842), .A2(new_n780), .B1(new_n783), .B2(new_n255), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n1252), .B(new_n1253), .C1(G159), .C2(new_n773), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n270), .B1(new_n794), .B2(new_n223), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n769), .A2(G132), .B1(KEYINPUT123), .B2(new_n1255), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1254), .B(new_n1256), .C1(KEYINPUT123), .C2(new_n1255), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n839), .A2(new_n1128), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n839), .A2(new_n530), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n319), .B1(new_n787), .B2(new_n835), .C1(new_n202), .C2(new_n794), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n1260), .B(new_n1054), .C1(G97), .C2(new_n773), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(G107), .A2(new_n784), .B1(new_n781), .B2(G283), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1261), .B(new_n1262), .C1(new_n831), .C2(new_n836), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n1257), .A2(new_n1258), .B1(new_n1259), .B2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1251), .B1(new_n1264), .B2(new_n763), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n760), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1265), .B1(new_n896), .B2(new_n1266), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1003), .B(KEYINPUT122), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1267), .B1(new_n1248), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1250), .A2(new_n1270), .ZN(G381));
  OR3_X1    g1071(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1272));
  NOR3_X1   g1072(.A1(G378), .A2(new_n1272), .A3(G381), .ZN(new_n1273));
  AOI21_X1  g1073(.A(G390), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1273), .A2(new_n1218), .A3(new_n1246), .A4(new_n1274), .ZN(G407));
  NOR2_X1   g1075(.A1(new_n679), .A2(G343), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1170), .A2(new_n1276), .ZN(new_n1277));
  OAI211_X1 g1077(.A(G407), .B(G213), .C1(G375), .C2(new_n1277), .ZN(G409));
  INV_X1    g1078(.A(KEYINPUT62), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(G384), .A2(KEYINPUT124), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1280), .A2(new_n1269), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT60), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1165), .B(new_n708), .C1(new_n1249), .C2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT60), .B1(new_n1284), .B2(new_n1248), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1281), .B1(new_n1283), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(G384), .A2(KEYINPUT124), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(new_n1286), .B(new_n1287), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1197), .A2(new_n1203), .ZN(new_n1289));
  NOR3_X1   g1089(.A1(new_n1115), .A2(new_n1116), .A3(new_n1248), .ZN(new_n1290));
  OAI21_X1  g1090(.A(KEYINPUT121), .B1(new_n1290), .B2(new_n1284), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1208), .A2(new_n1209), .A3(new_n1211), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1289), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n708), .B1(new_n1293), .B2(KEYINPUT57), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1217), .ZN(new_n1295));
  OAI211_X1 g1095(.A(G378), .B(new_n1246), .C1(new_n1294), .C2(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1025), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1289), .B1(new_n1297), .B2(new_n1268), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1170), .B1(new_n1298), .B2(new_n1245), .ZN(new_n1299));
  AOI211_X1 g1099(.A(new_n1276), .B(new_n1288), .C1(new_n1296), .C2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1279), .B1(new_n1300), .B2(KEYINPUT126), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1276), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1246), .ZN(new_n1303));
  AOI211_X1 g1103(.A(new_n1303), .B(new_n1170), .C1(new_n1216), .C2(new_n1217), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1297), .A2(new_n1268), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1204), .ZN(new_n1306));
  AOI21_X1  g1106(.A(G378), .B1(new_n1306), .B2(new_n1244), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1302), .B1(new_n1304), .B2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(G2897), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1302), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1288), .A2(new_n1310), .ZN(new_n1311));
  AND3_X1   g1111(.A1(new_n1286), .A2(KEYINPUT124), .A3(G384), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1281), .B(new_n1287), .C1(new_n1283), .C2(new_n1285), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  OAI22_X1  g1114(.A1(new_n1312), .A2(new_n1314), .B1(new_n1309), .B2(new_n1302), .ZN(new_n1315));
  AND2_X1   g1115(.A1(new_n1311), .A2(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(KEYINPUT61), .B1(new_n1308), .B2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1288), .ZN(new_n1318));
  OAI211_X1 g1118(.A(new_n1302), .B(new_n1318), .C1(new_n1304), .C2(new_n1307), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT126), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1319), .A2(new_n1320), .A3(KEYINPUT62), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1301), .A2(new_n1317), .A3(new_n1321), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(G393), .B(new_n812), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(G390), .A2(new_n1027), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1325), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1324), .B1(new_n1274), .B2(new_n1326), .ZN(new_n1327));
  OR2_X1    g1127(.A1(G390), .A2(new_n1027), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1328), .A2(new_n1323), .A3(new_n1325), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1327), .A2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1322), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT61), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1276), .B1(new_n1296), .B2(new_n1299), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1311), .A2(new_n1315), .ZN(new_n1335));
  OAI211_X1 g1135(.A(new_n1330), .B(new_n1333), .C1(new_n1334), .C2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1300), .A2(KEYINPUT63), .ZN(new_n1338));
  NOR3_X1   g1138(.A1(new_n1300), .A2(KEYINPUT125), .A3(KEYINPUT63), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT125), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT63), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1340), .B1(new_n1319), .B2(new_n1341), .ZN(new_n1342));
  OAI211_X1 g1142(.A(new_n1337), .B(new_n1338), .C1(new_n1339), .C2(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1332), .A2(new_n1343), .ZN(G405));
  AOI21_X1  g1144(.A(G378), .B1(new_n1218), .B2(new_n1246), .ZN(new_n1345));
  NOR2_X1   g1145(.A1(new_n1345), .A2(new_n1304), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1318), .A2(KEYINPUT127), .ZN(new_n1347));
  OR2_X1    g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1349));
  AND3_X1   g1149(.A1(new_n1348), .A2(new_n1331), .A3(new_n1349), .ZN(new_n1350));
  AOI21_X1  g1150(.A(new_n1331), .B1(new_n1348), .B2(new_n1349), .ZN(new_n1351));
  NOR2_X1   g1151(.A1(new_n1350), .A2(new_n1351), .ZN(G402));
endmodule


