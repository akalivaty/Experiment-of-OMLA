//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 0 1 0 1 0 1 1 1 1 0 0 0 1 1 0 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 0 1 1 0 0 1 1 0 1 1 1 0 1 0 0 1 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n799, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n999, new_n1000, new_n1001, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1044,
    new_n1045, new_n1046;
  INV_X1    g000(.A(KEYINPUT68), .ZN(new_n202));
  INV_X1    g001(.A(G113gat), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G120gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(G120gat), .ZN(new_n205));
  INV_X1    g004(.A(G120gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n206), .A2(KEYINPUT68), .A3(G113gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n204), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT69), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND4_X1  g009(.A1(new_n204), .A2(new_n207), .A3(KEYINPUT69), .A4(new_n205), .ZN(new_n211));
  INV_X1    g010(.A(G134gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G127gat), .ZN(new_n213));
  INV_X1    g012(.A(G127gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G134gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n213), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n210), .A2(new_n211), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n206), .A2(G113gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(new_n205), .ZN(new_n221));
  AOI22_X1  g020(.A1(new_n221), .A2(new_n216), .B1(new_n213), .B2(new_n215), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n219), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT82), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n217), .B1(new_n208), .B2(new_n209), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n222), .B1(new_n227), .B2(new_n211), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT82), .ZN(new_n229));
  OR2_X1    g028(.A1(KEYINPUT79), .A2(KEYINPUT2), .ZN(new_n230));
  NAND2_X1  g029(.A1(KEYINPUT79), .A2(KEYINPUT2), .ZN(new_n231));
  INV_X1    g030(.A(G141gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n232), .A2(G148gat), .ZN(new_n233));
  INV_X1    g032(.A(G148gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n234), .A2(G141gat), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n230), .B(new_n231), .C1(new_n233), .C2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G162gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G155gat), .ZN(new_n238));
  INV_X1    g037(.A(G155gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G162gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n236), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n241), .ZN(new_n243));
  AND2_X1   g042(.A1(KEYINPUT80), .A2(G141gat), .ZN(new_n244));
  NOR2_X1   g043(.A1(KEYINPUT80), .A2(G141gat), .ZN(new_n245));
  NOR3_X1   g044(.A1(new_n244), .A2(new_n245), .A3(new_n234), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n243), .B1(new_n246), .B2(new_n233), .ZN(new_n247));
  AND2_X1   g046(.A1(KEYINPUT81), .A2(G162gat), .ZN(new_n248));
  NOR2_X1   g047(.A1(KEYINPUT81), .A2(G162gat), .ZN(new_n249));
  OAI21_X1  g048(.A(G155gat), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n250), .A2(KEYINPUT2), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n242), .B1(new_n247), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n250), .A2(KEYINPUT2), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT80), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(new_n232), .ZN(new_n256));
  NAND2_X1  g055(.A1(KEYINPUT80), .A2(G141gat), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n256), .A2(G148gat), .A3(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n233), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n254), .A2(new_n260), .A3(new_n243), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT3), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n261), .A2(new_n262), .A3(new_n242), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n226), .A2(new_n229), .A3(new_n253), .A4(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT83), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI211_X1 g065(.A(new_n225), .B(new_n222), .C1(new_n227), .C2(new_n211), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT82), .B1(new_n219), .B2(new_n223), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n261), .A2(new_n262), .A3(new_n242), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n262), .B1(new_n261), .B2(new_n242), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n269), .A2(new_n272), .A3(KEYINPUT83), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n266), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n275));
  NAND2_X1  g074(.A1(G225gat), .A2(G233gat), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n241), .B1(new_n258), .B2(new_n259), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n277), .A2(new_n254), .B1(new_n241), .B2(new_n236), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n228), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n228), .A2(KEYINPUT4), .A3(new_n278), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n274), .A2(new_n275), .A3(new_n276), .A4(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n276), .ZN(new_n286));
  AOI211_X1 g085(.A(new_n286), .B(new_n283), .C1(new_n266), .C2(new_n273), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n226), .A2(new_n229), .A3(new_n252), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(new_n279), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n275), .B1(new_n289), .B2(new_n286), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n285), .B1(new_n287), .B2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G1gat), .B(G29gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(KEYINPUT0), .ZN(new_n294));
  XNOR2_X1  g093(.A(G57gat), .B(G85gat), .ZN(new_n295));
  XOR2_X1   g094(.A(new_n294), .B(new_n295), .Z(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n292), .A2(KEYINPUT6), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT84), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n264), .A2(new_n265), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT83), .B1(new_n269), .B2(new_n272), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n276), .B(new_n284), .C1(new_n301), .C2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(new_n290), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n296), .B1(new_n304), .B2(new_n285), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n305), .A2(KEYINPUT84), .A3(KEYINPUT6), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n300), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(G226gat), .A2(G233gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G183gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT27), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT27), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G183gat), .ZN(new_n314));
  INV_X1    g113(.A(G190gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n312), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n310), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT27), .B(G183gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n317), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(new_n315), .A3(new_n320), .ZN(new_n321));
  AOI22_X1  g120(.A1(new_n318), .A2(new_n321), .B1(G183gat), .B2(G190gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT64), .ZN(new_n323));
  INV_X1    g122(.A(G169gat), .ZN(new_n324));
  INV_X1    g123(.A(G176gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT26), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT67), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT67), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n326), .A2(new_n331), .A3(new_n327), .A4(new_n328), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n327), .B1(new_n324), .B2(new_n325), .ZN(new_n333));
  NOR2_X1   g132(.A1(G169gat), .A2(G176gat), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n330), .A2(new_n332), .A3(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(G183gat), .A2(G190gat), .ZN(new_n338));
  AND2_X1   g137(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n338), .B1(new_n339), .B2(G190gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(G183gat), .A2(G190gat), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT24), .ZN(new_n342));
  AND3_X1   g141(.A1(new_n341), .A2(KEYINPUT65), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT65), .B1(new_n341), .B2(new_n342), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n340), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n326), .A2(KEYINPUT23), .A3(new_n328), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT25), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT23), .B1(new_n324), .B2(new_n325), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n347), .B1(new_n348), .B2(new_n335), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n345), .A2(new_n346), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n334), .A2(KEYINPUT23), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT23), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n352), .B1(G169gat), .B2(G176gat), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n351), .B1(new_n353), .B2(new_n334), .ZN(new_n354));
  AND3_X1   g153(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n356));
  NOR3_X1   g155(.A1(new_n355), .A2(new_n356), .A3(new_n338), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n347), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n322), .A2(new_n337), .B1(new_n350), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n308), .B1(new_n359), .B2(KEYINPUT29), .ZN(new_n360));
  XNOR2_X1  g159(.A(G197gat), .B(G204gat), .ZN(new_n361));
  INV_X1    g160(.A(G218gat), .ZN(new_n362));
  INV_X1    g161(.A(G211gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT74), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT74), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(G211gat), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n362), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT73), .B(KEYINPUT22), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n361), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G211gat), .B(G218gat), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT75), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  OAI221_X1 g172(.A(new_n361), .B1(new_n370), .B2(new_n371), .C1(new_n367), .C2(new_n368), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n316), .A2(new_n317), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n376), .A2(new_n321), .A3(new_n309), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n337), .A2(new_n341), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n350), .A2(new_n358), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n308), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT76), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT76), .ZN(new_n383));
  AOI211_X1 g182(.A(new_n383), .B(new_n308), .C1(new_n378), .C2(new_n379), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n360), .B(new_n375), .C1(new_n382), .C2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n375), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n381), .B1(new_n380), .B2(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n359), .A2(new_n308), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n386), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT37), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n385), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n360), .B(new_n386), .C1(new_n382), .C2(new_n384), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n375), .B1(new_n388), .B2(new_n389), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(KEYINPUT37), .A3(new_n394), .ZN(new_n395));
  XOR2_X1   g194(.A(G8gat), .B(G36gat), .Z(new_n396));
  XNOR2_X1  g195(.A(new_n396), .B(KEYINPUT77), .ZN(new_n397));
  XNOR2_X1  g196(.A(G64gat), .B(G92gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n397), .B(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT78), .ZN(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT88), .B(KEYINPUT38), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n392), .A2(new_n395), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n380), .A2(new_n381), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n375), .B1(new_n360), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n383), .B1(new_n359), .B2(new_n308), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n380), .A2(KEYINPUT76), .A3(new_n381), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n388), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n404), .B1(new_n407), .B2(new_n375), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n399), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n402), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n399), .ZN(new_n411));
  OAI211_X1 g210(.A(KEYINPUT89), .B(new_n411), .C1(new_n408), .C2(new_n391), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT89), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n391), .B1(new_n385), .B2(new_n390), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n413), .B1(new_n414), .B2(new_n399), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n412), .A2(new_n415), .A3(new_n392), .ZN(new_n416));
  INV_X1    g215(.A(new_n401), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n410), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT6), .B1(new_n292), .B2(new_n297), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n304), .A2(new_n296), .A3(new_n285), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n307), .A2(new_n418), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(G228gat), .A2(G233gat), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT29), .B1(new_n278), .B2(new_n262), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n424), .A2(new_n375), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n369), .A2(new_n370), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n363), .A2(G218gat), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n362), .A2(G211gat), .ZN(new_n428));
  OAI221_X1 g227(.A(new_n361), .B1(new_n427), .B2(new_n428), .C1(new_n367), .C2(new_n368), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n426), .A2(new_n429), .A3(new_n387), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n278), .B1(new_n430), .B2(new_n262), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n423), .B1(new_n425), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT29), .B1(new_n373), .B2(new_n374), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n252), .B1(new_n433), .B2(KEYINPUT3), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n263), .A2(new_n387), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n386), .ZN(new_n436));
  INV_X1    g235(.A(new_n423), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n434), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n432), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(G22gat), .ZN(new_n440));
  INV_X1    g239(.A(G22gat), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n432), .A2(new_n441), .A3(new_n438), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT86), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n442), .A2(KEYINPUT85), .ZN(new_n445));
  XNOR2_X1  g244(.A(G78gat), .B(G106gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(KEYINPUT31), .B(G50gat), .ZN(new_n447));
  XOR2_X1   g246(.A(new_n446), .B(new_n447), .Z(new_n448));
  AOI21_X1  g247(.A(new_n444), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n448), .ZN(new_n450));
  AOI211_X1 g249(.A(KEYINPUT86), .B(new_n450), .C1(new_n442), .C2(KEYINPUT85), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n443), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT85), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT29), .B1(new_n369), .B2(new_n370), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT3), .B1(new_n454), .B2(new_n429), .ZN(new_n455));
  OAI22_X1  g254(.A1(new_n455), .A2(new_n278), .B1(new_n424), .B2(new_n375), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n423), .B1(new_n435), .B2(new_n386), .ZN(new_n457));
  AOI22_X1  g256(.A1(new_n456), .A2(new_n423), .B1(new_n457), .B2(new_n434), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n453), .B1(new_n458), .B2(new_n441), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT86), .B1(new_n459), .B2(new_n450), .ZN(new_n460));
  INV_X1    g259(.A(new_n443), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n444), .A3(new_n448), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n452), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n276), .B1(new_n274), .B2(new_n284), .ZN(new_n465));
  XOR2_X1   g264(.A(KEYINPUT87), .B(KEYINPUT39), .Z(new_n466));
  AOI21_X1  g265(.A(new_n297), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT39), .ZN(new_n468));
  INV_X1    g267(.A(new_n279), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n469), .B1(new_n269), .B2(new_n252), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n468), .B1(new_n470), .B2(new_n276), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n283), .B1(new_n266), .B2(new_n273), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n471), .B1(new_n472), .B2(new_n276), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT40), .B1(new_n467), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n284), .B1(new_n301), .B2(new_n302), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n475), .A2(new_n286), .A3(new_n466), .ZN(new_n476));
  AND4_X1   g275(.A1(KEYINPUT40), .A2(new_n476), .A3(new_n473), .A4(new_n296), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT30), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n385), .A2(new_n390), .ZN(new_n480));
  AOI22_X1  g279(.A1(new_n409), .A2(new_n479), .B1(new_n480), .B2(new_n400), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n408), .A2(KEYINPUT30), .A3(new_n399), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n305), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n464), .B1(new_n478), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n422), .A2(new_n484), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n300), .A2(new_n306), .B1(new_n420), .B2(new_n419), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n481), .A2(new_n482), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n464), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n378), .A2(new_n228), .A3(new_n379), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT70), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n380), .A2(new_n224), .ZN(new_n492));
  NAND2_X1  g291(.A1(G227gat), .A2(G233gat), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT70), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n378), .A2(new_n379), .A3(new_n494), .A4(new_n228), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n491), .A2(new_n492), .A3(new_n493), .A4(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT34), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n496), .B(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT32), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n491), .A2(new_n495), .A3(new_n492), .ZN(new_n501));
  INV_X1    g300(.A(new_n493), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT33), .B1(new_n501), .B2(new_n502), .ZN(new_n504));
  XOR2_X1   g303(.A(G15gat), .B(G43gat), .Z(new_n505));
  XNOR2_X1  g304(.A(G71gat), .B(G99gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NOR3_X1   g307(.A1(new_n503), .A2(new_n504), .A3(new_n508), .ZN(new_n509));
  AOI221_X4 g308(.A(new_n500), .B1(KEYINPUT33), .B2(new_n507), .C1(new_n501), .C2(new_n502), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n499), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n501), .A2(new_n502), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT33), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n508), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n503), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n503), .B1(new_n504), .B2(new_n508), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n498), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n511), .A2(KEYINPUT71), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT71), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n520), .B(new_n499), .C1(new_n509), .C2(new_n510), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT36), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n511), .A2(KEYINPUT72), .A3(new_n518), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT36), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT72), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n516), .A2(new_n526), .A3(new_n498), .A4(new_n517), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n524), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  AND2_X1   g327(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT35), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n487), .B1(new_n307), .B2(new_n421), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n464), .B1(new_n521), .B2(new_n519), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AND4_X1   g332(.A1(KEYINPUT84), .A2(new_n292), .A3(KEYINPUT6), .A4(new_n297), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT84), .B1(new_n305), .B2(KEYINPUT6), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n421), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n524), .A2(new_n527), .ZN(new_n537));
  INV_X1    g336(.A(new_n487), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n452), .A2(new_n530), .A3(new_n463), .ZN(new_n539));
  AND4_X1   g338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  OAI22_X1  g339(.A1(new_n489), .A2(new_n529), .B1(new_n533), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT93), .ZN(new_n543));
  XNOR2_X1  g342(.A(G15gat), .B(G22gat), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n544), .A2(G1gat), .ZN(new_n545));
  INV_X1    g344(.A(G8gat), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT16), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n544), .B1(new_n547), .B2(G1gat), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n546), .B1(new_n545), .B2(new_n548), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n543), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n551), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n553), .A2(KEYINPUT93), .A3(new_n549), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT21), .ZN(new_n556));
  INV_X1    g355(.A(G64gat), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n557), .A2(G57gat), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n557), .A2(G57gat), .ZN(new_n559));
  OAI21_X1  g358(.A(KEYINPUT9), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(G71gat), .A2(G78gat), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT94), .ZN(new_n563));
  INV_X1    g362(.A(G71gat), .ZN(new_n564));
  INV_X1    g363(.A(G78gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n562), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n560), .B(new_n567), .C1(new_n563), .C2(new_n566), .ZN(new_n568));
  NAND2_X1  g367(.A1(KEYINPUT95), .A2(G57gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(G64gat), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT96), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT9), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n561), .B1(new_n566), .B2(new_n572), .ZN(new_n573));
  AND3_X1   g372(.A1(new_n570), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n571), .B1(new_n570), .B2(new_n573), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n568), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n555), .B1(new_n556), .B2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(KEYINPUT98), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n569), .B(new_n557), .ZN(new_n579));
  NOR2_X1   g378(.A1(G71gat), .A2(G78gat), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n562), .B1(KEYINPUT9), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(KEYINPUT96), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n570), .A2(new_n571), .A3(new_n573), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(KEYINPUT21), .B1(new_n584), .B2(new_n568), .ZN(new_n585));
  NAND2_X1  g384(.A1(G231gat), .A2(G233gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G127gat), .B(G155gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT20), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n587), .B(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n578), .B(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G183gat), .B(G211gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  OR2_X1    g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n591), .A2(new_n594), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(KEYINPUT92), .B(KEYINPUT17), .Z(new_n598));
  XNOR2_X1  g397(.A(G43gat), .B(G50gat), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT90), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT15), .ZN(new_n602));
  INV_X1    g401(.A(G43gat), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n603), .A2(KEYINPUT90), .A3(G50gat), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n601), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT91), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n599), .A2(KEYINPUT15), .ZN(new_n607));
  INV_X1    g406(.A(G29gat), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n608), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n609));
  AND2_X1   g408(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n610));
  NOR2_X1   g409(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n609), .B1(new_n612), .B2(G36gat), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n605), .A2(new_n606), .A3(new_n607), .A4(new_n613), .ZN(new_n614));
  OR2_X1    g413(.A1(new_n613), .A2(new_n607), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n613), .A2(new_n607), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n606), .B1(new_n617), .B2(new_n605), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n598), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n605), .A2(new_n607), .A3(new_n613), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(KEYINPUT91), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n621), .A2(KEYINPUT17), .A3(new_n615), .A4(new_n614), .ZN(new_n622));
  NAND2_X1  g421(.A1(G85gat), .A2(G92gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT7), .ZN(new_n624));
  NAND2_X1  g423(.A1(G99gat), .A2(G106gat), .ZN(new_n625));
  INV_X1    g424(.A(G85gat), .ZN(new_n626));
  INV_X1    g425(.A(G92gat), .ZN(new_n627));
  AOI22_X1  g426(.A1(KEYINPUT8), .A2(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  OR2_X1    g428(.A1(G99gat), .A2(G106gat), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n629), .A2(new_n625), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n625), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n624), .A2(new_n632), .A3(new_n628), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n619), .A2(new_n622), .A3(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(G190gat), .B(G218gat), .Z(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n621), .A2(new_n615), .A3(new_n614), .ZN(new_n638));
  INV_X1    g437(.A(new_n634), .ZN(new_n639));
  AND2_X1   g438(.A1(G232gat), .A2(G233gat), .ZN(new_n640));
  AOI22_X1  g439(.A1(new_n638), .A2(new_n639), .B1(KEYINPUT41), .B2(new_n640), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n635), .A2(new_n637), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n637), .B1(new_n635), .B2(new_n641), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n640), .A2(KEYINPUT41), .ZN(new_n644));
  XNOR2_X1  g443(.A(G134gat), .B(G162gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  OR3_X1    g446(.A1(new_n642), .A2(new_n643), .A3(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n647), .B1(new_n642), .B2(new_n643), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n597), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n619), .A2(new_n553), .A3(new_n549), .A4(new_n622), .ZN(new_n653));
  NAND2_X1  g452(.A1(G229gat), .A2(G233gat), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n638), .A2(new_n554), .A3(new_n552), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT18), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n653), .A2(KEYINPUT18), .A3(new_n654), .A4(new_n655), .ZN(new_n659));
  INV_X1    g458(.A(new_n638), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(new_n555), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n655), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n654), .B(KEYINPUT13), .Z(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n658), .A2(new_n659), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(G113gat), .B(G141gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G197gat), .ZN(new_n667));
  XOR2_X1   g466(.A(KEYINPUT11), .B(G169gat), .Z(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT12), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n665), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n658), .A2(new_n670), .A3(new_n659), .A4(new_n664), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n576), .A2(new_n634), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n584), .A2(new_n568), .A3(new_n633), .A4(new_n631), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n675), .A2(new_n676), .A3(KEYINPUT99), .ZN(new_n677));
  INV_X1    g476(.A(G230gat), .ZN(new_n678));
  INV_X1    g477(.A(G233gat), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT99), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n576), .A2(new_n634), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n677), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n683), .A2(KEYINPUT100), .ZN(new_n684));
  INV_X1    g483(.A(new_n680), .ZN(new_n685));
  AOI21_X1  g484(.A(KEYINPUT10), .B1(new_n677), .B2(new_n682), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT10), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n676), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n685), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n683), .A2(KEYINPUT100), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n684), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(G120gat), .B(G148gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(G176gat), .B(G204gat), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n692), .B(new_n693), .Z(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n684), .A2(new_n689), .A3(new_n694), .A4(new_n690), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n652), .A2(new_n674), .A3(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n542), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n486), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(G1gat), .ZN(G1324gat));
  OR2_X1    g502(.A1(new_n542), .A2(new_n700), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n704), .A2(new_n538), .ZN(new_n705));
  XOR2_X1   g504(.A(KEYINPUT16), .B(G8gat), .Z(new_n706));
  AND4_X1   g505(.A1(KEYINPUT101), .A2(new_n705), .A3(KEYINPUT42), .A4(new_n706), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n705), .A2(new_n706), .ZN(new_n708));
  AOI21_X1  g507(.A(KEYINPUT101), .B1(new_n708), .B2(KEYINPUT42), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT42), .B1(new_n705), .B2(new_n546), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n705), .A2(new_n706), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n707), .B1(new_n709), .B2(new_n712), .ZN(G1325gat));
  INV_X1    g512(.A(new_n537), .ZN(new_n714));
  OR3_X1    g513(.A1(new_n704), .A2(G15gat), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n523), .A2(new_n528), .ZN(new_n716));
  OAI21_X1  g515(.A(G15gat), .B1(new_n704), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(G1326gat));
  NAND2_X1  g517(.A1(new_n701), .A2(new_n464), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT102), .ZN(new_n720));
  XOR2_X1   g519(.A(KEYINPUT43), .B(G22gat), .Z(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1327gat));
  INV_X1    g521(.A(new_n464), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n536), .A2(new_n522), .A3(new_n538), .A4(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT35), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n531), .A2(new_n537), .A3(new_n539), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n716), .A2(new_n485), .A3(new_n488), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n650), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n674), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n597), .A2(new_n730), .A3(new_n698), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n733), .A2(new_n608), .A3(new_n486), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT45), .ZN(new_n735));
  INV_X1    g534(.A(new_n728), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT103), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(new_n533), .B2(new_n540), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n725), .A2(KEYINPUT103), .A3(new_n726), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n736), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n650), .A2(KEYINPUT44), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT44), .ZN(new_n743));
  OAI22_X1  g542(.A1(new_n740), .A2(new_n742), .B1(new_n743), .B2(new_n729), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n731), .ZN(new_n745));
  OAI21_X1  g544(.A(G29gat), .B1(new_n745), .B2(new_n536), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n735), .A2(new_n746), .ZN(G1328gat));
  AOI21_X1  g546(.A(G36gat), .B1(KEYINPUT104), .B2(KEYINPUT46), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n733), .A2(new_n487), .A3(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(G36gat), .B1(new_n745), .B2(new_n538), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(G1329gat));
  INV_X1    g552(.A(new_n650), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n714), .A2(G43gat), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n541), .A2(new_n754), .A3(new_n731), .A4(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT105), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n729), .A2(KEYINPUT105), .A3(new_n731), .A4(new_n755), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n738), .A2(new_n739), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n742), .B1(new_n761), .B2(new_n728), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n743), .B1(new_n541), .B2(new_n754), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n529), .B(new_n731), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n760), .B1(new_n764), .B2(G43gat), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT47), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n765), .A2(KEYINPUT106), .A3(new_n766), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n766), .A2(KEYINPUT106), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n766), .A2(KEYINPUT106), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n765), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n767), .A2(new_n770), .ZN(G1330gat));
  INV_X1    g570(.A(KEYINPUT48), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT107), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n723), .A2(G50gat), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n732), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n744), .A2(new_n464), .A3(new_n731), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n776), .B1(new_n777), .B2(G50gat), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n772), .A2(KEYINPUT107), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n778), .B(new_n779), .ZN(G1331gat));
  NAND2_X1  g579(.A1(new_n761), .A2(new_n728), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n651), .A2(new_n674), .A3(new_n699), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n486), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g585(.A1(new_n783), .A2(new_n538), .ZN(new_n787));
  NOR2_X1   g586(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n788));
  AND2_X1   g587(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n790), .B1(new_n787), .B2(new_n788), .ZN(G1333gat));
  XNOR2_X1  g590(.A(new_n537), .B(KEYINPUT108), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(G71gat), .B1(new_n784), .B2(new_n793), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n783), .A2(new_n564), .A3(new_n716), .ZN(new_n795));
  OR3_X1    g594(.A1(new_n794), .A2(new_n795), .A3(KEYINPUT50), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT50), .B1(new_n794), .B2(new_n795), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(G1334gat));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n723), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(new_n565), .ZN(G1335gat));
  NOR2_X1   g599(.A1(new_n597), .A2(new_n674), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n801), .A2(KEYINPUT109), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n801), .A2(KEYINPUT109), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n754), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT51), .B1(new_n781), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT51), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n740), .A2(new_n807), .A3(new_n804), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n809), .A2(new_n626), .A3(new_n486), .A4(new_n698), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n802), .A2(new_n803), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n811), .A2(new_n699), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n744), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(G85gat), .B1(new_n813), .B2(new_n536), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n810), .A2(new_n814), .ZN(G1336gat));
  OAI211_X1 g614(.A(new_n487), .B(new_n812), .C1(new_n762), .C2(new_n763), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT110), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n744), .A2(KEYINPUT110), .A3(new_n487), .A4(new_n812), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n818), .A2(G92gat), .A3(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n538), .A2(G92gat), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n698), .B(new_n822), .C1(new_n806), .C2(new_n808), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n820), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n816), .A2(G92gat), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT52), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n824), .A2(new_n827), .ZN(G1337gat));
  NOR3_X1   g627(.A1(new_n714), .A2(G99gat), .A3(new_n699), .ZN(new_n829));
  XOR2_X1   g628(.A(new_n829), .B(KEYINPUT111), .Z(new_n830));
  NAND2_X1  g629(.A1(new_n809), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(G99gat), .B1(new_n813), .B2(new_n716), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(G1338gat));
  NAND3_X1  g632(.A1(new_n744), .A2(new_n464), .A3(new_n812), .ZN(new_n834));
  XNOR2_X1  g633(.A(KEYINPUT112), .B(G106gat), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n723), .A2(G106gat), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n698), .B(new_n837), .C1(new_n806), .C2(new_n808), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(KEYINPUT53), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n836), .A2(new_n838), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(G1339gat));
  INV_X1    g642(.A(new_n597), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n845), .B(new_n685), .C1(new_n686), .C2(new_n688), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n846), .A2(new_n695), .ZN(new_n847));
  INV_X1    g646(.A(new_n688), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n677), .A2(new_n682), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n680), .B(new_n848), .C1(new_n849), .C2(KEYINPUT10), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(KEYINPUT54), .A3(new_n689), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n847), .A2(KEYINPUT55), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n697), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT55), .B1(new_n847), .B2(new_n851), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT113), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT55), .ZN(new_n856));
  INV_X1    g655(.A(new_n851), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n846), .A2(new_n695), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT113), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n859), .A2(new_n860), .A3(new_n697), .A4(new_n852), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n855), .A2(new_n674), .A3(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n662), .A2(new_n663), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n654), .B1(new_n653), .B2(new_n655), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n669), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n673), .A2(new_n865), .ZN(new_n866));
  AND3_X1   g665(.A1(new_n866), .A2(KEYINPUT114), .A3(new_n698), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT114), .B1(new_n866), .B2(new_n698), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n754), .B1(new_n862), .B2(new_n869), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n754), .A2(new_n866), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n855), .A2(new_n871), .A3(new_n861), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n844), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n652), .A2(new_n730), .A3(new_n699), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n877), .A2(new_n536), .ZN(new_n878));
  INV_X1    g677(.A(new_n532), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(new_n487), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n203), .A3(new_n674), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n486), .A2(new_n538), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n883), .A2(new_n714), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT115), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n885), .B1(new_n876), .B2(new_n723), .ZN(new_n886));
  AOI211_X1 g685(.A(KEYINPUT115), .B(new_n464), .C1(new_n874), .C2(new_n875), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n674), .B(new_n884), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT116), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n888), .A2(new_n889), .A3(G113gat), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n889), .B1(new_n888), .B2(G113gat), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n882), .B1(new_n890), .B2(new_n891), .ZN(G1340gat));
  NOR2_X1   g691(.A1(new_n699), .A2(G120gat), .ZN(new_n893));
  AND4_X1   g692(.A1(new_n486), .A2(new_n876), .A3(new_n880), .A4(new_n893), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n698), .B(new_n884), .C1(new_n886), .C2(new_n887), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n894), .B1(new_n895), .B2(G120gat), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT117), .ZN(G1341gat));
  NAND3_X1  g696(.A1(new_n881), .A2(new_n214), .A3(new_n597), .ZN(new_n898));
  OR2_X1    g697(.A1(new_n886), .A2(new_n887), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n899), .A2(new_n597), .A3(new_n884), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n898), .B1(new_n901), .B2(new_n214), .ZN(G1342gat));
  NAND3_X1  g701(.A1(new_n899), .A2(new_n754), .A3(new_n884), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(G134gat), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n878), .A2(new_n212), .A3(new_n754), .A4(new_n880), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT56), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n905), .A2(KEYINPUT56), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n904), .A2(new_n906), .A3(new_n907), .ZN(G1343gat));
  INV_X1    g707(.A(KEYINPUT120), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(KEYINPUT58), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n529), .A2(new_n883), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT57), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n723), .A2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n651), .A2(new_n674), .A3(new_n698), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT118), .B1(new_n857), .B2(new_n858), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n847), .A2(new_n918), .A3(new_n851), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n917), .A2(new_n856), .A3(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n853), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n920), .A2(new_n921), .A3(new_n674), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n866), .A2(new_n698), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n650), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n597), .B1(new_n925), .B2(new_n872), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n916), .B1(new_n926), .B2(KEYINPUT119), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n754), .B1(new_n922), .B2(new_n923), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n844), .B1(new_n928), .B2(new_n873), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT119), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n915), .B1(new_n927), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(KEYINPUT57), .B1(new_n876), .B2(new_n464), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n674), .B(new_n912), .C1(new_n932), .C2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n256), .A2(new_n257), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n529), .A2(new_n723), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(new_n538), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n730), .A2(G141gat), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n939), .A2(new_n876), .A3(new_n486), .A4(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT58), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(KEYINPUT120), .B2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n911), .B1(new_n936), .B2(new_n944), .ZN(new_n945));
  AOI211_X1 g744(.A(new_n910), .B(new_n943), .C1(new_n934), .C2(new_n935), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n945), .A2(new_n946), .ZN(G1344gat));
  INV_X1    g746(.A(KEYINPUT121), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n878), .A2(new_n939), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n698), .A2(new_n234), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n877), .A2(new_n536), .A3(new_n938), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n952), .A2(KEYINPUT121), .A3(new_n234), .A4(new_n698), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n853), .A2(new_n854), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n871), .A2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g755(.A(KEYINPUT122), .B1(new_n928), .B2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT122), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n730), .A2(new_n853), .ZN(new_n959));
  AOI22_X1  g758(.A1(new_n959), .A2(new_n920), .B1(new_n698), .B2(new_n866), .ZN(new_n960));
  OAI211_X1 g759(.A(new_n958), .B(new_n955), .C1(new_n960), .C2(new_n754), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n957), .A2(new_n961), .A3(new_n844), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n723), .B1(new_n962), .B2(new_n875), .ZN(new_n963));
  OAI22_X1  g762(.A1(new_n963), .A2(KEYINPUT57), .B1(new_n877), .B2(new_n915), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n964), .A2(new_n698), .A3(new_n912), .ZN(new_n965));
  AND2_X1   g764(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n966));
  AOI22_X1  g765(.A1(new_n951), .A2(new_n953), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(new_n912), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n876), .A2(new_n464), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(new_n913), .ZN(new_n970));
  INV_X1    g769(.A(new_n931), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n875), .B1(new_n929), .B2(new_n930), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n914), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n968), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n234), .B1(new_n974), .B2(new_n698), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n967), .B1(KEYINPUT59), .B2(new_n975), .ZN(G1345gat));
  AOI21_X1  g775(.A(new_n239), .B1(new_n974), .B2(new_n597), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n952), .A2(new_n239), .A3(new_n597), .ZN(new_n978));
  INV_X1    g777(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g778(.A(KEYINPUT123), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n912), .B1(new_n932), .B2(new_n933), .ZN(new_n981));
  OAI21_X1  g780(.A(G155gat), .B1(new_n981), .B2(new_n844), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT123), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n982), .A2(new_n983), .A3(new_n978), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n980), .A2(new_n984), .ZN(G1346gat));
  XNOR2_X1  g784(.A(KEYINPUT81), .B(G162gat), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n986), .B1(new_n952), .B2(new_n754), .ZN(new_n987));
  AND2_X1   g786(.A1(new_n754), .A2(new_n986), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n987), .B1(new_n974), .B2(new_n988), .ZN(G1347gat));
  NOR2_X1   g788(.A1(new_n879), .A2(new_n538), .ZN(new_n990));
  AND3_X1   g789(.A1(new_n876), .A2(new_n536), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g790(.A(G169gat), .B1(new_n991), .B2(new_n674), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n486), .A2(new_n538), .ZN(new_n993));
  INV_X1    g792(.A(new_n993), .ZN(new_n994));
  NOR2_X1   g793(.A1(new_n792), .A2(new_n994), .ZN(new_n995));
  AND2_X1   g794(.A1(new_n899), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g795(.A1(new_n730), .A2(new_n324), .ZN(new_n997));
  AOI21_X1  g796(.A(new_n992), .B1(new_n996), .B2(new_n997), .ZN(G1348gat));
  NAND3_X1  g797(.A1(new_n991), .A2(new_n325), .A3(new_n698), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n899), .A2(new_n698), .A3(new_n995), .ZN(new_n1000));
  INV_X1    g799(.A(new_n1000), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n999), .B1(new_n1001), .B2(new_n325), .ZN(G1349gat));
  INV_X1    g801(.A(KEYINPUT124), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(KEYINPUT60), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n876), .A2(new_n536), .A3(new_n990), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n597), .A2(new_n319), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n1004), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g806(.A(new_n597), .B(new_n995), .C1(new_n886), .C2(new_n887), .ZN(new_n1008));
  AOI21_X1  g807(.A(new_n1007), .B1(new_n1008), .B2(G183gat), .ZN(new_n1009));
  NOR2_X1   g808(.A1(new_n1003), .A2(KEYINPUT60), .ZN(new_n1010));
  XNOR2_X1  g809(.A(new_n1009), .B(new_n1010), .ZN(G1350gat));
  NAND3_X1  g810(.A1(new_n991), .A2(new_n315), .A3(new_n754), .ZN(new_n1012));
  OAI211_X1 g811(.A(new_n754), .B(new_n995), .C1(new_n886), .C2(new_n887), .ZN(new_n1013));
  INV_X1    g812(.A(KEYINPUT61), .ZN(new_n1014));
  AND3_X1   g813(.A1(new_n1013), .A2(new_n1014), .A3(G190gat), .ZN(new_n1015));
  AOI21_X1  g814(.A(new_n1014), .B1(new_n1013), .B2(G190gat), .ZN(new_n1016));
  OAI21_X1  g815(.A(new_n1012), .B1(new_n1015), .B2(new_n1016), .ZN(G1351gat));
  AND4_X1   g816(.A1(new_n536), .A2(new_n876), .A3(new_n487), .A4(new_n937), .ZN(new_n1018));
  AOI21_X1  g817(.A(G197gat), .B1(new_n1018), .B2(new_n674), .ZN(new_n1019));
  INV_X1    g818(.A(new_n964), .ZN(new_n1020));
  NOR2_X1   g819(.A1(new_n529), .A2(new_n994), .ZN(new_n1021));
  INV_X1    g820(.A(new_n1021), .ZN(new_n1022));
  NOR2_X1   g821(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  AND2_X1   g822(.A1(new_n674), .A2(G197gat), .ZN(new_n1024));
  AOI21_X1  g823(.A(new_n1019), .B1(new_n1023), .B2(new_n1024), .ZN(G1352gat));
  INV_X1    g824(.A(G204gat), .ZN(new_n1026));
  NAND3_X1  g825(.A1(new_n1018), .A2(new_n1026), .A3(new_n698), .ZN(new_n1027));
  INV_X1    g826(.A(KEYINPUT62), .ZN(new_n1028));
  NAND2_X1  g827(.A1(new_n1028), .A2(KEYINPUT125), .ZN(new_n1029));
  NAND2_X1  g828(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g829(.A(new_n1030), .B1(KEYINPUT125), .B2(new_n1028), .ZN(new_n1031));
  INV_X1    g830(.A(KEYINPUT125), .ZN(new_n1032));
  NAND3_X1  g831(.A1(new_n1027), .A2(new_n1032), .A3(KEYINPUT62), .ZN(new_n1033));
  NOR3_X1   g832(.A1(new_n1020), .A2(new_n699), .A3(new_n1022), .ZN(new_n1034));
  OAI211_X1 g833(.A(new_n1031), .B(new_n1033), .C1(new_n1026), .C2(new_n1034), .ZN(G1353gat));
  NAND4_X1  g834(.A1(new_n1018), .A2(new_n364), .A3(new_n366), .A4(new_n597), .ZN(new_n1036));
  NAND3_X1  g835(.A1(new_n964), .A2(new_n597), .A3(new_n1021), .ZN(new_n1037));
  AND2_X1   g836(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n1038));
  OAI21_X1  g837(.A(G211gat), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n1039));
  INV_X1    g838(.A(new_n1039), .ZN(new_n1040));
  AND3_X1   g839(.A1(new_n1037), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g840(.A(new_n1038), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1042));
  OAI21_X1  g841(.A(new_n1036), .B1(new_n1041), .B2(new_n1042), .ZN(G1354gat));
  AOI21_X1  g842(.A(G218gat), .B1(new_n1018), .B2(new_n754), .ZN(new_n1044));
  NAND2_X1  g843(.A1(new_n754), .A2(G218gat), .ZN(new_n1045));
  XNOR2_X1  g844(.A(new_n1045), .B(KEYINPUT127), .ZN(new_n1046));
  AOI21_X1  g845(.A(new_n1044), .B1(new_n1023), .B2(new_n1046), .ZN(G1355gat));
endmodule


