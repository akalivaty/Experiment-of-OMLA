

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779;

  AND2_X2 U376 ( .A1(n444), .A2(n383), .ZN(n361) );
  AND2_X2 U377 ( .A1(n628), .A2(n627), .ZN(n419) );
  AND2_X2 U378 ( .A1(n384), .A2(n564), .ZN(n632) );
  XNOR2_X2 U379 ( .A(n395), .B(KEYINPUT32), .ZN(n778) );
  NOR2_X2 U380 ( .A1(n394), .A2(n559), .ZN(n561) );
  XNOR2_X2 U381 ( .A(n546), .B(KEYINPUT4), .ZN(n510) );
  INV_X2 U382 ( .A(n762), .ZN(n444) );
  XNOR2_X1 U383 ( .A(n498), .B(n497), .ZN(n713) );
  NOR2_X2 U384 ( .A1(n664), .A2(n454), .ZN(n375) );
  NOR2_X1 U385 ( .A1(n673), .A2(n659), .ZN(n556) );
  INV_X1 U386 ( .A(n562), .ZN(n605) );
  NOR2_X1 U387 ( .A1(n568), .A2(n567), .ZN(n555) );
  INV_X1 U388 ( .A(n443), .ZN(n374) );
  INV_X2 U389 ( .A(G953), .ZN(n766) );
  NAND2_X1 U390 ( .A1(n393), .A2(n355), .ZN(n395) );
  AND2_X1 U391 ( .A1(n428), .A2(n426), .ZN(n425) );
  OR2_X1 U392 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U393 ( .A1(n356), .A2(n434), .ZN(n602) );
  XNOR2_X1 U394 ( .A(n601), .B(n367), .ZN(n422) );
  XNOR2_X1 U395 ( .A(n555), .B(KEYINPUT101), .ZN(n673) );
  AND2_X1 U396 ( .A1(n414), .A2(n413), .ZN(n412) );
  XNOR2_X1 U397 ( .A(n504), .B(n503), .ZN(n752) );
  XNOR2_X1 U398 ( .A(n392), .B(n391), .ZN(n503) );
  XNOR2_X1 U399 ( .A(n508), .B(n400), .ZN(n530) );
  XNOR2_X1 U400 ( .A(n536), .B(G475), .ZN(n537) );
  XNOR2_X1 U401 ( .A(G110), .B(G107), .ZN(n501) );
  XNOR2_X1 U402 ( .A(n472), .B(G125), .ZN(n508) );
  AND2_X1 U403 ( .A1(n422), .A2(n657), .ZN(n372) );
  XNOR2_X1 U404 ( .A(KEYINPUT82), .B(KEYINPUT39), .ZN(n637) );
  NAND2_X1 U405 ( .A1(n440), .A2(n363), .ZN(n439) );
  NOR2_X1 U406 ( .A1(n779), .A2(n773), .ZN(n639) );
  XNOR2_X1 U407 ( .A(G101), .B(KEYINPUT3), .ZN(n465) );
  XNOR2_X1 U408 ( .A(KEYINPUT10), .B(KEYINPUT67), .ZN(n400) );
  XNOR2_X1 U409 ( .A(n399), .B(n462), .ZN(n398) );
  XNOR2_X1 U410 ( .A(n528), .B(n527), .ZN(n399) );
  XNOR2_X1 U411 ( .A(KEYINPUT11), .B(KEYINPUT95), .ZN(n527) );
  XNOR2_X1 U412 ( .A(G113), .B(G131), .ZN(n532) );
  XOR2_X1 U413 ( .A(G140), .B(G143), .Z(n533) );
  XOR2_X1 U414 ( .A(G137), .B(G140), .Z(n492) );
  AND2_X1 U415 ( .A1(n427), .A2(n613), .ZN(n426) );
  NAND2_X1 U416 ( .A1(n454), .A2(KEYINPUT34), .ZN(n427) );
  NAND2_X1 U417 ( .A1(n424), .A2(KEYINPUT34), .ZN(n423) );
  NAND2_X1 U418 ( .A1(n415), .A2(G902), .ZN(n413) );
  XNOR2_X1 U419 ( .A(n498), .B(n469), .ZN(n650) );
  XNOR2_X1 U420 ( .A(n511), .B(n752), .ZN(n743) );
  INV_X1 U421 ( .A(n611), .ZN(n450) );
  INV_X1 U422 ( .A(KEYINPUT30), .ZN(n452) );
  XNOR2_X1 U423 ( .A(n385), .B(n600), .ZN(n384) );
  XNOR2_X1 U424 ( .A(n599), .B(KEYINPUT28), .ZN(n600) );
  NAND2_X1 U425 ( .A1(n387), .A2(n386), .ZN(n385) );
  XNOR2_X1 U426 ( .A(n485), .B(n460), .ZN(n486) );
  NAND2_X1 U427 ( .A1(n744), .A2(G478), .ZN(n459) );
  NAND2_X1 U428 ( .A1(n744), .A2(G475), .ZN(n449) );
  NAND2_X1 U429 ( .A1(n744), .A2(G210), .ZN(n433) );
  NAND2_X1 U430 ( .A1(n403), .A2(n550), .ZN(n402) );
  INV_X1 U431 ( .A(n500), .ZN(n403) );
  XOR2_X1 U432 ( .A(KEYINPUT12), .B(KEYINPUT94), .Z(n528) );
  NOR2_X1 U433 ( .A1(G953), .A2(G237), .ZN(n529) );
  XNOR2_X1 U434 ( .A(G134), .B(G131), .ZN(n463) );
  XNOR2_X1 U435 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n506) );
  NAND2_X1 U436 ( .A1(G234), .A2(G237), .ZN(n518) );
  NAND2_X1 U437 ( .A1(n516), .A2(n706), .ZN(n442) );
  OR2_X1 U438 ( .A1(n743), .A2(n441), .ZN(n440) );
  INV_X1 U439 ( .A(G237), .ZN(n513) );
  XNOR2_X1 U440 ( .A(G116), .B(G113), .ZN(n391) );
  XNOR2_X1 U441 ( .A(n465), .B(n464), .ZN(n392) );
  INV_X1 U442 ( .A(G119), .ZN(n464) );
  XOR2_X1 U443 ( .A(KEYINPUT98), .B(KEYINPUT7), .Z(n542) );
  XNOR2_X1 U444 ( .A(KEYINPUT97), .B(KEYINPUT9), .ZN(n541) );
  XNOR2_X1 U445 ( .A(G116), .B(G134), .ZN(n539) );
  XOR2_X1 U446 ( .A(G122), .B(G107), .Z(n540) );
  XNOR2_X1 U447 ( .A(n397), .B(n535), .ZN(n745) );
  XNOR2_X1 U448 ( .A(n534), .B(n354), .ZN(n535) );
  XNOR2_X1 U449 ( .A(n530), .B(n398), .ZN(n397) );
  XNOR2_X1 U450 ( .A(n429), .B(n554), .ZN(n587) );
  NAND2_X1 U451 ( .A1(n425), .A2(n423), .ZN(n429) );
  XNOR2_X1 U452 ( .A(n375), .B(KEYINPUT31), .ZN(n734) );
  NOR2_X1 U453 ( .A1(n374), .A2(KEYINPUT19), .ZN(n435) );
  OR2_X1 U454 ( .A1(n650), .A2(n411), .ZN(n410) );
  NAND2_X1 U455 ( .A1(n471), .A2(n550), .ZN(n411) );
  XNOR2_X1 U456 ( .A(G119), .B(G110), .ZN(n481) );
  XNOR2_X1 U457 ( .A(n638), .B(KEYINPUT40), .ZN(n779) );
  XNOR2_X1 U458 ( .A(n389), .B(n388), .ZN(n608) );
  INV_X1 U459 ( .A(KEYINPUT36), .ZN(n388) );
  INV_X1 U460 ( .A(G122), .ZN(n709) );
  BUF_X1 U461 ( .A(n587), .Z(n710) );
  AND2_X1 U462 ( .A1(n563), .A2(n605), .ZN(n717) );
  XNOR2_X1 U463 ( .A(n459), .B(n370), .ZN(n458) );
  INV_X1 U464 ( .A(KEYINPUT60), .ZN(n446) );
  XNOR2_X1 U465 ( .A(n449), .B(n368), .ZN(n448) );
  INV_X1 U466 ( .A(KEYINPUT56), .ZN(n430) );
  NAND2_X1 U467 ( .A1(n707), .A2(n706), .ZN(n711) );
  XOR2_X1 U468 ( .A(n533), .B(n532), .Z(n354) );
  AND2_X1 U469 ( .A1(n576), .A2(n396), .ZN(n355) );
  AND2_X1 U470 ( .A1(n438), .A2(n437), .ZN(n356) );
  INV_X1 U471 ( .A(n387), .ZN(n598) );
  AND2_X1 U472 ( .A1(n377), .A2(n376), .ZN(n357) );
  OR2_X1 U473 ( .A1(n644), .A2(n420), .ZN(n358) );
  OR2_X2 U474 ( .A1(n404), .A2(n401), .ZN(n601) );
  AND2_X1 U475 ( .A1(n657), .A2(n387), .ZN(n359) );
  AND2_X1 U476 ( .A1(n436), .A2(n443), .ZN(n360) );
  AND2_X1 U477 ( .A1(n565), .A2(n526), .ZN(n362) );
  AND2_X1 U478 ( .A1(n442), .A2(n675), .ZN(n363) );
  AND2_X1 U479 ( .A1(n440), .A2(n442), .ZN(n364) );
  AND2_X1 U480 ( .A1(n444), .A2(n648), .ZN(n365) );
  XOR2_X1 U481 ( .A(KEYINPUT100), .B(KEYINPUT6), .Z(n366) );
  XNOR2_X1 U482 ( .A(KEYINPUT65), .B(KEYINPUT1), .ZN(n367) );
  XNOR2_X1 U483 ( .A(n747), .B(n746), .ZN(n368) );
  XOR2_X1 U484 ( .A(n743), .B(n742), .Z(n369) );
  XNOR2_X1 U485 ( .A(n708), .B(KEYINPUT124), .ZN(n370) );
  INV_X1 U486 ( .A(KEYINPUT2), .ZN(n383) );
  AND2_X1 U487 ( .A1(n653), .A2(G953), .ZN(n751) );
  INV_X1 U488 ( .A(n751), .ZN(n457) );
  NAND2_X1 U489 ( .A1(n439), .A2(KEYINPUT19), .ZN(n438) );
  NAND2_X1 U490 ( .A1(n448), .A2(n457), .ZN(n447) );
  XNOR2_X2 U491 ( .A(n371), .B(KEYINPUT33), .ZN(n669) );
  NAND2_X1 U492 ( .A1(n372), .A2(n606), .ZN(n371) );
  NOR2_X1 U493 ( .A1(G902), .A2(n748), .ZN(n487) );
  NOR2_X1 U494 ( .A1(n605), .A2(n461), .ZN(n386) );
  NAND2_X1 U495 ( .A1(n713), .A2(n500), .ZN(n406) );
  NAND2_X1 U496 ( .A1(n406), .A2(n405), .ZN(n404) );
  NAND2_X1 U497 ( .A1(n373), .A2(KEYINPUT47), .ZN(n618) );
  NAND2_X1 U498 ( .A1(n604), .A2(n672), .ZN(n373) );
  XNOR2_X2 U499 ( .A(n387), .B(n366), .ZN(n606) );
  NOR2_X1 U500 ( .A1(n607), .A2(n735), .ZN(n390) );
  NAND2_X1 U501 ( .A1(n643), .A2(n360), .ZN(n389) );
  NAND2_X1 U502 ( .A1(n374), .A2(KEYINPUT19), .ZN(n437) );
  NAND2_X4 U503 ( .A1(n412), .A2(n410), .ZN(n387) );
  INV_X1 U504 ( .A(n636), .ZN(n376) );
  NOR2_X1 U505 ( .A1(n635), .A2(n670), .ZN(n377) );
  XNOR2_X1 U506 ( .A(n453), .B(n452), .ZN(n451) );
  NAND2_X1 U507 ( .A1(n381), .A2(n692), .ZN(n707) );
  AND2_X1 U508 ( .A1(n445), .A2(n444), .ZN(n689) );
  NAND2_X1 U509 ( .A1(n365), .A2(n445), .ZN(n692) );
  NAND2_X1 U510 ( .A1(n378), .A2(KEYINPUT2), .ZN(n380) );
  NAND2_X1 U511 ( .A1(n445), .A2(n444), .ZN(n378) );
  NAND2_X1 U512 ( .A1(n380), .A2(n379), .ZN(n382) );
  NAND2_X1 U513 ( .A1(n361), .A2(n445), .ZN(n379) );
  NAND2_X1 U514 ( .A1(n382), .A2(n690), .ZN(n381) );
  NAND2_X1 U515 ( .A1(n387), .A2(n675), .ZN(n453) );
  NOR2_X1 U516 ( .A1(n610), .A2(n387), .ZN(n566) );
  NOR2_X1 U517 ( .A1(n661), .A2(n387), .ZN(n662) );
  AND2_X1 U518 ( .A1(n606), .A2(n390), .ZN(n643) );
  INV_X1 U519 ( .A(n394), .ZN(n393) );
  NOR2_X1 U520 ( .A1(n394), .A2(n578), .ZN(n579) );
  XNOR2_X2 U521 ( .A(n558), .B(KEYINPUT22), .ZN(n394) );
  XNOR2_X1 U522 ( .A(n575), .B(KEYINPUT103), .ZN(n396) );
  NOR2_X1 U523 ( .A1(n713), .A2(n402), .ZN(n401) );
  NAND2_X1 U524 ( .A1(n500), .A2(G902), .ZN(n405) );
  XNOR2_X1 U525 ( .A(n407), .B(KEYINPUT85), .ZN(n582) );
  NAND2_X1 U526 ( .A1(n573), .A2(n574), .ZN(n407) );
  NAND2_X1 U527 ( .A1(n436), .A2(n435), .ZN(n434) );
  INV_X2 U528 ( .A(G146), .ZN(n472) );
  NOR2_X2 U529 ( .A1(G902), .A2(n745), .ZN(n538) );
  OR2_X2 U530 ( .A1(n732), .A2(n408), .ZN(n604) );
  INV_X1 U531 ( .A(KEYINPUT78), .ZN(n408) );
  XNOR2_X2 U532 ( .A(n603), .B(n409), .ZN(n732) );
  INV_X1 U533 ( .A(KEYINPUT74), .ZN(n409) );
  NAND2_X1 U534 ( .A1(n650), .A2(n415), .ZN(n414) );
  INV_X1 U535 ( .A(n471), .ZN(n415) );
  NAND2_X1 U536 ( .A1(n416), .A2(n647), .ZN(n762) );
  XNOR2_X1 U537 ( .A(n418), .B(n417), .ZN(n416) );
  INV_X1 U538 ( .A(KEYINPUT48), .ZN(n417) );
  NAND2_X1 U539 ( .A1(n419), .A2(n640), .ZN(n418) );
  BUF_X2 U540 ( .A(n422), .Z(n420) );
  INV_X1 U541 ( .A(n420), .ZN(n577) );
  NAND2_X1 U542 ( .A1(n562), .A2(n420), .ZN(n575) );
  NAND2_X1 U543 ( .A1(n421), .A2(n577), .ZN(n559) );
  INV_X1 U544 ( .A(n606), .ZN(n421) );
  NOR2_X1 U545 ( .A1(n657), .A2(n420), .ZN(n658) );
  NAND2_X1 U546 ( .A1(n359), .A2(n420), .ZN(n664) );
  NAND2_X1 U547 ( .A1(n608), .A2(n420), .ZN(n609) );
  INV_X1 U548 ( .A(n669), .ZN(n424) );
  NAND2_X1 U549 ( .A1(n669), .A2(n362), .ZN(n428) );
  XNOR2_X1 U550 ( .A(n431), .B(n430), .ZN(G51) );
  NAND2_X1 U551 ( .A1(n432), .A2(n457), .ZN(n431) );
  XNOR2_X1 U552 ( .A(n433), .B(n369), .ZN(n432) );
  INV_X1 U553 ( .A(n439), .ZN(n436) );
  NAND2_X1 U554 ( .A1(n443), .A2(n364), .ZN(n645) );
  OR2_X1 U555 ( .A1(n516), .A2(n706), .ZN(n441) );
  NAND2_X1 U556 ( .A1(n743), .A2(n516), .ZN(n443) );
  XNOR2_X2 U557 ( .A(n592), .B(KEYINPUT45), .ZN(n445) );
  AND2_X1 U558 ( .A1(n445), .A2(n766), .ZN(n755) );
  XNOR2_X1 U559 ( .A(n447), .B(n446), .ZN(G60) );
  NAND2_X1 U560 ( .A1(n451), .A2(n450), .ZN(n635) );
  INV_X1 U561 ( .A(n565), .ZN(n454) );
  XNOR2_X2 U562 ( .A(n525), .B(n524), .ZN(n565) );
  XNOR2_X2 U563 ( .A(n455), .B(G143), .ZN(n546) );
  XNOR2_X2 U564 ( .A(G128), .B(KEYINPUT75), .ZN(n455) );
  NOR2_X2 U565 ( .A1(n562), .A2(n659), .ZN(n657) );
  XNOR2_X1 U566 ( .A(n456), .B(KEYINPUT125), .ZN(G63) );
  NAND2_X1 U567 ( .A1(n458), .A2(n457), .ZN(n456) );
  NOR2_X1 U568 ( .A1(n654), .A2(n751), .ZN(n656) );
  XNOR2_X1 U569 ( .A(n357), .B(n637), .ZN(n642) );
  NOR2_X1 U570 ( .A1(n711), .A2(n649), .ZN(n652) );
  XNOR2_X1 U571 ( .A(KEYINPUT72), .B(n484), .ZN(n460) );
  OR2_X1 U572 ( .A1(n611), .A2(n659), .ZN(n461) );
  AND2_X1 U573 ( .A1(G214), .A2(n529), .ZN(n462) );
  NOR2_X1 U574 ( .A1(n717), .A2(n572), .ZN(n573) );
  INV_X1 U575 ( .A(KEYINPUT84), .ZN(n583) );
  INV_X1 U576 ( .A(KEYINPUT108), .ZN(n599) );
  INV_X1 U577 ( .A(n492), .ZN(n477) );
  XNOR2_X1 U578 ( .A(n470), .B(G472), .ZN(n471) );
  INV_X1 U579 ( .A(KEYINPUT63), .ZN(n655) );
  XNOR2_X1 U580 ( .A(n704), .B(n703), .ZN(G75) );
  XNOR2_X2 U581 ( .A(n510), .B(n463), .ZN(n765) );
  XNOR2_X2 U582 ( .A(n765), .B(n472), .ZN(n498) );
  XOR2_X1 U583 ( .A(G137), .B(KEYINPUT5), .Z(n467) );
  NAND2_X1 U584 ( .A1(n529), .A2(G210), .ZN(n466) );
  XNOR2_X1 U585 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U586 ( .A(n503), .B(n468), .ZN(n469) );
  XNOR2_X1 U587 ( .A(KEYINPUT69), .B(KEYINPUT92), .ZN(n470) );
  XOR2_X1 U588 ( .A(KEYINPUT80), .B(KEYINPUT23), .Z(n474) );
  XNOR2_X1 U589 ( .A(G128), .B(KEYINPUT24), .ZN(n473) );
  XNOR2_X1 U590 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U591 ( .A(n530), .B(n475), .Z(n480) );
  NAND2_X1 U592 ( .A1(G234), .A2(n766), .ZN(n476) );
  XOR2_X1 U593 ( .A(KEYINPUT8), .B(n476), .Z(n545) );
  NAND2_X1 U594 ( .A1(G221), .A2(n545), .ZN(n478) );
  XNOR2_X1 U595 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U596 ( .A(n480), .B(n479), .ZN(n482) );
  XNOR2_X1 U597 ( .A(n482), .B(n481), .ZN(n748) );
  XNOR2_X1 U598 ( .A(KEYINPUT15), .B(G902), .ZN(n512) );
  NAND2_X1 U599 ( .A1(G234), .A2(n512), .ZN(n483) );
  XNOR2_X1 U600 ( .A(KEYINPUT20), .B(n483), .ZN(n488) );
  NAND2_X1 U601 ( .A1(n488), .A2(G217), .ZN(n485) );
  XOR2_X1 U602 ( .A(KEYINPUT90), .B(KEYINPUT25), .Z(n484) );
  XNOR2_X2 U603 ( .A(n487), .B(n486), .ZN(n562) );
  NAND2_X1 U604 ( .A1(G221), .A2(n488), .ZN(n489) );
  XNOR2_X1 U605 ( .A(n489), .B(KEYINPUT91), .ZN(n491) );
  INV_X1 U606 ( .A(KEYINPUT21), .ZN(n490) );
  XNOR2_X1 U607 ( .A(n491), .B(n490), .ZN(n659) );
  XOR2_X1 U608 ( .A(KEYINPUT89), .B(n492), .Z(n763) );
  NAND2_X1 U609 ( .A1(G227), .A2(n766), .ZN(n493) );
  XNOR2_X1 U610 ( .A(G104), .B(n493), .ZN(n494) );
  XNOR2_X1 U611 ( .A(n494), .B(G101), .ZN(n495) );
  XNOR2_X1 U612 ( .A(n501), .B(n495), .ZN(n496) );
  XNOR2_X1 U613 ( .A(n763), .B(n496), .ZN(n497) );
  INV_X1 U614 ( .A(KEYINPUT68), .ZN(n499) );
  XNOR2_X1 U615 ( .A(n499), .B(G469), .ZN(n500) );
  XNOR2_X1 U616 ( .A(n501), .B(KEYINPUT16), .ZN(n502) );
  XNOR2_X1 U617 ( .A(n709), .B(G104), .ZN(n531) );
  XNOR2_X1 U618 ( .A(n502), .B(n531), .ZN(n504) );
  NAND2_X1 U619 ( .A1(n766), .A2(G224), .ZN(n505) );
  XNOR2_X1 U620 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U621 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U622 ( .A(n510), .B(n509), .ZN(n511) );
  INV_X1 U623 ( .A(n512), .ZN(n706) );
  INV_X1 U624 ( .A(G902), .ZN(n550) );
  NAND2_X1 U625 ( .A1(n550), .A2(n513), .ZN(n517) );
  NAND2_X1 U626 ( .A1(n517), .A2(G210), .ZN(n515) );
  INV_X1 U627 ( .A(KEYINPUT87), .ZN(n514) );
  XNOR2_X1 U628 ( .A(n515), .B(n514), .ZN(n516) );
  NAND2_X1 U629 ( .A1(n517), .A2(G214), .ZN(n675) );
  XNOR2_X1 U630 ( .A(n518), .B(KEYINPUT14), .ZN(n520) );
  NAND2_X1 U631 ( .A1(G952), .A2(n520), .ZN(n519) );
  XNOR2_X1 U632 ( .A(KEYINPUT88), .B(n519), .ZN(n684) );
  NOR2_X1 U633 ( .A1(n684), .A2(G953), .ZN(n597) );
  NOR2_X1 U634 ( .A1(G898), .A2(n766), .ZN(n753) );
  INV_X1 U635 ( .A(n753), .ZN(n521) );
  NAND2_X1 U636 ( .A1(G902), .A2(n520), .ZN(n593) );
  NOR2_X1 U637 ( .A1(n521), .A2(n593), .ZN(n522) );
  OR2_X1 U638 ( .A1(n597), .A2(n522), .ZN(n523) );
  NAND2_X1 U639 ( .A1(n602), .A2(n523), .ZN(n525) );
  INV_X1 U640 ( .A(KEYINPUT0), .ZN(n524) );
  INV_X1 U641 ( .A(KEYINPUT34), .ZN(n526) );
  XNOR2_X1 U642 ( .A(n531), .B(KEYINPUT93), .ZN(n534) );
  XNOR2_X1 U643 ( .A(KEYINPUT96), .B(KEYINPUT13), .ZN(n536) );
  XNOR2_X2 U644 ( .A(n538), .B(n537), .ZN(n568) );
  XNOR2_X1 U645 ( .A(n540), .B(n539), .ZN(n544) );
  XNOR2_X1 U646 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U647 ( .A(n544), .B(n543), .Z(n549) );
  NAND2_X1 U648 ( .A1(G217), .A2(n545), .ZN(n547) );
  XNOR2_X1 U649 ( .A(n546), .B(n547), .ZN(n548) );
  XNOR2_X1 U650 ( .A(n549), .B(n548), .ZN(n708) );
  NAND2_X1 U651 ( .A1(n708), .A2(n550), .ZN(n551) );
  XNOR2_X1 U652 ( .A(n551), .B(G478), .ZN(n567) );
  AND2_X1 U653 ( .A1(n568), .A2(n567), .ZN(n552) );
  XNOR2_X1 U654 ( .A(n552), .B(KEYINPUT104), .ZN(n613) );
  INV_X1 U655 ( .A(KEYINPUT81), .ZN(n553) );
  XNOR2_X1 U656 ( .A(n553), .B(KEYINPUT35), .ZN(n554) );
  NAND2_X1 U657 ( .A1(n587), .A2(KEYINPUT44), .ZN(n574) );
  XNOR2_X1 U658 ( .A(n556), .B(KEYINPUT102), .ZN(n557) );
  NAND2_X1 U659 ( .A1(n557), .A2(n565), .ZN(n558) );
  INV_X1 U660 ( .A(KEYINPUT83), .ZN(n560) );
  XNOR2_X1 U661 ( .A(n561), .B(n560), .ZN(n563) );
  INV_X1 U662 ( .A(n601), .ZN(n564) );
  NAND2_X1 U663 ( .A1(n657), .A2(n564), .ZN(n610) );
  NAND2_X1 U664 ( .A1(n566), .A2(n565), .ZN(n720) );
  NAND2_X1 U665 ( .A1(n734), .A2(n720), .ZN(n571) );
  INV_X1 U666 ( .A(n567), .ZN(n569) );
  NOR2_X1 U667 ( .A1(n569), .A2(n568), .ZN(n728) );
  INV_X1 U668 ( .A(n728), .ZN(n737) );
  XOR2_X1 U669 ( .A(KEYINPUT99), .B(n737), .Z(n641) );
  NAND2_X1 U670 ( .A1(n569), .A2(n568), .ZN(n735) );
  NAND2_X1 U671 ( .A1(n641), .A2(n735), .ZN(n672) );
  INV_X1 U672 ( .A(KEYINPUT79), .ZN(n570) );
  XNOR2_X1 U673 ( .A(n672), .B(n570), .ZN(n619) );
  AND2_X1 U674 ( .A1(n571), .A2(n619), .ZN(n572) );
  XNOR2_X1 U675 ( .A(n606), .B(KEYINPUT73), .ZN(n576) );
  NAND2_X1 U676 ( .A1(n598), .A2(n577), .ZN(n578) );
  NAND2_X1 U677 ( .A1(n562), .A2(n579), .ZN(n727) );
  NAND2_X1 U678 ( .A1(n778), .A2(n727), .ZN(n585) );
  NAND2_X1 U679 ( .A1(n585), .A2(KEYINPUT44), .ZN(n580) );
  XNOR2_X1 U680 ( .A(n580), .B(KEYINPUT64), .ZN(n581) );
  NAND2_X1 U681 ( .A1(n582), .A2(n581), .ZN(n584) );
  XNOR2_X1 U682 ( .A(n584), .B(n583), .ZN(n591) );
  XNOR2_X1 U683 ( .A(KEYINPUT86), .B(n585), .ZN(n586) );
  NOR2_X1 U684 ( .A1(n586), .A2(KEYINPUT44), .ZN(n589) );
  INV_X1 U685 ( .A(n710), .ZN(n588) );
  NAND2_X1 U686 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U687 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U688 ( .A1(G900), .A2(n593), .ZN(n594) );
  NAND2_X1 U689 ( .A1(G953), .A2(n594), .ZN(n595) );
  XNOR2_X1 U690 ( .A(KEYINPUT105), .B(n595), .ZN(n596) );
  NOR2_X1 U691 ( .A1(n597), .A2(n596), .ZN(n611) );
  NAND2_X1 U692 ( .A1(n632), .A2(n602), .ZN(n603) );
  OR2_X1 U693 ( .A1(n605), .A2(n461), .ZN(n607) );
  INV_X1 U694 ( .A(n735), .ZN(n731) );
  XNOR2_X1 U695 ( .A(n609), .B(KEYINPUT111), .ZN(n775) );
  XNOR2_X1 U696 ( .A(n610), .B(KEYINPUT106), .ZN(n636) );
  OR2_X1 U697 ( .A1(n636), .A2(n635), .ZN(n615) );
  INV_X1 U698 ( .A(n645), .ZN(n612) );
  NAND2_X1 U699 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U700 ( .A(KEYINPUT107), .B(n616), .ZN(n774) );
  NOR2_X1 U701 ( .A1(n775), .A2(n774), .ZN(n617) );
  AND2_X1 U702 ( .A1(n618), .A2(n617), .ZN(n628) );
  INV_X1 U703 ( .A(KEYINPUT70), .ZN(n622) );
  INV_X1 U704 ( .A(KEYINPUT47), .ZN(n623) );
  AND2_X1 U705 ( .A1(n623), .A2(n619), .ZN(n620) );
  NAND2_X1 U706 ( .A1(n732), .A2(n620), .ZN(n621) );
  XNOR2_X1 U707 ( .A(n622), .B(n621), .ZN(n626) );
  NOR2_X1 U708 ( .A1(n732), .A2(n623), .ZN(n624) );
  NOR2_X1 U709 ( .A1(KEYINPUT78), .A2(n624), .ZN(n625) );
  NOR2_X1 U710 ( .A1(n626), .A2(n625), .ZN(n627) );
  XOR2_X1 U711 ( .A(KEYINPUT109), .B(KEYINPUT41), .Z(n631) );
  INV_X1 U712 ( .A(KEYINPUT38), .ZN(n629) );
  XNOR2_X1 U713 ( .A(n645), .B(n629), .ZN(n670) );
  NOR2_X1 U714 ( .A1(n673), .A2(n670), .ZN(n677) );
  NAND2_X1 U715 ( .A1(n677), .A2(n675), .ZN(n630) );
  XNOR2_X1 U716 ( .A(n631), .B(n630), .ZN(n697) );
  NAND2_X1 U717 ( .A1(n697), .A2(n632), .ZN(n634) );
  XOR2_X1 U718 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n633) );
  XNOR2_X1 U719 ( .A(n634), .B(n633), .ZN(n773) );
  NOR2_X1 U720 ( .A1(n642), .A2(n735), .ZN(n638) );
  XNOR2_X1 U721 ( .A(n639), .B(KEYINPUT46), .ZN(n640) );
  NOR2_X1 U722 ( .A1(n642), .A2(n641), .ZN(n739) );
  NAND2_X1 U723 ( .A1(n643), .A2(n675), .ZN(n644) );
  XNOR2_X1 U724 ( .A(n358), .B(KEYINPUT43), .ZN(n646) );
  AND2_X1 U725 ( .A1(n646), .A2(n645), .ZN(n705) );
  NOR2_X1 U726 ( .A1(n739), .A2(n705), .ZN(n647) );
  INV_X1 U727 ( .A(KEYINPUT71), .ZN(n690) );
  AND2_X1 U728 ( .A1(KEYINPUT2), .A2(KEYINPUT71), .ZN(n648) );
  INV_X1 U729 ( .A(G472), .ZN(n649) );
  XOR2_X1 U730 ( .A(KEYINPUT62), .B(n650), .Z(n651) );
  XNOR2_X1 U731 ( .A(n652), .B(n651), .ZN(n654) );
  INV_X1 U732 ( .A(G952), .ZN(n653) );
  XNOR2_X1 U733 ( .A(n656), .B(n655), .ZN(G57) );
  XOR2_X1 U734 ( .A(KEYINPUT50), .B(n658), .Z(n663) );
  AND2_X1 U735 ( .A1(n659), .A2(n562), .ZN(n660) );
  XOR2_X1 U736 ( .A(KEYINPUT49), .B(n660), .Z(n661) );
  NAND2_X1 U737 ( .A1(n663), .A2(n662), .ZN(n665) );
  NAND2_X1 U738 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U739 ( .A(KEYINPUT51), .B(n666), .Z(n667) );
  NAND2_X1 U740 ( .A1(n697), .A2(n667), .ZN(n668) );
  XOR2_X1 U741 ( .A(KEYINPUT118), .B(n668), .Z(n681) );
  INV_X1 U742 ( .A(n670), .ZN(n671) );
  NAND2_X1 U743 ( .A1(n672), .A2(n671), .ZN(n674) );
  NAND2_X1 U744 ( .A1(n674), .A2(n673), .ZN(n676) );
  AND2_X1 U745 ( .A1(n676), .A2(n675), .ZN(n678) );
  NOR2_X1 U746 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U747 ( .A1(n424), .A2(n679), .ZN(n680) );
  NOR2_X1 U748 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U749 ( .A(n682), .B(KEYINPUT52), .ZN(n683) );
  NOR2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U751 ( .A(KEYINPUT119), .B(n685), .ZN(n702) );
  INV_X1 U752 ( .A(n689), .ZN(n687) );
  XOR2_X1 U753 ( .A(KEYINPUT77), .B(n383), .Z(n686) );
  NAND2_X1 U754 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U755 ( .A(n688), .B(KEYINPUT76), .ZN(n695) );
  NAND2_X1 U756 ( .A1(n689), .A2(KEYINPUT2), .ZN(n691) );
  NAND2_X1 U757 ( .A1(n691), .A2(n690), .ZN(n693) );
  NAND2_X1 U758 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U759 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U760 ( .A1(n696), .A2(n766), .ZN(n700) );
  NAND2_X1 U761 ( .A1(n697), .A2(n669), .ZN(n698) );
  XOR2_X1 U762 ( .A(n698), .B(KEYINPUT120), .Z(n699) );
  NOR2_X1 U763 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U764 ( .A1(n702), .A2(n701), .ZN(n704) );
  XNOR2_X1 U765 ( .A(KEYINPUT53), .B(KEYINPUT121), .ZN(n703) );
  XOR2_X1 U766 ( .A(n705), .B(G140), .Z(G42) );
  AND2_X2 U767 ( .A1(n707), .A2(n706), .ZN(n744) );
  XNOR2_X1 U768 ( .A(n710), .B(n709), .ZN(G24) );
  NAND2_X1 U769 ( .A1(n744), .A2(G469), .ZN(n715) );
  XOR2_X1 U770 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n712) );
  XNOR2_X1 U771 ( .A(n713), .B(n712), .ZN(n714) );
  XNOR2_X1 U772 ( .A(n715), .B(n714), .ZN(n716) );
  NOR2_X1 U773 ( .A1(n716), .A2(n751), .ZN(G54) );
  XOR2_X1 U774 ( .A(n717), .B(G101), .Z(n718) );
  XNOR2_X1 U775 ( .A(KEYINPUT112), .B(n718), .ZN(G3) );
  NOR2_X1 U776 ( .A1(n735), .A2(n720), .ZN(n719) );
  XOR2_X1 U777 ( .A(G104), .B(n719), .Z(G6) );
  NOR2_X1 U778 ( .A1(n737), .A2(n720), .ZN(n725) );
  XOR2_X1 U779 ( .A(KEYINPUT27), .B(KEYINPUT114), .Z(n722) );
  XNOR2_X1 U780 ( .A(G107), .B(KEYINPUT26), .ZN(n721) );
  XNOR2_X1 U781 ( .A(n722), .B(n721), .ZN(n723) );
  XNOR2_X1 U782 ( .A(KEYINPUT113), .B(n723), .ZN(n724) );
  XNOR2_X1 U783 ( .A(n725), .B(n724), .ZN(G9) );
  XOR2_X1 U784 ( .A(G110), .B(KEYINPUT115), .Z(n726) );
  XNOR2_X1 U785 ( .A(n727), .B(n726), .ZN(G12) );
  XOR2_X1 U786 ( .A(G128), .B(KEYINPUT29), .Z(n730) );
  NAND2_X1 U787 ( .A1(n728), .A2(n732), .ZN(n729) );
  XNOR2_X1 U788 ( .A(n730), .B(n729), .ZN(G30) );
  NAND2_X1 U789 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U790 ( .A(n733), .B(G146), .ZN(G48) );
  NOR2_X1 U791 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U792 ( .A(G113), .B(n736), .Z(G15) );
  NOR2_X1 U793 ( .A1(n737), .A2(n734), .ZN(n738) );
  XOR2_X1 U794 ( .A(G116), .B(n738), .Z(G18) );
  XNOR2_X1 U795 ( .A(G134), .B(n739), .ZN(n740) );
  XNOR2_X1 U796 ( .A(n740), .B(KEYINPUT117), .ZN(G36) );
  XOR2_X1 U797 ( .A(KEYINPUT55), .B(KEYINPUT54), .Z(n741) );
  XNOR2_X1 U798 ( .A(n741), .B(KEYINPUT122), .ZN(n742) );
  XOR2_X1 U799 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n747) );
  XNOR2_X1 U800 ( .A(n745), .B(KEYINPUT66), .ZN(n746) );
  NAND2_X1 U801 ( .A1(n744), .A2(G217), .ZN(n749) );
  XNOR2_X1 U802 ( .A(n749), .B(n748), .ZN(n750) );
  NOR2_X1 U803 ( .A1(n751), .A2(n750), .ZN(G66) );
  XOR2_X1 U804 ( .A(KEYINPUT127), .B(n752), .Z(n754) );
  NOR2_X1 U805 ( .A1(n754), .A2(n753), .ZN(n761) );
  XOR2_X1 U806 ( .A(KEYINPUT126), .B(n755), .Z(n759) );
  NAND2_X1 U807 ( .A1(G953), .A2(G224), .ZN(n756) );
  XNOR2_X1 U808 ( .A(KEYINPUT61), .B(n756), .ZN(n757) );
  NAND2_X1 U809 ( .A1(n757), .A2(G898), .ZN(n758) );
  NAND2_X1 U810 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U811 ( .A(n761), .B(n760), .ZN(G69) );
  XNOR2_X1 U812 ( .A(n530), .B(n763), .ZN(n764) );
  XOR2_X1 U813 ( .A(n765), .B(n764), .Z(n768) );
  XNOR2_X1 U814 ( .A(n762), .B(n768), .ZN(n767) );
  NAND2_X1 U815 ( .A1(n767), .A2(n766), .ZN(n772) );
  XNOR2_X1 U816 ( .A(n768), .B(G227), .ZN(n769) );
  NAND2_X1 U817 ( .A1(n769), .A2(G900), .ZN(n770) );
  NAND2_X1 U818 ( .A1(n770), .A2(G953), .ZN(n771) );
  NAND2_X1 U819 ( .A1(n772), .A2(n771), .ZN(G72) );
  XOR2_X1 U820 ( .A(G137), .B(n773), .Z(G39) );
  XOR2_X1 U821 ( .A(G143), .B(n774), .Z(G45) );
  XNOR2_X1 U822 ( .A(n775), .B(KEYINPUT37), .ZN(n776) );
  XNOR2_X1 U823 ( .A(n776), .B(KEYINPUT116), .ZN(n777) );
  XNOR2_X1 U824 ( .A(G125), .B(n777), .ZN(G27) );
  XNOR2_X1 U825 ( .A(G119), .B(n778), .ZN(G21) );
  XOR2_X1 U826 ( .A(G131), .B(n779), .Z(G33) );
endmodule

