//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 0 1 0 1 1 1 0 0 0 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1243, new_n1244, new_n1245, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1306, new_n1307, new_n1308, new_n1309;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G107), .A2(G264), .ZN(new_n208));
  INV_X1    g0008(.A(G97), .ZN(new_n209));
  INV_X1    g0009(.A(G257), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n207), .B(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  OR2_X1    g0011(.A1(new_n211), .A2(KEYINPUT65), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(KEYINPUT65), .ZN(new_n213));
  INV_X1    g0013(.A(G226), .ZN(new_n214));
  INV_X1    g0014(.A(G116), .ZN(new_n215));
  INV_X1    g0015(.A(G270), .ZN(new_n216));
  OAI22_X1  g0016(.A1(new_n202), .A2(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT64), .B(G77), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n217), .B1(G244), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n212), .A2(new_n213), .A3(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n206), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT1), .Z(new_n225));
  NOR2_X1   g0025(.A1(new_n206), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT0), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G20), .ZN(new_n231));
  OAI21_X1  g0031(.A(G50), .B1(G58), .B2(G68), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n225), .B(new_n228), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT2), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n214), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G264), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n216), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G58), .ZN(new_n245));
  INV_X1    g0045(.A(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(G107), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(new_n215), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(new_n218), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT3), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT3), .B(G33), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G222), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G223), .A2(G1698), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n260), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  AND3_X1   g0064(.A1(new_n258), .A2(new_n259), .A3(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G41), .A2(G45), .ZN(new_n266));
  INV_X1    g0066(.A(G274), .ZN(new_n267));
  NOR3_X1   g0067(.A1(new_n266), .A2(G1), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G41), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n230), .B1(new_n255), .B2(new_n270), .ZN(new_n271));
  AND2_X1   g0071(.A1(KEYINPUT66), .A2(G1), .ZN(new_n272));
  NOR2_X1   g0072(.A1(KEYINPUT66), .A2(G1), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n271), .B1(new_n274), .B2(new_n266), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n269), .B1(new_n275), .B2(new_n214), .ZN(new_n276));
  OAI21_X1  g0076(.A(G200), .B1(new_n265), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n203), .A2(G20), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G20), .A2(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G150), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT8), .B(G58), .ZN(new_n281));
  INV_X1    g0081(.A(G20), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G33), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n278), .B(new_n280), .C1(new_n281), .C2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n229), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  OR2_X1    g0087(.A1(KEYINPUT66), .A2(G1), .ZN(new_n288));
  NAND2_X1  g0088(.A1(KEYINPUT66), .A2(G1), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n286), .B1(new_n290), .B2(G20), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G50), .ZN(new_n292));
  OAI211_X1 g0092(.A(G13), .B(G20), .C1(new_n272), .C2(new_n273), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n202), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n287), .A2(new_n292), .A3(KEYINPUT9), .A4(new_n295), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n277), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT10), .ZN(new_n298));
  INV_X1    g0098(.A(new_n266), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n259), .B1(new_n290), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n268), .B1(new_n300), .B2(G226), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n258), .A2(new_n259), .A3(new_n264), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n301), .A2(G190), .A3(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n287), .A2(new_n295), .A3(new_n292), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT9), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n297), .A2(new_n298), .A3(new_n303), .A4(new_n306), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n306), .A2(new_n303), .A3(new_n277), .A4(new_n296), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT10), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT11), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n221), .A2(G20), .ZN(new_n312));
  INV_X1    g0112(.A(new_n279), .ZN(new_n313));
  OAI221_X1 g0113(.A(new_n312), .B1(new_n283), .B2(new_n246), .C1(new_n313), .C2(new_n202), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT69), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n314), .A2(new_n315), .A3(new_n286), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n315), .B1(new_n314), .B2(new_n286), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n311), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n318), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n320), .A2(KEYINPUT11), .A3(new_n316), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n294), .A2(new_n221), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n322), .B(KEYINPUT12), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n291), .A2(G68), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n319), .A2(new_n321), .A3(new_n323), .A4(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n214), .A2(new_n261), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n236), .A2(G1698), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n254), .A2(new_n327), .A3(new_n256), .A4(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(G33), .A2(G97), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT68), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n329), .A2(KEYINPUT68), .A3(new_n330), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n333), .A2(new_n259), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT13), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n268), .B1(new_n300), .B2(G238), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n336), .B1(new_n335), .B2(new_n337), .ZN(new_n340));
  OAI21_X1  g0140(.A(G200), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n340), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(G190), .A3(new_n338), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n326), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n265), .A2(new_n276), .ZN(new_n345));
  INV_X1    g0145(.A(G179), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n347), .B(new_n304), .C1(G169), .C2(new_n345), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n310), .A2(new_n344), .A3(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(G169), .B1(new_n339), .B2(new_n340), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT14), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n342), .A2(G179), .A3(new_n338), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT14), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n353), .B(G169), .C1(new_n339), .C2(new_n340), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n351), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n325), .ZN(new_n356));
  OAI22_X1  g0156(.A1(new_n252), .A2(new_n282), .B1(new_n281), .B2(new_n313), .ZN(new_n357));
  XNOR2_X1  g0157(.A(KEYINPUT15), .B(G87), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(new_n283), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n286), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n291), .A2(G77), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n360), .B(new_n361), .C1(new_n218), .C2(new_n293), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT67), .ZN(new_n363));
  OR2_X1    g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n363), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n260), .A2(G1698), .ZN(new_n367));
  INV_X1    g0167(.A(G107), .ZN(new_n368));
  OAI22_X1  g0168(.A1(new_n367), .A2(new_n222), .B1(new_n368), .B2(new_n260), .ZN(new_n369));
  NOR3_X1   g0169(.A1(new_n257), .A2(new_n236), .A3(G1698), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n259), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n300), .A2(G244), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(new_n269), .A3(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G169), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n366), .B(new_n375), .C1(G179), .C2(new_n373), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n349), .A2(new_n356), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n366), .ZN(new_n378));
  INV_X1    g0178(.A(new_n373), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(G190), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n373), .A2(G200), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n378), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n293), .A2(new_n281), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n291), .B2(new_n281), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n271), .B(G232), .C1(new_n274), .C2(new_n266), .ZN(new_n385));
  INV_X1    g0185(.A(G190), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n385), .A2(new_n386), .A3(new_n269), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n254), .A2(new_n256), .A3(G223), .A4(new_n261), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n254), .A2(new_n256), .A3(G226), .A4(G1698), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G33), .A2(G87), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT73), .ZN(new_n392));
  AND3_X1   g0192(.A1(new_n391), .A2(new_n392), .A3(new_n259), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n392), .B1(new_n391), .B2(new_n259), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n387), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n391), .A2(new_n259), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(new_n385), .A3(new_n269), .ZN(new_n397));
  INV_X1    g0197(.A(G200), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT71), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n255), .B2(KEYINPUT3), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n253), .A2(KEYINPUT71), .A3(G33), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(new_n256), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT7), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n405), .A2(G20), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT72), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n405), .B1(new_n260), .B2(G20), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT72), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n404), .A2(new_n410), .A3(new_n406), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n408), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(G68), .ZN(new_n413));
  XNOR2_X1  g0213(.A(G58), .B(G68), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(G20), .B1(G159), .B2(new_n279), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT16), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT70), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n417), .B(new_n405), .C1(new_n260), .C2(G20), .ZN(new_n418));
  AOI21_X1  g0218(.A(G20), .B1(new_n254), .B2(new_n256), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT70), .B1(new_n419), .B2(KEYINPUT7), .ZN(new_n420));
  NOR3_X1   g0220(.A1(new_n260), .A2(new_n405), .A3(G20), .ZN(new_n421));
  OAI211_X1 g0221(.A(G68), .B(new_n418), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n422), .A2(KEYINPUT16), .A3(new_n415), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n286), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n384), .B(new_n400), .C1(new_n416), .C2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT17), .ZN(new_n426));
  INV_X1    g0226(.A(new_n415), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(new_n412), .B2(G68), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n286), .B(new_n423), .C1(new_n428), .C2(KEYINPUT16), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT17), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n429), .A2(new_n430), .A3(new_n384), .A4(new_n400), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n429), .A2(new_n384), .ZN(new_n433));
  AND3_X1   g0233(.A1(new_n385), .A2(new_n346), .A3(new_n269), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n393), .B2(new_n394), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n397), .A2(new_n374), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT18), .B1(new_n433), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT18), .ZN(new_n440));
  AOI211_X1 g0240(.A(new_n440), .B(new_n437), .C1(new_n429), .C2(new_n384), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n382), .B(new_n432), .C1(new_n439), .C2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT74), .ZN(new_n443));
  OR3_X1    g0243(.A1(new_n377), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n443), .B1(new_n377), .B2(new_n442), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(G45), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n447), .B1(new_n288), .B2(new_n289), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n259), .B1(new_n448), .B2(new_n267), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(G250), .B2(new_n448), .ZN(new_n450));
  NOR3_X1   g0250(.A1(new_n257), .A2(new_n222), .A3(G1698), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n254), .A2(new_n256), .A3(G244), .A4(G1698), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G33), .A2(G116), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n259), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n450), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(KEYINPUT76), .B1(new_n456), .B2(G179), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT19), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n282), .B1(new_n330), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(G97), .A2(G107), .ZN(new_n460));
  INV_X1    g0260(.A(G87), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT77), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n260), .A2(new_n282), .A3(G68), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT77), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n459), .A2(new_n462), .A3(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n458), .B1(new_n283), .B2(new_n209), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n464), .A2(new_n465), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n469), .A2(new_n286), .B1(new_n294), .B2(new_n358), .ZN(new_n470));
  INV_X1    g0270(.A(new_n286), .ZN(new_n471));
  OAI21_X1  g0271(.A(G33), .B1(new_n272), .B2(new_n273), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n293), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  OR2_X1    g0273(.A1(new_n473), .A2(new_n358), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n456), .A2(new_n374), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT76), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n450), .A2(new_n455), .A3(new_n477), .A4(new_n346), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n457), .A2(new_n475), .A3(new_n476), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n456), .A2(G200), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n450), .A2(new_n455), .A3(G190), .ZN(new_n481));
  INV_X1    g0281(.A(new_n473), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G87), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n480), .A2(new_n481), .A3(new_n470), .A4(new_n483), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT24), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n254), .A2(new_n256), .A3(new_n282), .A4(G87), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT81), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT81), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n260), .A2(new_n489), .A3(new_n282), .A4(G87), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n488), .A2(new_n490), .A3(KEYINPUT22), .ZN(new_n491));
  AOI21_X1  g0291(.A(KEYINPUT22), .B1(new_n488), .B2(new_n490), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT23), .B1(new_n282), .B2(G107), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT23), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n495), .A2(new_n368), .A3(G20), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n282), .A2(G33), .A3(G116), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n494), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT82), .ZN(new_n499));
  XNOR2_X1  g0299(.A(new_n498), .B(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n486), .B1(new_n493), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n488), .A2(new_n490), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT22), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n488), .A2(new_n490), .A3(KEYINPUT22), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n504), .A2(new_n500), .A3(new_n486), .A4(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n286), .B1(new_n501), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n260), .A2(G250), .A3(new_n261), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n367), .B2(new_n210), .ZN(new_n510));
  XOR2_X1   g0310(.A(KEYINPUT84), .B(G294), .Z(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n512), .A2(new_n255), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n259), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(G45), .B1(new_n272), .B2(new_n273), .ZN(new_n515));
  AND2_X1   g0315(.A1(KEYINPUT5), .A2(G41), .ZN(new_n516));
  NOR2_X1   g0316(.A1(KEYINPUT5), .A2(G41), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n271), .B(G264), .C1(new_n515), .C2(new_n518), .ZN(new_n519));
  OR2_X1    g0319(.A1(new_n516), .A2(new_n517), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n448), .A2(new_n520), .A3(new_n271), .A4(G274), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n514), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n398), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n514), .A2(new_n386), .A3(new_n519), .A4(new_n521), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n473), .A2(new_n368), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT83), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n528), .A2(KEYINPUT25), .ZN(new_n529));
  NOR3_X1   g0329(.A1(new_n293), .A2(G107), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(KEYINPUT25), .ZN(new_n531));
  XNOR2_X1  g0331(.A(new_n530), .B(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n508), .A2(new_n525), .A3(new_n527), .A4(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n485), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n522), .A2(new_n374), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(G179), .B2(new_n522), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n504), .A2(new_n500), .A3(new_n505), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT24), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n506), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n526), .B1(new_n540), .B2(new_n286), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n537), .B1(new_n541), .B2(new_n533), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n535), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n368), .A2(KEYINPUT6), .A3(G97), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n209), .A2(new_n368), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n545), .A2(new_n460), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n544), .B1(new_n546), .B2(KEYINPUT6), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(G20), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n313), .A2(new_n246), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n404), .A2(new_n410), .A3(new_n406), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n410), .B1(new_n404), .B2(new_n406), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n419), .A2(KEYINPUT7), .ZN(new_n553));
  NOR3_X1   g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n548), .B(new_n550), .C1(new_n554), .C2(new_n368), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n555), .A2(new_n286), .B1(new_n209), .B2(new_n294), .ZN(new_n556));
  NAND2_X1  g0356(.A1(G33), .A2(G283), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n254), .A2(new_n256), .A3(G244), .A4(new_n261), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT4), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n260), .A2(KEYINPUT4), .A3(G244), .A4(new_n261), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n254), .A2(new_n256), .A3(G250), .A4(G1698), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(KEYINPUT75), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT75), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n260), .A2(new_n565), .A3(G250), .A4(G1698), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n561), .A2(new_n562), .A3(new_n564), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n259), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n271), .B(G257), .C1(new_n515), .C2(new_n518), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n568), .A2(new_n386), .A3(new_n521), .A4(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n569), .ZN(new_n571));
  INV_X1    g0371(.A(new_n521), .ZN(new_n572));
  AOI211_X1 g0372(.A(new_n571), .B(new_n572), .C1(new_n567), .C2(new_n259), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n570), .B1(new_n573), .B2(G200), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n482), .A2(G97), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n556), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n568), .A2(new_n346), .A3(new_n521), .A4(new_n569), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n573), .B2(G169), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n578), .B1(new_n556), .B2(new_n575), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n285), .A2(new_n229), .B1(G20), .B2(new_n215), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n557), .B(new_n282), .C1(G33), .C2(new_n209), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT20), .ZN(new_n584));
  OR2_X1    g0384(.A1(new_n584), .A2(KEYINPUT78), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(KEYINPUT78), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n583), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n581), .A2(KEYINPUT78), .A3(new_n582), .A4(new_n584), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n290), .A2(G13), .A3(G20), .A4(new_n215), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n293), .A2(new_n471), .A3(new_n472), .A4(G116), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n587), .A2(new_n588), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n261), .A2(G257), .ZN(new_n592));
  NAND2_X1  g0392(.A1(G264), .A2(G1698), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n254), .A2(new_n256), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n594), .B(new_n259), .C1(G303), .C2(new_n260), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n271), .B(G270), .C1(new_n515), .C2(new_n518), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(new_n521), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n591), .A2(G169), .A3(new_n597), .ZN(new_n598));
  XOR2_X1   g0398(.A(KEYINPUT80), .B(KEYINPUT21), .Z(new_n599));
  NOR2_X1   g0399(.A1(new_n597), .A2(new_n346), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n598), .A2(new_n599), .B1(new_n600), .B2(new_n591), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n591), .A2(KEYINPUT21), .A3(new_n597), .A4(G169), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT79), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n602), .A2(new_n603), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n601), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n591), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n597), .A2(new_n386), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n609), .B1(G200), .B2(new_n597), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n607), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  AND4_X1   g0411(.A1(new_n446), .A2(new_n543), .A3(new_n580), .A4(new_n611), .ZN(G372));
  NOR2_X1   g0412(.A1(new_n439), .A2(new_n441), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n356), .A2(new_n376), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n432), .A2(new_n344), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n310), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n348), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n446), .ZN(new_n620));
  OAI21_X1  g0420(.A(KEYINPUT85), .B1(new_n542), .B2(new_n607), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT85), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n598), .A2(new_n599), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n600), .A2(new_n591), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n606), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n625), .B1(new_n626), .B2(new_n604), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n471), .B1(new_n539), .B2(new_n506), .ZN(new_n628));
  NOR3_X1   g0428(.A1(new_n628), .A2(new_n526), .A3(new_n532), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n622), .B(new_n627), .C1(new_n629), .C2(new_n537), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n475), .B(new_n476), .C1(G179), .C2(new_n456), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n484), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n632), .B1(new_n629), .B2(new_n525), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n621), .A2(new_n580), .A3(new_n630), .A4(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n555), .A2(new_n286), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n294), .A2(new_n209), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(new_n636), .A3(new_n575), .ZN(new_n637));
  INV_X1    g0437(.A(new_n578), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n479), .A2(new_n484), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT26), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n631), .A2(new_n484), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT26), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n579), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n641), .A2(new_n631), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n634), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n619), .B1(new_n620), .B2(new_n647), .ZN(G369));
  INV_X1    g0448(.A(G13), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(G20), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n290), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n651), .B(KEYINPUT86), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT27), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(G213), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(G343), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n591), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n611), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n607), .A2(new_n591), .A3(new_n658), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G330), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT87), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n508), .A2(new_n527), .A3(new_n533), .ZN(new_n666));
  INV_X1    g0466(.A(new_n537), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(new_n658), .ZN(new_n669));
  INV_X1    g0469(.A(new_n658), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n534), .B1(new_n629), .B2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n669), .B1(new_n668), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n665), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n627), .A2(new_n658), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT88), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(new_n669), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n673), .A2(new_n678), .ZN(G399));
  NOR2_X1   g0479(.A1(new_n462), .A2(G116), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n226), .A2(new_n270), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G1), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n232), .B2(new_n681), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT28), .ZN(new_n684));
  OAI21_X1  g0484(.A(KEYINPUT26), .B1(new_n639), .B2(new_n632), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n579), .A2(new_n485), .A3(new_n643), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(new_n631), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT89), .B1(new_n576), .B2(new_n579), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT89), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n556), .A2(new_n574), .A3(new_n575), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n639), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n668), .A2(new_n627), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n693), .A2(new_n633), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n687), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT29), .B1(new_n695), .B2(new_n658), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n658), .B1(new_n634), .B2(new_n645), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT29), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n543), .A2(new_n580), .A3(new_n611), .A4(new_n670), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n514), .A2(new_n519), .ZN(new_n703));
  INV_X1    g0503(.A(new_n456), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n573), .A2(new_n703), .A3(new_n704), .A4(new_n600), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT30), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n573), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n597), .A2(new_n346), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n708), .A2(new_n456), .A3(new_n522), .A4(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n705), .A2(new_n706), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n707), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n658), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT31), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n712), .A2(KEYINPUT31), .A3(new_n658), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n702), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G330), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n701), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n684), .B1(new_n720), .B2(G1), .ZN(G364));
  INV_X1    g0521(.A(G1), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n722), .B1(new_n650), .B2(G45), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n681), .ZN(new_n724));
  OAI211_X1 g0524(.A(new_n664), .B(new_n724), .C1(G330), .C2(new_n662), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n282), .A2(G190), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT94), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n398), .A2(G179), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n729), .A2(KEYINPUT95), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(KEYINPUT95), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n368), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT93), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n386), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n736), .A2(G190), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI22_X1  g0540(.A1(new_n202), .A2(new_n738), .B1(new_n740), .B2(new_n221), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G179), .A2(G200), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n727), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(KEYINPUT32), .A3(G159), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT32), .ZN(new_n746));
  INV_X1    g0546(.A(G159), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n746), .B1(new_n743), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n741), .B1(new_n745), .B2(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n282), .B1(new_n742), .B2(G190), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT96), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G97), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n282), .A2(new_n386), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n346), .A2(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G58), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n754), .A2(new_n728), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n260), .B1(new_n756), .B2(new_n757), .C1(new_n461), .C2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n755), .A2(new_n726), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n760), .A2(KEYINPUT92), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(KEYINPUT92), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n759), .B1(new_n764), .B2(new_n218), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n734), .A2(new_n749), .A3(new_n753), .A4(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n732), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n743), .A2(KEYINPUT97), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n743), .A2(KEYINPUT97), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n767), .A2(G283), .B1(new_n771), .B2(G329), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n737), .A2(G326), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n512), .A2(new_n750), .ZN(new_n774));
  INV_X1    g0574(.A(G311), .ZN(new_n775));
  INV_X1    g0575(.A(G303), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n257), .B1(new_n760), .B2(new_n775), .C1(new_n776), .C2(new_n758), .ZN(new_n777));
  XNOR2_X1  g0577(.A(KEYINPUT33), .B(G317), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n774), .B(new_n777), .C1(new_n739), .C2(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n772), .A2(new_n773), .A3(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G322), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n756), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n766), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n229), .B1(G20), .B2(new_n374), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G13), .A2(G33), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G20), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n784), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n260), .A2(G355), .A3(new_n226), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n257), .A2(new_n226), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT90), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(G45), .B2(new_n232), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT91), .Z(new_n793));
  NOR2_X1   g0593(.A1(new_n247), .A2(new_n447), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n789), .B1(G116), .B2(new_n226), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n783), .A2(new_n784), .B1(new_n788), .B2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n724), .ZN(new_n797));
  INV_X1    g0597(.A(new_n787), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n796), .B(new_n797), .C1(new_n662), .C2(new_n798), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n725), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(G396));
  NOR2_X1   g0601(.A1(new_n376), .A2(new_n658), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n382), .B1(new_n378), .B2(new_n670), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n802), .B1(new_n803), .B2(new_n376), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n697), .B(new_n804), .Z(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(new_n718), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(new_n724), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n764), .A2(G116), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G283), .A2(new_n739), .B1(new_n737), .B2(G303), .ZN(new_n809));
  INV_X1    g0609(.A(new_n756), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n260), .B1(new_n810), .B2(G294), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n808), .A2(new_n809), .A3(new_n753), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n767), .A2(G87), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n775), .B2(new_n770), .ZN(new_n814));
  INV_X1    g0614(.A(new_n758), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n812), .B(new_n814), .C1(G107), .C2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(G50), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n767), .A2(G68), .ZN(new_n818));
  INV_X1    g0618(.A(new_n750), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n257), .B1(new_n819), .B2(G58), .ZN(new_n820));
  INV_X1    g0620(.A(G132), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n818), .B(new_n820), .C1(new_n821), .C2(new_n770), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n764), .A2(G159), .B1(G137), .B2(new_n737), .ZN(new_n823));
  INV_X1    g0623(.A(G143), .ZN(new_n824));
  INV_X1    g0624(.A(G150), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n823), .B1(new_n824), .B2(new_n756), .C1(new_n825), .C2(new_n740), .ZN(new_n826));
  XNOR2_X1  g0626(.A(KEYINPUT98), .B(KEYINPUT34), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n826), .A2(new_n827), .ZN(new_n829));
  NOR3_X1   g0629(.A1(new_n822), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n816), .B1(new_n817), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n784), .A2(new_n785), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n832), .A2(new_n784), .B1(new_n246), .B2(new_n833), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n834), .B(new_n797), .C1(new_n786), .C2(new_n804), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n807), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(G384));
  OAI211_X1 g0637(.A(G20), .B(new_n230), .C1(new_n547), .C2(KEYINPUT35), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n215), .B(new_n838), .C1(KEYINPUT35), .C2(new_n547), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT36), .Z(new_n840));
  OAI21_X1  g0640(.A(new_n218), .B1(new_n757), .B2(new_n221), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n841), .A2(new_n232), .B1(G50), .B2(new_n221), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n842), .A2(new_n649), .A3(new_n274), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT99), .Z(new_n845));
  NAND3_X1  g0645(.A1(new_n713), .A2(KEYINPUT103), .A3(new_n714), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n714), .A2(KEYINPUT103), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n712), .A2(new_n658), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n702), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n356), .A2(new_n344), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n850), .A2(new_n325), .A3(new_n658), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n356), .B(new_n344), .C1(new_n326), .C2(new_n670), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT40), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n849), .A2(new_n853), .A3(new_n854), .A4(new_n804), .ZN(new_n855));
  INV_X1    g0655(.A(new_n425), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n429), .A2(new_n384), .B1(new_n656), .B2(new_n437), .ZN(new_n857));
  NOR3_X1   g0657(.A1(new_n856), .A2(new_n857), .A3(KEYINPUT37), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT16), .B1(new_n422), .B2(new_n415), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n384), .B1(new_n424), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n656), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT100), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n860), .A2(new_n861), .A3(KEYINPUT100), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n860), .A2(new_n438), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n864), .A2(new_n425), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n858), .B1(new_n867), .B2(KEYINPUT37), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n384), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n415), .B1(new_n554), .B2(new_n221), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT16), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n423), .A2(new_n286), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n870), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n440), .B1(new_n875), .B2(new_n437), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n433), .A2(KEYINPUT18), .A3(new_n438), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n876), .A2(new_n877), .B1(new_n426), .B2(new_n431), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n864), .A2(new_n865), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n878), .A2(new_n879), .A3(KEYINPUT101), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT101), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n432), .B1(new_n439), .B2(new_n441), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n864), .A2(new_n865), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n869), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT101), .B1(new_n878), .B2(new_n879), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n882), .A2(new_n881), .A3(new_n883), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n868), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT38), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n855), .B1(new_n887), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n882), .A2(new_n433), .A3(new_n861), .ZN(new_n894));
  INV_X1    g0694(.A(new_n858), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT37), .B1(new_n856), .B2(new_n857), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT38), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n890), .B2(KEYINPUT38), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n849), .A2(new_n853), .A3(new_n804), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT40), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n893), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n446), .A2(new_n849), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n902), .B(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(G330), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n618), .B1(new_n700), .B2(new_n446), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n906), .B(KEYINPUT104), .Z(new_n907));
  XNOR2_X1  g0707(.A(new_n905), .B(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n887), .A2(new_n891), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n851), .A2(new_n852), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n607), .B1(new_n666), .B2(new_n667), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n580), .B1(new_n911), .B2(new_n622), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n630), .A2(new_n633), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n641), .A2(new_n631), .A3(new_n644), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n670), .B(new_n804), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n802), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n910), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n909), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n613), .A2(new_n656), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT102), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT102), .ZN(new_n922));
  INV_X1    g0722(.A(new_n920), .ZN(new_n923));
  AOI211_X1 g0723(.A(new_n922), .B(new_n923), .C1(new_n909), .C2(new_n918), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n356), .A2(new_n658), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  AOI211_X1 g0726(.A(new_n886), .B(new_n868), .C1(new_n888), .C2(new_n889), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n888), .A2(new_n889), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT38), .B1(new_n928), .B2(new_n869), .ZN(new_n929));
  OAI21_X1  g0729(.A(KEYINPUT39), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT39), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n899), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n926), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n921), .A2(new_n924), .A3(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n908), .B(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n290), .A2(new_n650), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n845), .B1(new_n935), .B2(new_n936), .ZN(G367));
  INV_X1    g0737(.A(new_n673), .ZN(new_n938));
  INV_X1    g0738(.A(new_n637), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n692), .B1(new_n939), .B2(new_n670), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n579), .A2(new_n658), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n677), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT42), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n940), .A2(new_n668), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n658), .B1(new_n945), .B2(new_n639), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n470), .A2(new_n483), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n658), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n642), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n631), .B2(new_n949), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(KEYINPUT43), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n938), .B(new_n942), .C1(new_n947), .C2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n938), .A2(new_n942), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n955), .B(new_n952), .C1(new_n946), .C2(new_n944), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n951), .A2(KEYINPUT43), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n957), .B(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n681), .B(KEYINPUT41), .Z(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n664), .A2(KEYINPUT106), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n672), .A2(new_n675), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n962), .A2(new_n676), .A3(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n664), .A2(KEYINPUT106), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n964), .B(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(KEYINPUT107), .B1(new_n967), .B2(new_n719), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n964), .B(new_n965), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT107), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n969), .A2(new_n970), .A3(new_n720), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n678), .A2(new_n942), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT44), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n678), .A2(new_n942), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT45), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n977), .A2(KEYINPUT105), .A3(new_n938), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n938), .A2(KEYINPUT105), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n973), .A2(new_n979), .A3(new_n976), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n968), .A2(new_n971), .A3(new_n978), .A4(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n961), .B1(new_n981), .B2(new_n720), .ZN(new_n982));
  INV_X1    g0782(.A(new_n723), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n959), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n260), .B1(new_n764), .B2(G283), .ZN(new_n985));
  INV_X1    g0785(.A(G317), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n985), .B1(new_n368), .B2(new_n750), .C1(new_n986), .C2(new_n743), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(new_n511), .B2(new_n739), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n815), .A2(G116), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT46), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n737), .A2(G311), .B1(G303), .B2(new_n810), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT108), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n767), .A2(G97), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n988), .A2(new_n990), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT109), .Z(new_n995));
  AOI21_X1  g0795(.A(new_n257), .B1(new_n815), .B2(G58), .ZN(new_n996));
  INV_X1    g0796(.A(G137), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n996), .B1(new_n743), .B2(new_n997), .C1(new_n763), .C2(new_n202), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(new_n767), .B2(new_n218), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n751), .A2(new_n221), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n747), .B2(new_n740), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(G143), .B2(new_n737), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n999), .B(new_n1003), .C1(new_n825), .C2(new_n756), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT110), .Z(new_n1005));
  NOR2_X1   g0805(.A1(new_n995), .A2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT47), .Z(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n784), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n791), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n788), .B1(new_n226), .B2(new_n358), .C1(new_n242), .C2(new_n1009), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n951), .A2(new_n798), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1008), .A2(new_n797), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n984), .A2(new_n1012), .ZN(G387));
  NAND2_X1  g0813(.A1(new_n968), .A2(new_n971), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n681), .B(KEYINPUT113), .Z(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1014), .B(new_n1016), .C1(new_n720), .C2(new_n969), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n764), .A2(G303), .B1(G322), .B2(new_n737), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n775), .B2(new_n740), .C1(new_n986), .C2(new_n756), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT48), .ZN(new_n1020));
  INV_X1    g0820(.A(G283), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1020), .B1(new_n1021), .B2(new_n750), .C1(new_n512), .C2(new_n758), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT49), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n744), .A2(G326), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n260), .B1(new_n767), .B2(G116), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n760), .A2(new_n221), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n751), .A2(new_n358), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G159), .B2(new_n737), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n257), .B1(new_n810), .B2(G50), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n815), .A2(new_n218), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1032), .B(new_n1033), .C1(new_n743), .C2(new_n825), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n281), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1034), .B1(new_n1035), .B2(new_n739), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n993), .A2(new_n1031), .A3(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1028), .B1(new_n1029), .B2(new_n1037), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT112), .Z(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n784), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n672), .A2(new_n798), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n791), .B1(new_n239), .B2(new_n447), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n680), .B(new_n447), .C1(new_n221), .C2(new_n246), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT50), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n281), .B2(G50), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1035), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1043), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1042), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n260), .A2(new_n226), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n1049), .A2(new_n680), .B1(G107), .B2(new_n226), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT111), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n724), .B(new_n1041), .C1(new_n788), .C2(new_n1052), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n1040), .A2(new_n1053), .B1(new_n969), .B2(new_n983), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1017), .A2(new_n1054), .ZN(G393));
  NAND2_X1  g0855(.A1(new_n977), .A2(new_n938), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n973), .A2(new_n673), .A3(new_n976), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1058), .A2(new_n723), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n788), .B1(new_n209), .B2(new_n226), .C1(new_n250), .C2(new_n1009), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n260), .B1(new_n743), .B2(new_n824), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n740), .A2(new_n202), .B1(new_n246), .B2(new_n751), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(new_n1035), .C2(new_n764), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n815), .A2(G68), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n737), .A2(G150), .B1(G159), .B2(new_n810), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT51), .Z(new_n1066));
  NAND4_X1  g0866(.A1(new_n813), .A2(new_n1063), .A3(new_n1064), .A4(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n260), .B1(new_n815), .B2(G283), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(new_n215), .B2(new_n750), .C1(new_n743), .C2(new_n781), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(G303), .B2(new_n739), .ZN(new_n1070));
  INV_X1    g0870(.A(G294), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n734), .B(new_n1070), .C1(new_n1071), .C2(new_n760), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n737), .A2(G317), .B1(G311), .B2(new_n810), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT114), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT52), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1067), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n724), .B1(new_n1076), .B2(new_n784), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1060), .B(new_n1077), .C1(new_n942), .C2(new_n798), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1059), .A2(new_n1079), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n1014), .A2(new_n1058), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n981), .A2(new_n1016), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(G390));
  AOI21_X1  g0883(.A(new_n802), .B1(new_n697), .B2(new_n804), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n926), .B1(new_n1084), .B2(new_n910), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1085), .A2(new_n930), .A3(new_n932), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n898), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n891), .A2(new_n1087), .ZN(new_n1088));
  AND3_X1   g0888(.A1(new_n685), .A2(new_n631), .A3(new_n686), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n688), .A2(new_n693), .A3(new_n633), .A4(new_n691), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n658), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n803), .A2(new_n376), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n802), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1088), .B(new_n926), .C1(new_n910), .C2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n717), .A2(new_n853), .A3(G330), .A4(new_n804), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1086), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT115), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1086), .A2(new_n1094), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n849), .A2(new_n853), .A3(G330), .A4(new_n804), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1086), .A2(KEYINPUT115), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1098), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1084), .ZN(new_n1105));
  AND3_X1   g0905(.A1(new_n717), .A2(G330), .A3(new_n804), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1100), .B1(new_n1106), .B2(new_n853), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1095), .A2(new_n1093), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n849), .A2(G330), .A3(new_n804), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n910), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1105), .A2(new_n1107), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n445), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n377), .A2(new_n442), .A3(new_n443), .ZN(new_n1113));
  OAI211_X1 g0913(.A(G330), .B(new_n849), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT116), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n446), .A2(KEYINPUT116), .A3(G330), .A4(new_n849), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n906), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1111), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1104), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1098), .A2(new_n1120), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1122), .A2(new_n1016), .A3(new_n1123), .ZN(new_n1124));
  OR2_X1    g0924(.A1(new_n1104), .A2(new_n723), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n930), .A2(new_n932), .A3(new_n785), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n833), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1127), .A2(new_n1035), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n771), .A2(G294), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n257), .B1(new_n215), .B2(new_n756), .C1(new_n763), .C2(new_n209), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(G87), .B2(new_n815), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n368), .A2(new_n740), .B1(new_n738), .B2(new_n1021), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(G77), .B2(new_n752), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n818), .A2(new_n1129), .A3(new_n1131), .A4(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n758), .A2(new_n825), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT53), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(KEYINPUT54), .B(G143), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1136), .B(new_n260), .C1(new_n763), .C2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n771), .B2(G125), .ZN(new_n1139));
  INV_X1    g0939(.A(G128), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n738), .A2(new_n1140), .B1(new_n747), .B2(new_n751), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(G137), .B2(new_n739), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1139), .B(new_n1142), .C1(new_n202), .C2(new_n732), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n756), .A2(new_n821), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1134), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n724), .B(new_n1128), .C1(new_n1145), .C2(new_n784), .ZN(new_n1146));
  XOR2_X1   g0946(.A(new_n1146), .B(KEYINPUT117), .Z(new_n1147));
  NAND2_X1  g0947(.A1(new_n1126), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1124), .A2(new_n1125), .A3(new_n1148), .ZN(G378));
  NAND2_X1  g0949(.A1(new_n861), .A2(new_n304), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n310), .A2(new_n348), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n1152), .A2(KEYINPUT55), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1152), .A2(KEYINPUT55), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1151), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  OR2_X1    g0955(.A1(new_n1152), .A2(KEYINPUT55), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1152), .A2(KEYINPUT55), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1156), .A2(new_n1157), .A3(new_n1150), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1155), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1159), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT121), .ZN(new_n1163));
  NOR3_X1   g0963(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1159), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(KEYINPUT121), .B1(new_n1167), .B2(new_n1160), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1164), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n785), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n833), .A2(new_n202), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1001), .B1(new_n770), .B2(new_n1021), .C1(new_n732), .C2(new_n757), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n737), .A2(G116), .ZN(new_n1173));
  AOI21_X1  g0973(.A(G41), .B1(new_n810), .B2(G107), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1173), .A2(new_n257), .A3(new_n1033), .A4(new_n1174), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n740), .A2(new_n209), .B1(new_n358), .B2(new_n760), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT118), .ZN(new_n1177));
  NOR3_X1   g0977(.A1(new_n1172), .A2(new_n1175), .A3(new_n1177), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT58), .Z(new_n1179));
  AOI21_X1  g0979(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1180));
  AOI21_X1  g0980(.A(G33), .B1(new_n744), .B2(G124), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1181), .B(new_n270), .C1(new_n732), .C2(new_n747), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT119), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n1140), .A2(new_n756), .B1(new_n758), .B2(new_n1137), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n752), .B2(G150), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(G125), .A2(new_n737), .B1(new_n739), .B2(G132), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1185), .B(new_n1186), .C1(new_n997), .C2(new_n760), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT59), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1179), .B1(G50), .B2(new_n1180), .C1(new_n1183), .C2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n724), .B1(new_n1189), .B2(new_n784), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1170), .A2(new_n1171), .A3(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n900), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n854), .B1(new_n1088), .B2(new_n1193), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1169), .B(G330), .C1(new_n1194), .C2(new_n892), .ZN(new_n1195));
  INV_X1    g0995(.A(G330), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n893), .B2(new_n901), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1195), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT122), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1200), .B1(new_n934), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n919), .A2(new_n920), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n922), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n933), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n919), .A2(KEYINPUT102), .A3(new_n920), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(G330), .B1(new_n1194), .B2(new_n892), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n1198), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1207), .A2(KEYINPUT122), .A3(new_n1209), .A4(new_n1195), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1202), .A2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1192), .B1(new_n1211), .B2(new_n983), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1119), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1123), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n934), .A2(new_n1209), .A3(new_n1195), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1200), .A2(new_n1207), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1216), .A2(new_n1217), .A3(KEYINPUT57), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1016), .B1(new_n1215), .B2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(KEYINPUT57), .B1(new_n1211), .B2(new_n1214), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1212), .B1(new_n1219), .B2(new_n1220), .ZN(G375));
  AOI22_X1  g1021(.A1(new_n767), .A2(G77), .B1(new_n771), .B2(G303), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n257), .B1(new_n209), .B2(new_n758), .C1(new_n763), .C2(new_n368), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n215), .A2(new_n740), .B1(new_n738), .B2(new_n1071), .ZN(new_n1224));
  NOR3_X1   g1024(.A1(new_n1223), .A2(new_n1224), .A3(new_n1030), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1222), .B(new_n1225), .C1(new_n1021), .C2(new_n756), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n756), .A2(new_n997), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n767), .A2(G58), .B1(new_n771), .B2(G128), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n751), .A2(new_n202), .B1(new_n825), .B2(new_n760), .ZN(new_n1229));
  XOR2_X1   g1029(.A(new_n1229), .B(KEYINPUT123), .Z(new_n1230));
  OAI221_X1 g1030(.A(new_n260), .B1(new_n758), .B2(new_n747), .C1(new_n740), .C2(new_n1137), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(G132), .B2(new_n737), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1228), .A2(new_n1230), .A3(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1226), .B1(new_n1227), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n784), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(G68), .B2(new_n1127), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n724), .B(new_n1236), .C1(new_n910), .C2(new_n785), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1111), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1237), .B1(new_n1238), .B2(new_n983), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1111), .A2(new_n1119), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n960), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1239), .B1(new_n1241), .B2(new_n1120), .ZN(G381));
  NOR4_X1   g1042(.A1(G387), .A2(G396), .A3(G393), .A4(G390), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(G375), .A2(G378), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(G384), .A2(G381), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .ZN(G407));
  NAND2_X1  g1046(.A1(new_n657), .A2(G213), .ZN(new_n1247));
  XOR2_X1   g1047(.A(new_n1247), .B(KEYINPUT124), .Z(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1244), .A2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(G407), .A2(G213), .A3(new_n1250), .ZN(G409));
  OAI211_X1 g1051(.A(G378), .B(new_n1212), .C1(new_n1219), .C2(new_n1220), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1124), .A2(new_n1125), .A3(new_n1148), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1211), .A2(new_n960), .A3(new_n1214), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1216), .A2(new_n1217), .A3(new_n983), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1254), .A2(new_n1191), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1252), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT60), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1015), .B1(new_n1240), .B2(new_n1259), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1260), .B(new_n1121), .C1(new_n1259), .C2(new_n1240), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1261), .A2(G384), .A3(new_n1239), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(G384), .B1(new_n1261), .B2(new_n1239), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1258), .A2(KEYINPUT63), .A3(new_n1248), .A4(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT127), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1249), .B1(new_n1252), .B2(new_n1257), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1269), .A2(KEYINPUT127), .A3(KEYINPUT63), .A4(new_n1265), .ZN(new_n1270));
  AOI21_X1  g1070(.A(KEYINPUT61), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT63), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT125), .ZN(new_n1273));
  AND4_X1   g1073(.A1(new_n1273), .A2(new_n1258), .A3(new_n1247), .A4(new_n1265), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1247), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(new_n1252), .B2(new_n1257), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1273), .B1(new_n1276), .B2(new_n1265), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1272), .B1(new_n1274), .B2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(G390), .B1(new_n984), .B2(new_n1012), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(G393), .A2(G396), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n800), .B1(new_n1017), .B2(new_n1054), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n984), .A2(new_n1012), .A3(G390), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1280), .A2(new_n1283), .A3(new_n1284), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n984), .A2(new_n1012), .A3(G390), .ZN(new_n1286));
  OAI22_X1  g1086(.A1(new_n1286), .A2(new_n1279), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT126), .ZN(new_n1289));
  OR2_X1    g1089(.A1(new_n1276), .A2(new_n1289), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1265), .A2(new_n1248), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1275), .A2(G2897), .ZN(new_n1292));
  AOI22_X1  g1092(.A1(new_n1291), .A2(G2897), .B1(new_n1265), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1276), .A2(new_n1289), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1290), .A2(new_n1293), .A3(new_n1294), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1271), .A2(new_n1278), .A3(new_n1288), .A4(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1269), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1293), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT61), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT62), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1301), .B1(new_n1274), .B2(new_n1277), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1269), .A2(KEYINPUT62), .A3(new_n1265), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1300), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1296), .B1(new_n1304), .B2(new_n1288), .ZN(G405));
  NAND2_X1  g1105(.A1(G375), .A2(new_n1253), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1252), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1265), .ZN(new_n1308));
  XNOR2_X1  g1108(.A(new_n1307), .B(new_n1308), .ZN(new_n1309));
  XNOR2_X1  g1109(.A(new_n1288), .B(new_n1309), .ZN(G402));
endmodule


