

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585;

  NOR2_X1 U324 ( .A1(n549), .A2(n525), .ZN(n531) );
  XNOR2_X1 U325 ( .A(n430), .B(n429), .ZN(n547) );
  XNOR2_X1 U326 ( .A(KEYINPUT101), .B(KEYINPUT37), .ZN(n473) );
  XNOR2_X1 U327 ( .A(KEYINPUT90), .B(n467), .ZN(n518) );
  XOR2_X1 U328 ( .A(n305), .B(n304), .Z(n292) );
  XNOR2_X1 U329 ( .A(KEYINPUT54), .B(KEYINPUT124), .ZN(n432) );
  XNOR2_X1 U330 ( .A(KEYINPUT48), .B(KEYINPUT117), .ZN(n429) );
  XNOR2_X1 U331 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U332 ( .A(n306), .B(n292), .ZN(n307) );
  XNOR2_X1 U333 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U334 ( .A(n474), .B(n473), .ZN(n517) );
  NOR2_X1 U335 ( .A1(n533), .A2(n452), .ZN(n568) );
  XOR2_X1 U336 ( .A(n363), .B(n362), .Z(n521) );
  XNOR2_X1 U337 ( .A(KEYINPUT126), .B(G183GAT), .ZN(n453) );
  XNOR2_X1 U338 ( .A(n478), .B(G43GAT), .ZN(n479) );
  XNOR2_X1 U339 ( .A(n454), .B(n453), .ZN(G1350GAT) );
  XNOR2_X1 U340 ( .A(n480), .B(n479), .ZN(G1330GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT76), .B(KEYINPUT79), .Z(n294) );
  XNOR2_X1 U342 ( .A(KEYINPUT75), .B(KEYINPUT78), .ZN(n293) );
  XNOR2_X1 U343 ( .A(n294), .B(n293), .ZN(n310) );
  XOR2_X1 U344 ( .A(KEYINPUT77), .B(KEYINPUT12), .Z(n296) );
  NAND2_X1 U345 ( .A1(G231GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U346 ( .A(n296), .B(n295), .ZN(n298) );
  INV_X1 U347 ( .A(KEYINPUT15), .ZN(n297) );
  XNOR2_X1 U348 ( .A(n298), .B(n297), .ZN(n303) );
  XOR2_X1 U349 ( .A(G57GAT), .B(G155GAT), .Z(n300) );
  XNOR2_X1 U350 ( .A(G1GAT), .B(G127GAT), .ZN(n299) );
  XNOR2_X1 U351 ( .A(n300), .B(n299), .ZN(n347) );
  XNOR2_X1 U352 ( .A(G78GAT), .B(KEYINPUT13), .ZN(n301) );
  XNOR2_X1 U353 ( .A(n301), .B(KEYINPUT67), .ZN(n380) );
  XNOR2_X1 U354 ( .A(n347), .B(n380), .ZN(n302) );
  XNOR2_X1 U355 ( .A(n303), .B(n302), .ZN(n308) );
  XOR2_X1 U356 ( .A(G15GAT), .B(G22GAT), .Z(n366) );
  XOR2_X1 U357 ( .A(G8GAT), .B(G211GAT), .Z(n354) );
  XNOR2_X1 U358 ( .A(n366), .B(n354), .ZN(n306) );
  XOR2_X1 U359 ( .A(KEYINPUT14), .B(G64GAT), .Z(n305) );
  XNOR2_X1 U360 ( .A(G183GAT), .B(G71GAT), .ZN(n304) );
  XOR2_X1 U361 ( .A(n310), .B(n309), .Z(n555) );
  XNOR2_X1 U362 ( .A(n555), .B(KEYINPUT114), .ZN(n539) );
  XOR2_X1 U363 ( .A(G176GAT), .B(G183GAT), .Z(n312) );
  XNOR2_X1 U364 ( .A(G169GAT), .B(KEYINPUT82), .ZN(n311) );
  XNOR2_X1 U365 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U366 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n314) );
  XNOR2_X1 U367 ( .A(G190GAT), .B(KEYINPUT19), .ZN(n313) );
  XNOR2_X1 U368 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U369 ( .A(n316), .B(n315), .Z(n361) );
  XOR2_X1 U370 ( .A(KEYINPUT83), .B(KEYINPUT81), .Z(n318) );
  XNOR2_X1 U371 ( .A(G127GAT), .B(KEYINPUT80), .ZN(n317) );
  XNOR2_X1 U372 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U373 ( .A(n361), .B(n319), .ZN(n327) );
  XNOR2_X1 U374 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n320) );
  XNOR2_X1 U375 ( .A(n320), .B(G120GAT), .ZN(n331) );
  XOR2_X1 U376 ( .A(G43GAT), .B(G134GAT), .Z(n398) );
  XNOR2_X1 U377 ( .A(n331), .B(n398), .ZN(n322) );
  AND2_X1 U378 ( .A1(G227GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U379 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U380 ( .A(n323), .B(KEYINPUT20), .ZN(n325) );
  XOR2_X1 U381 ( .A(G99GAT), .B(G71GAT), .Z(n381) );
  XOR2_X1 U382 ( .A(G15GAT), .B(n381), .Z(n324) );
  XNOR2_X1 U383 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U384 ( .A(n327), .B(n326), .ZN(n533) );
  XOR2_X1 U385 ( .A(KEYINPUT1), .B(KEYINPUT89), .Z(n333) );
  XOR2_X1 U386 ( .A(KEYINPUT6), .B(KEYINPUT5), .Z(n329) );
  XNOR2_X1 U387 ( .A(KEYINPUT86), .B(KEYINPUT87), .ZN(n328) );
  XNOR2_X1 U388 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U390 ( .A(n333), .B(n332), .ZN(n340) );
  XOR2_X1 U391 ( .A(G29GAT), .B(G85GAT), .Z(n397) );
  XOR2_X1 U392 ( .A(KEYINPUT4), .B(KEYINPUT88), .Z(n335) );
  XNOR2_X1 U393 ( .A(G134GAT), .B(G162GAT), .ZN(n334) );
  XNOR2_X1 U394 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U395 ( .A(n397), .B(n336), .Z(n338) );
  NAND2_X1 U396 ( .A1(G225GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U397 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U398 ( .A(n340), .B(n339), .Z(n349) );
  INV_X1 U399 ( .A(KEYINPUT2), .ZN(n341) );
  NAND2_X1 U400 ( .A1(G148GAT), .A2(n341), .ZN(n344) );
  INV_X1 U401 ( .A(G148GAT), .ZN(n342) );
  NAND2_X1 U402 ( .A1(n342), .A2(KEYINPUT2), .ZN(n343) );
  NAND2_X1 U403 ( .A1(n344), .A2(n343), .ZN(n346) );
  XNOR2_X1 U404 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n345) );
  XNOR2_X1 U405 ( .A(n346), .B(n345), .ZN(n436) );
  XNOR2_X1 U406 ( .A(n436), .B(n347), .ZN(n348) );
  XNOR2_X1 U407 ( .A(n349), .B(n348), .ZN(n467) );
  XNOR2_X1 U408 ( .A(KEYINPUT91), .B(KEYINPUT93), .ZN(n351) );
  AND2_X1 U409 ( .A1(G226GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U410 ( .A(n351), .B(n350), .ZN(n353) );
  INV_X1 U411 ( .A(KEYINPUT92), .ZN(n352) );
  XNOR2_X1 U412 ( .A(n353), .B(n352), .ZN(n356) );
  XOR2_X1 U413 ( .A(G197GAT), .B(KEYINPUT21), .Z(n435) );
  XNOR2_X1 U414 ( .A(n435), .B(n354), .ZN(n355) );
  XOR2_X1 U415 ( .A(n356), .B(n355), .Z(n358) );
  XNOR2_X1 U416 ( .A(G36GAT), .B(G218GAT), .ZN(n357) );
  XNOR2_X1 U417 ( .A(n357), .B(KEYINPUT74), .ZN(n414) );
  XNOR2_X1 U418 ( .A(n358), .B(n414), .ZN(n363) );
  XOR2_X1 U419 ( .A(G64GAT), .B(KEYINPUT68), .Z(n360) );
  XNOR2_X1 U420 ( .A(G204GAT), .B(G92GAT), .ZN(n359) );
  XNOR2_X1 U421 ( .A(n360), .B(n359), .ZN(n384) );
  XNOR2_X1 U422 ( .A(n361), .B(n384), .ZN(n362) );
  XOR2_X1 U423 ( .A(KEYINPUT123), .B(n521), .Z(n431) );
  XOR2_X1 U424 ( .A(G50GAT), .B(G43GAT), .Z(n365) );
  XNOR2_X1 U425 ( .A(G29GAT), .B(G36GAT), .ZN(n364) );
  XNOR2_X1 U426 ( .A(n365), .B(n364), .ZN(n379) );
  XOR2_X1 U427 ( .A(KEYINPUT30), .B(n366), .Z(n368) );
  NAND2_X1 U428 ( .A1(G229GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U429 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U430 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n405) );
  XOR2_X1 U431 ( .A(n369), .B(n405), .Z(n377) );
  XOR2_X1 U432 ( .A(G197GAT), .B(G141GAT), .Z(n371) );
  XNOR2_X1 U433 ( .A(G169GAT), .B(G113GAT), .ZN(n370) );
  XNOR2_X1 U434 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U435 ( .A(KEYINPUT66), .B(KEYINPUT29), .Z(n373) );
  XNOR2_X1 U436 ( .A(G1GAT), .B(G8GAT), .ZN(n372) );
  XNOR2_X1 U437 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U438 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U439 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U440 ( .A(n379), .B(n378), .Z(n573) );
  INV_X1 U441 ( .A(n573), .ZN(n560) );
  XOR2_X1 U442 ( .A(n380), .B(G85GAT), .Z(n383) );
  XNOR2_X1 U443 ( .A(n381), .B(G106GAT), .ZN(n382) );
  XNOR2_X1 U444 ( .A(n383), .B(n382), .ZN(n388) );
  XOR2_X1 U445 ( .A(KEYINPUT69), .B(n384), .Z(n386) );
  NAND2_X1 U446 ( .A1(G230GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U447 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U448 ( .A(n388), .B(n387), .Z(n396) );
  XOR2_X1 U449 ( .A(G57GAT), .B(G148GAT), .Z(n390) );
  XNOR2_X1 U450 ( .A(G176GAT), .B(G120GAT), .ZN(n389) );
  XNOR2_X1 U451 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U452 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n392) );
  XNOR2_X1 U453 ( .A(KEYINPUT31), .B(KEYINPUT70), .ZN(n391) );
  XNOR2_X1 U454 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U455 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n396), .B(n395), .ZN(n577) );
  XOR2_X1 U457 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n400) );
  XNOR2_X1 U458 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U459 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U460 ( .A(KEYINPUT73), .B(G92GAT), .Z(n402) );
  NAND2_X1 U461 ( .A1(G232GAT), .A2(G233GAT), .ZN(n401) );
  XOR2_X1 U462 ( .A(n402), .B(n401), .Z(n403) );
  XNOR2_X1 U463 ( .A(n404), .B(n403), .ZN(n407) );
  XNOR2_X1 U464 ( .A(n405), .B(G190GAT), .ZN(n406) );
  XNOR2_X1 U465 ( .A(n407), .B(n406), .ZN(n411) );
  XOR2_X1 U466 ( .A(KEYINPUT9), .B(KEYINPUT64), .Z(n409) );
  XNOR2_X1 U467 ( .A(G99GAT), .B(KEYINPUT11), .ZN(n408) );
  XNOR2_X1 U468 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U469 ( .A(n411), .B(n410), .Z(n416) );
  XOR2_X1 U470 ( .A(G106GAT), .B(G162GAT), .Z(n413) );
  XNOR2_X1 U471 ( .A(G50GAT), .B(KEYINPUT72), .ZN(n412) );
  XNOR2_X1 U472 ( .A(n413), .B(n412), .ZN(n440) );
  XNOR2_X1 U473 ( .A(n440), .B(n414), .ZN(n415) );
  XNOR2_X1 U474 ( .A(n416), .B(n415), .ZN(n481) );
  XNOR2_X1 U475 ( .A(KEYINPUT36), .B(n481), .ZN(n583) );
  INV_X1 U476 ( .A(n555), .ZN(n417) );
  NOR2_X1 U477 ( .A1(n583), .A2(n417), .ZN(n419) );
  XNOR2_X1 U478 ( .A(KEYINPUT45), .B(KEYINPUT115), .ZN(n418) );
  XOR2_X1 U479 ( .A(n419), .B(n418), .Z(n420) );
  NAND2_X1 U480 ( .A1(n577), .A2(n420), .ZN(n421) );
  XNOR2_X1 U481 ( .A(n421), .B(KEYINPUT116), .ZN(n422) );
  NOR2_X1 U482 ( .A1(n560), .A2(n422), .ZN(n428) );
  XOR2_X1 U483 ( .A(n577), .B(KEYINPUT41), .Z(n536) );
  NOR2_X1 U484 ( .A1(n573), .A2(n536), .ZN(n423) );
  XNOR2_X1 U485 ( .A(n423), .B(KEYINPUT46), .ZN(n424) );
  NOR2_X1 U486 ( .A1(n539), .A2(n424), .ZN(n425) );
  NAND2_X1 U487 ( .A1(n481), .A2(n425), .ZN(n426) );
  XNOR2_X1 U488 ( .A(n426), .B(KEYINPUT47), .ZN(n427) );
  NOR2_X1 U489 ( .A1(n428), .A2(n427), .ZN(n430) );
  NAND2_X1 U490 ( .A1(n431), .A2(n547), .ZN(n433) );
  NOR2_X1 U491 ( .A1(n518), .A2(n434), .ZN(n572) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n438) );
  AND2_X1 U493 ( .A1(G228GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U495 ( .A(n439), .B(G78GAT), .Z(n442) );
  XNOR2_X1 U496 ( .A(G22GAT), .B(n440), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n442), .B(n441), .ZN(n450) );
  XOR2_X1 U498 ( .A(KEYINPUT23), .B(KEYINPUT85), .Z(n444) );
  XNOR2_X1 U499 ( .A(G218GAT), .B(KEYINPUT22), .ZN(n443) );
  XNOR2_X1 U500 ( .A(n444), .B(n443), .ZN(n448) );
  XOR2_X1 U501 ( .A(G155GAT), .B(G204GAT), .Z(n446) );
  XNOR2_X1 U502 ( .A(KEYINPUT24), .B(G211GAT), .ZN(n445) );
  XNOR2_X1 U503 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U504 ( .A(n448), .B(n447), .Z(n449) );
  XNOR2_X1 U505 ( .A(n450), .B(n449), .ZN(n456) );
  AND2_X1 U506 ( .A1(n572), .A2(n456), .ZN(n451) );
  XNOR2_X1 U507 ( .A(n451), .B(KEYINPUT55), .ZN(n452) );
  NAND2_X1 U508 ( .A1(n539), .A2(n568), .ZN(n454) );
  NAND2_X1 U509 ( .A1(n560), .A2(n577), .ZN(n455) );
  XNOR2_X1 U510 ( .A(n455), .B(KEYINPUT71), .ZN(n485) );
  INV_X1 U511 ( .A(KEYINPUT100), .ZN(n471) );
  XNOR2_X1 U512 ( .A(n521), .B(KEYINPUT27), .ZN(n463) );
  NAND2_X1 U513 ( .A1(n463), .A2(n518), .ZN(n549) );
  XOR2_X1 U514 ( .A(KEYINPUT28), .B(n456), .Z(n525) );
  XNOR2_X1 U515 ( .A(n531), .B(KEYINPUT94), .ZN(n458) );
  XNOR2_X1 U516 ( .A(n533), .B(KEYINPUT84), .ZN(n457) );
  NAND2_X1 U517 ( .A1(n458), .A2(n457), .ZN(n459) );
  XNOR2_X1 U518 ( .A(n459), .B(KEYINPUT95), .ZN(n469) );
  INV_X1 U519 ( .A(n533), .ZN(n523) );
  NAND2_X1 U520 ( .A1(n523), .A2(n521), .ZN(n460) );
  NAND2_X1 U521 ( .A1(n456), .A2(n460), .ZN(n461) );
  XNOR2_X1 U522 ( .A(n461), .B(KEYINPUT25), .ZN(n465) );
  NOR2_X1 U523 ( .A1(n523), .A2(n456), .ZN(n462) );
  XNOR2_X1 U524 ( .A(KEYINPUT26), .B(n462), .ZN(n571) );
  AND2_X1 U525 ( .A1(n463), .A2(n571), .ZN(n464) );
  NOR2_X1 U526 ( .A1(n465), .A2(n464), .ZN(n466) );
  NOR2_X1 U527 ( .A1(n467), .A2(n466), .ZN(n468) );
  NOR2_X1 U528 ( .A1(n469), .A2(n468), .ZN(n484) );
  NOR2_X1 U529 ( .A1(n555), .A2(n484), .ZN(n470) );
  XNOR2_X1 U530 ( .A(n471), .B(n470), .ZN(n472) );
  NOR2_X1 U531 ( .A1(n472), .A2(n583), .ZN(n474) );
  NAND2_X1 U532 ( .A1(n485), .A2(n517), .ZN(n476) );
  XOR2_X1 U533 ( .A(KEYINPUT103), .B(KEYINPUT38), .Z(n475) );
  XNOR2_X1 U534 ( .A(n476), .B(n475), .ZN(n477) );
  XOR2_X1 U535 ( .A(KEYINPUT102), .B(n477), .Z(n501) );
  NAND2_X1 U536 ( .A1(n501), .A2(n523), .ZN(n480) );
  XOR2_X1 U537 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n478) );
  INV_X1 U538 ( .A(n481), .ZN(n567) );
  NOR2_X1 U539 ( .A1(n567), .A2(n417), .ZN(n482) );
  XOR2_X1 U540 ( .A(KEYINPUT16), .B(n482), .Z(n483) );
  NOR2_X1 U541 ( .A1(n484), .A2(n483), .ZN(n503) );
  AND2_X1 U542 ( .A1(n485), .A2(n503), .ZN(n493) );
  NAND2_X1 U543 ( .A1(n518), .A2(n493), .ZN(n488) );
  XNOR2_X1 U544 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n486), .B(KEYINPUT96), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n488), .B(n487), .ZN(G1324GAT) );
  XOR2_X1 U547 ( .A(G8GAT), .B(KEYINPUT97), .Z(n490) );
  NAND2_X1 U548 ( .A1(n493), .A2(n521), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n490), .B(n489), .ZN(G1325GAT) );
  XOR2_X1 U550 ( .A(G15GAT), .B(KEYINPUT35), .Z(n492) );
  NAND2_X1 U551 ( .A1(n493), .A2(n523), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(G1326GAT) );
  NAND2_X1 U553 ( .A1(n525), .A2(n493), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n494), .B(KEYINPUT98), .ZN(n495) );
  XNOR2_X1 U555 ( .A(G22GAT), .B(n495), .ZN(G1327GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT99), .B(KEYINPUT104), .Z(n497) );
  XNOR2_X1 U557 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n497), .B(n496), .ZN(n499) );
  NAND2_X1 U559 ( .A1(n518), .A2(n501), .ZN(n498) );
  XOR2_X1 U560 ( .A(n499), .B(n498), .Z(G1328GAT) );
  NAND2_X1 U561 ( .A1(n501), .A2(n521), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n500), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U563 ( .A1(n525), .A2(n501), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n502), .B(G50GAT), .ZN(G1331GAT) );
  NOR2_X1 U565 ( .A1(n536), .A2(n560), .ZN(n516) );
  NAND2_X1 U566 ( .A1(n516), .A2(n503), .ZN(n504) );
  XOR2_X1 U567 ( .A(KEYINPUT106), .B(n504), .Z(n512) );
  NAND2_X1 U568 ( .A1(n512), .A2(n518), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n505), .B(KEYINPUT42), .ZN(n506) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(n506), .ZN(G1332GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n508) );
  NAND2_X1 U572 ( .A1(n512), .A2(n521), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U574 ( .A(G64GAT), .B(n509), .ZN(G1333GAT) );
  XOR2_X1 U575 ( .A(G71GAT), .B(KEYINPUT109), .Z(n511) );
  NAND2_X1 U576 ( .A1(n512), .A2(n523), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(G1334GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT43), .B(KEYINPUT110), .Z(n514) );
  NAND2_X1 U579 ( .A1(n512), .A2(n525), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U581 ( .A(G78GAT), .B(n515), .ZN(G1335GAT) );
  XOR2_X1 U582 ( .A(G85GAT), .B(KEYINPUT111), .Z(n520) );
  AND2_X1 U583 ( .A1(n517), .A2(n516), .ZN(n526) );
  NAND2_X1 U584 ( .A1(n526), .A2(n518), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(G1336GAT) );
  NAND2_X1 U586 ( .A1(n521), .A2(n526), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n522), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U588 ( .A1(n523), .A2(n526), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n524), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U590 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n530) );
  XOR2_X1 U591 ( .A(KEYINPUT113), .B(KEYINPUT112), .Z(n528) );
  NAND2_X1 U592 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n530), .B(n529), .ZN(G1339GAT) );
  NAND2_X1 U595 ( .A1(n547), .A2(n531), .ZN(n532) );
  NOR2_X1 U596 ( .A1(n533), .A2(n532), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n560), .A2(n543), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n534), .B(KEYINPUT118), .ZN(n535) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(n535), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT49), .Z(n538) );
  INV_X1 U601 ( .A(n536), .ZN(n562) );
  NAND2_X1 U602 ( .A1(n543), .A2(n562), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n541) );
  NAND2_X1 U605 ( .A1(n543), .A2(n539), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n542), .ZN(G1342GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT120), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U609 ( .A1(n543), .A2(n567), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U611 ( .A(G134GAT), .B(n546), .ZN(G1343GAT) );
  NAND2_X1 U612 ( .A1(n547), .A2(n571), .ZN(n548) );
  NOR2_X1 U613 ( .A1(n549), .A2(n548), .ZN(n557) );
  NAND2_X1 U614 ( .A1(n560), .A2(n557), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n550), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT121), .B(KEYINPUT52), .Z(n552) );
  NAND2_X1 U617 ( .A1(n557), .A2(n562), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(n554) );
  XOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT53), .Z(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  NAND2_X1 U621 ( .A1(n557), .A2(n555), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U623 ( .A1(n567), .A2(n557), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(KEYINPUT122), .ZN(n559) );
  XNOR2_X1 U625 ( .A(G162GAT), .B(n559), .ZN(G1347GAT) );
  NAND2_X1 U626 ( .A1(n560), .A2(n568), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U628 ( .A1(n568), .A2(n562), .ZN(n564) );
  XOR2_X1 U629 ( .A(G176GAT), .B(KEYINPUT125), .Z(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n566) );
  XOR2_X1 U631 ( .A(KEYINPUT57), .B(KEYINPUT56), .Z(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1349GAT) );
  XNOR2_X1 U633 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n570) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1351GAT) );
  NAND2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n582) );
  NOR2_X1 U637 ( .A1(n573), .A2(n582), .ZN(n575) );
  XNOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(n576), .ZN(G1352GAT) );
  NOR2_X1 U641 ( .A1(n577), .A2(n582), .ZN(n579) );
  XNOR2_X1 U642 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(n580) );
  XOR2_X1 U644 ( .A(G204GAT), .B(n580), .Z(G1353GAT) );
  NOR2_X1 U645 ( .A1(n417), .A2(n582), .ZN(n581) );
  XOR2_X1 U646 ( .A(G211GAT), .B(n581), .Z(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(KEYINPUT62), .B(n584), .Z(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

