//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 1 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 0 1 0 1 1 0 0 1 0 0 0 0 0 1 1 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n872, new_n873, new_n874, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G119), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT23), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G128), .ZN(new_n191));
  AND2_X1   g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G110), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(KEYINPUT71), .A3(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n189), .A2(new_n193), .A3(new_n191), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT71), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n191), .A2(new_n188), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT24), .B(G110), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n194), .A2(new_n197), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  INV_X1    g016(.A(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(G125), .A2(G140), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AND2_X1   g022(.A1(G125), .A2(G140), .ZN(new_n209));
  NOR2_X1   g023(.A1(G125), .A2(G140), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT16), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  OR3_X1    g025(.A1(new_n202), .A2(KEYINPUT16), .A3(G140), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(G146), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT72), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT72), .A4(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n201), .A2(new_n208), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n211), .A2(new_n212), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n220), .B(G146), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n198), .A2(new_n199), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n223), .B1(new_n193), .B2(new_n192), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT22), .B(G137), .ZN(new_n226));
  INV_X1    g040(.A(G221), .ZN(new_n227));
  INV_X1    g041(.A(G234), .ZN(new_n228));
  NOR3_X1   g042(.A1(new_n227), .A2(new_n228), .A3(G953), .ZN(new_n229));
  XOR2_X1   g043(.A(new_n226), .B(new_n229), .Z(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n225), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G902), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n219), .A2(new_n224), .A3(new_n230), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT25), .ZN(new_n236));
  INV_X1    g050(.A(G217), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n237), .B1(G234), .B2(new_n233), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT25), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n232), .A2(new_n239), .A3(new_n233), .A4(new_n234), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n236), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  OR2_X1    g055(.A1(new_n235), .A2(new_n238), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT32), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT67), .B1(new_n190), .B2(G116), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT67), .ZN(new_n246));
  INV_X1    g060(.A(G116), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n247), .A3(G119), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n190), .A2(G116), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  XOR2_X1   g065(.A(KEYINPUT2), .B(G113), .Z(new_n252));
  XNOR2_X1  g066(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n187), .A2(KEYINPUT1), .ZN(new_n255));
  INV_X1    g069(.A(G143), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G146), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n207), .A2(G143), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n255), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n256), .A2(KEYINPUT1), .A3(G146), .ZN(new_n260));
  XNOR2_X1  g074(.A(G143), .B(G146), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n259), .B(new_n260), .C1(G128), .C2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G134), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G137), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n263), .A2(G137), .ZN(new_n266));
  OAI21_X1  g080(.A(G131), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT11), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n268), .B1(new_n263), .B2(G137), .ZN(new_n269));
  INV_X1    g083(.A(G137), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT11), .A3(G134), .ZN(new_n271));
  INV_X1    g085(.A(G131), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n269), .A2(new_n271), .A3(new_n272), .A4(new_n264), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n262), .A2(new_n267), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(KEYINPUT0), .A2(G128), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n276), .B1(new_n261), .B2(KEYINPUT65), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n257), .A2(new_n258), .ZN(new_n278));
  XNOR2_X1  g092(.A(KEYINPUT0), .B(G128), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT65), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT66), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n277), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n282), .B1(new_n277), .B2(new_n281), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n269), .A2(new_n264), .A3(new_n271), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G131), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n273), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n275), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n254), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n277), .A2(new_n281), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT68), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n288), .A2(new_n292), .A3(KEYINPUT68), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n295), .A2(KEYINPUT30), .A3(new_n274), .A4(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT69), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n288), .A2(KEYINPUT68), .A3(new_n292), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT68), .B1(new_n288), .B2(new_n292), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n302), .A2(KEYINPUT69), .A3(KEYINPUT30), .A4(new_n274), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n291), .B1(new_n299), .B2(new_n303), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n253), .A2(new_n274), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(G237), .A2(G953), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G210), .ZN(new_n308));
  INV_X1    g122(.A(G101), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n308), .B(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n310), .B(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n306), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT31), .B1(new_n304), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT28), .ZN(new_n316));
  INV_X1    g130(.A(new_n284), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n277), .A2(new_n281), .A3(new_n282), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n288), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n274), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n254), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n316), .B1(new_n321), .B2(new_n306), .ZN(new_n322));
  AOI21_X1  g136(.A(KEYINPUT28), .B1(new_n305), .B2(new_n293), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n312), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n303), .A2(new_n299), .ZN(new_n325));
  INV_X1    g139(.A(new_n290), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n253), .B1(new_n320), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT31), .ZN(new_n329));
  INV_X1    g143(.A(new_n314), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n315), .A2(new_n324), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT70), .ZN(new_n333));
  NOR2_X1   g147(.A1(G472), .A2(G902), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n333), .B1(new_n332), .B2(new_n334), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n244), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G472), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n321), .A2(new_n306), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT28), .ZN(new_n340));
  INV_X1    g154(.A(new_n323), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n341), .A3(new_n313), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT29), .ZN(new_n343));
  INV_X1    g157(.A(new_n306), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n344), .B1(new_n325), .B2(new_n327), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n342), .B(new_n343), .C1(new_n345), .C2(new_n313), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n302), .A2(new_n274), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n254), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n306), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n323), .B1(new_n349), .B2(KEYINPUT28), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n312), .A2(new_n343), .ZN(new_n351));
  AOI21_X1  g165(.A(G902), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n338), .B1(new_n346), .B2(new_n352), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n332), .A2(new_n334), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n353), .B1(new_n354), .B2(KEYINPUT32), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n243), .B1(new_n337), .B2(new_n355), .ZN(new_n356));
  XOR2_X1   g170(.A(KEYINPUT9), .B(G234), .Z(new_n357));
  INV_X1    g171(.A(G953), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(G217), .A3(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(G128), .B(G143), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n360), .B(G134), .ZN(new_n361));
  INV_X1    g175(.A(G122), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT90), .B1(new_n362), .B2(G116), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT90), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n364), .A2(new_n247), .A3(G122), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G107), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n247), .A2(G122), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n366), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT92), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n366), .A2(KEYINPUT92), .A3(new_n367), .A4(new_n369), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n366), .A2(KEYINPUT14), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(KEYINPUT93), .A3(new_n369), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT14), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n363), .A2(new_n365), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT93), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n377), .B1(new_n363), .B2(new_n365), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n379), .B1(new_n380), .B2(new_n368), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n376), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  AOI211_X1 g196(.A(new_n361), .B(new_n374), .C1(new_n382), .C2(G107), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n360), .A2(new_n263), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(KEYINPUT91), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n263), .B1(new_n360), .B2(KEYINPUT13), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n256), .A2(G128), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n386), .B1(KEYINPUT13), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n370), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n367), .B1(new_n366), .B2(new_n369), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n385), .B(new_n388), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n359), .B1(new_n383), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n361), .B1(new_n382), .B2(G107), .ZN(new_n394));
  INV_X1    g208(.A(new_n374), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n359), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(new_n391), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n393), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n233), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT15), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n400), .A2(new_n401), .A3(G478), .ZN(new_n402));
  INV_X1    g216(.A(G478), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n399), .B(new_n233), .C1(KEYINPUT15), .C2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(G113), .B(G122), .ZN(new_n405));
  INV_X1    g219(.A(G104), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n405), .B(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT84), .ZN(new_n408));
  AOI21_X1  g222(.A(KEYINPUT85), .B1(new_n408), .B2(new_n256), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT85), .ZN(new_n410));
  OAI21_X1  g224(.A(G214), .B1(new_n410), .B2(G143), .ZN(new_n411));
  INV_X1    g225(.A(G237), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n358), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n409), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n410), .B1(KEYINPUT84), .B2(G143), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n256), .A2(KEYINPUT85), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n415), .A2(G214), .A3(new_n416), .A4(new_n307), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n272), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT17), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n414), .A2(new_n417), .A3(G131), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n414), .A2(G131), .A3(new_n417), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT17), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n422), .A2(new_n221), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(KEYINPUT18), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n209), .A2(new_n210), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G146), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n208), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT18), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n418), .B1(new_n430), .B2(new_n272), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n426), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n407), .B1(new_n425), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT89), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n425), .A2(new_n432), .A3(new_n407), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT89), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n434), .B(new_n233), .C1(new_n437), .C2(new_n433), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G475), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n402), .A2(new_n404), .A3(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(G475), .A2(G902), .ZN(new_n441));
  INV_X1    g255(.A(new_n435), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT86), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT19), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n443), .B(new_n444), .C1(new_n427), .C2(KEYINPUT87), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT87), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT86), .B1(new_n206), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(KEYINPUT86), .B1(new_n209), .B2(new_n210), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT19), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n445), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n207), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n419), .A2(new_n421), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n218), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n407), .B1(new_n453), .B2(new_n432), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n442), .A2(new_n454), .A3(KEYINPUT88), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT88), .ZN(new_n456));
  INV_X1    g270(.A(new_n407), .ZN(new_n457));
  AOI21_X1  g271(.A(G131), .B1(new_n414), .B2(new_n417), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n423), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(KEYINPUT87), .B1(new_n204), .B2(new_n205), .ZN(new_n460));
  OAI211_X1 g274(.A(KEYINPUT19), .B(new_n448), .C1(new_n460), .C2(KEYINPUT86), .ZN(new_n461));
  AOI21_X1  g275(.A(G146), .B1(new_n461), .B2(new_n445), .ZN(new_n462));
  NOR3_X1   g276(.A1(new_n459), .A2(new_n462), .A3(new_n217), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n426), .A2(new_n429), .A3(new_n431), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n457), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n456), .B1(new_n465), .B2(new_n435), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n441), .B1(new_n455), .B2(new_n466), .ZN(new_n467));
  XOR2_X1   g281(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n441), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n470), .A2(KEYINPUT20), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n471), .B1(new_n442), .B2(new_n454), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n440), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  AND2_X1   g287(.A1(new_n358), .A2(G952), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n474), .B1(new_n228), .B2(new_n412), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  OAI211_X1 g290(.A(G902), .B(G953), .C1(new_n228), .C2(new_n412), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(KEYINPUT94), .ZN(new_n478));
  XOR2_X1   g292(.A(KEYINPUT21), .B(G898), .Z(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n476), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(G214), .B1(G237), .B2(G902), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(G210), .B1(G237), .B2(G902), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n485), .B(KEYINPUT82), .Z(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n292), .A2(G125), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n262), .A2(new_n202), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT80), .B(G224), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n358), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n488), .A2(new_n492), .A3(new_n489), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT7), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(G110), .B(G122), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(KEYINPUT8), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n249), .A2(KEYINPUT5), .A3(new_n250), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n501), .B(G113), .C1(KEYINPUT5), .C2(new_n250), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n406), .A2(G107), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n367), .A2(G104), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n309), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT3), .B1(new_n406), .B2(G107), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT3), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(new_n367), .A3(G104), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n506), .A2(new_n508), .A3(new_n503), .ZN(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT76), .B(G101), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n505), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n252), .A2(new_n249), .A3(new_n250), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n502), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n512), .B1(new_n502), .B2(new_n513), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n500), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n488), .A2(new_n489), .A3(new_n496), .A4(new_n492), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n498), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT81), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n498), .A2(new_n516), .A3(KEYINPUT81), .A4(new_n517), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n502), .A2(new_n512), .A3(new_n513), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n506), .A2(new_n508), .A3(new_n503), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT4), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n524), .A3(G101), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n509), .A2(new_n309), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT4), .B1(new_n523), .B2(new_n510), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n522), .B(new_n499), .C1(new_n528), .C2(new_n253), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n520), .A2(new_n521), .A3(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n522), .B1(new_n528), .B2(new_n253), .ZN(new_n531));
  INV_X1    g345(.A(new_n499), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(KEYINPUT6), .A3(new_n529), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n494), .A2(new_n495), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT6), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n531), .A2(new_n536), .A3(new_n532), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n534), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n233), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n487), .B1(new_n530), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n520), .A2(new_n521), .A3(new_n529), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n541), .A2(new_n233), .A3(new_n485), .A4(new_n538), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n484), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n473), .A2(new_n482), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(G469), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n512), .B(new_n262), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT77), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n547), .A3(new_n288), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n548), .A2(KEYINPUT12), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT12), .ZN(new_n550));
  OR2_X1    g364(.A1(new_n512), .A2(new_n262), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n512), .A2(new_n262), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT77), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n550), .B1(new_n553), .B2(new_n288), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT10), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n292), .B(new_n525), .C1(new_n526), .C2(new_n527), .ZN(new_n557));
  INV_X1    g371(.A(new_n288), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n512), .A2(KEYINPUT10), .A3(new_n262), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n556), .A2(new_n557), .A3(new_n558), .A4(new_n559), .ZN(new_n560));
  XOR2_X1   g374(.A(G110), .B(G140), .Z(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n561), .B(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G227), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(G953), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n563), .B(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n560), .A2(new_n566), .ZN(new_n567));
  NOR3_X1   g381(.A1(new_n549), .A2(new_n554), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n556), .A2(new_n559), .A3(new_n557), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n288), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n566), .B1(new_n570), .B2(new_n560), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n545), .B(new_n233), .C1(new_n568), .C2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n548), .A2(KEYINPUT12), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n553), .A2(new_n550), .A3(new_n288), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(new_n560), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n566), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT78), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n567), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n560), .A2(KEYINPUT78), .A3(new_n566), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n570), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n577), .A2(G469), .A3(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n545), .A2(new_n233), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n572), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n227), .B1(new_n357), .B2(new_n233), .ZN(new_n586));
  XOR2_X1   g400(.A(new_n586), .B(KEYINPUT73), .Z(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(KEYINPUT79), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT79), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n585), .A2(new_n590), .A3(new_n587), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n356), .A2(new_n544), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(new_n510), .ZN(G3));
  INV_X1    g408(.A(new_n336), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n332), .A2(new_n233), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n595), .A2(new_n596), .B1(G472), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n243), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n598), .A2(new_n592), .A3(new_n599), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n383), .A2(new_n359), .A3(new_n392), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n397), .B1(new_n396), .B2(new_n391), .ZN(new_n602));
  OAI21_X1  g416(.A(KEYINPUT33), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT33), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n393), .A2(new_n604), .A3(new_n398), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n603), .A2(G478), .A3(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n403), .A2(new_n233), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n399), .A2(new_n403), .A3(new_n233), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n606), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(KEYINPUT95), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT95), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n606), .A2(new_n612), .A3(new_n608), .A4(new_n609), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  AOI22_X1  g428(.A1(new_n469), .A2(new_n472), .B1(G475), .B2(new_n438), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n485), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n617), .B1(new_n530), .B2(new_n539), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n484), .B1(new_n618), .B2(new_n542), .ZN(new_n619));
  AND4_X1   g433(.A1(new_n482), .A2(new_n614), .A3(new_n616), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n600), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT34), .B(G104), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G6));
  NAND2_X1  g437(.A1(new_n402), .A2(new_n404), .ZN(new_n624));
  INV_X1    g438(.A(new_n468), .ZN(new_n625));
  OAI21_X1  g439(.A(KEYINPUT88), .B1(new_n442), .B2(new_n454), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n465), .A2(new_n456), .A3(new_n435), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n625), .B1(new_n628), .B2(new_n441), .ZN(new_n629));
  AOI211_X1 g443(.A(new_n470), .B(new_n468), .C1(new_n626), .C2(new_n627), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT96), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n470), .B1(new_n626), .B2(new_n627), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n625), .ZN(new_n634));
  AOI21_X1  g448(.A(KEYINPUT96), .B1(new_n469), .B2(new_n634), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n624), .B(new_n439), .C1(new_n632), .C2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n619), .A2(new_n482), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n600), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT35), .B(G107), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G9));
  NOR2_X1   g455(.A1(new_n231), .A2(KEYINPUT36), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n225), .B(new_n642), .ZN(new_n643));
  OAI211_X1 g457(.A(new_n643), .B(new_n233), .C1(new_n237), .C2(G234), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n241), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n646), .B1(new_n589), .B2(new_n591), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n544), .A2(new_n598), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G110), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT97), .B(KEYINPUT37), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G12));
  NAND2_X1  g465(.A1(new_n337), .A2(new_n355), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n631), .B1(new_n629), .B2(new_n630), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n469), .A2(new_n634), .A3(KEYINPUT96), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(G900), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n476), .B1(new_n478), .B2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  AND4_X1   g472(.A1(new_n624), .A2(new_n655), .A3(new_n439), .A4(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n652), .A2(new_n659), .A3(new_n619), .A4(new_n647), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G128), .ZN(G30));
  XNOR2_X1  g475(.A(new_n657), .B(KEYINPUT39), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n592), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n646), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n666), .B1(new_n664), .B2(new_n665), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n354), .A2(KEYINPUT32), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n344), .B1(new_n254), .B2(new_n347), .ZN(new_n669));
  AOI21_X1  g483(.A(G902), .B1(new_n669), .B2(new_n312), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n670), .B1(new_n312), .B2(new_n345), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n671), .A2(KEYINPUT98), .A3(G472), .ZN(new_n672));
  AOI21_X1  g486(.A(KEYINPUT98), .B1(new_n671), .B2(G472), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n337), .A2(new_n668), .A3(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT99), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n540), .A2(new_n542), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT38), .ZN(new_n679));
  INV_X1    g493(.A(new_n624), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n615), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n667), .A2(new_n677), .A3(new_n483), .A4(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT101), .B(G143), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G45));
  OAI21_X1  g499(.A(new_n472), .B1(new_n633), .B2(new_n625), .ZN(new_n686));
  AOI221_X4 g500(.A(new_n657), .B1(new_n439), .B2(new_n686), .C1(new_n611), .C2(new_n613), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n652), .A2(new_n619), .A3(new_n647), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT102), .B(G146), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G48));
  INV_X1    g504(.A(new_n572), .ZN(new_n691));
  INV_X1    g505(.A(new_n571), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n573), .A2(new_n560), .A3(new_n574), .A4(new_n566), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n545), .B1(new_n694), .B2(new_n233), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n691), .A2(new_n695), .A3(new_n586), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n356), .A2(new_n620), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT41), .B(G113), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G15));
  NAND4_X1  g513(.A1(new_n652), .A2(new_n638), .A3(new_n599), .A4(new_n696), .ZN(new_n700));
  XOR2_X1   g514(.A(KEYINPUT103), .B(G116), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G18));
  AND3_X1   g516(.A1(new_n619), .A2(new_n696), .A3(new_n482), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n652), .A2(new_n473), .A3(new_n645), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G119), .ZN(G21));
  NAND2_X1  g519(.A1(new_n597), .A2(G472), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n315), .A2(new_n331), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n350), .A2(new_n313), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n334), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n703), .A2(new_n710), .A3(new_n599), .A4(new_n681), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G122), .ZN(G24));
  INV_X1    g526(.A(new_n619), .ZN(new_n713));
  INV_X1    g527(.A(new_n696), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n706), .A2(new_n645), .A3(new_n709), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n715), .A2(new_n687), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G125), .ZN(G27));
  INV_X1    g532(.A(new_n586), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n585), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n678), .A2(new_n484), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n356), .A2(new_n687), .A3(new_n720), .A4(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT42), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n687), .A2(new_n721), .ZN(new_n725));
  OR2_X1    g539(.A1(new_n354), .A2(KEYINPUT32), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n243), .B1(new_n726), .B2(new_n355), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n725), .A2(KEYINPUT42), .A3(new_n720), .A4(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g543(.A(KEYINPUT104), .B(G131), .Z(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G33));
  INV_X1    g545(.A(new_n659), .ZN(new_n732));
  OR2_X1    g546(.A1(new_n732), .A2(KEYINPUT105), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n356), .A2(new_n721), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n732), .A2(KEYINPUT105), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n733), .A2(new_n734), .A3(new_n720), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G134), .ZN(G36));
  NAND2_X1  g551(.A1(new_n614), .A2(new_n615), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT43), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n598), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n740), .A2(new_n741), .A3(new_n645), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n740), .A2(KEYINPUT44), .A3(new_n741), .A4(new_n645), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT46), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n577), .A2(KEYINPUT45), .A3(new_n581), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT45), .B1(new_n577), .B2(new_n581), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n747), .A2(new_n748), .A3(new_n545), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n746), .B1(new_n749), .B2(new_n583), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n691), .B1(new_n750), .B2(KEYINPUT106), .ZN(new_n751));
  OR3_X1    g565(.A1(new_n749), .A2(new_n746), .A3(new_n583), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n751), .B(new_n752), .C1(KEYINPUT106), .C2(new_n750), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n753), .A2(new_n719), .A3(new_n663), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n721), .B(KEYINPUT107), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n744), .A2(new_n745), .A3(new_n754), .A4(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G137), .ZN(G39));
  NAND4_X1  g571(.A1(new_n725), .A2(new_n243), .A3(new_n337), .A4(new_n355), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(KEYINPUT109), .ZN(new_n759));
  XOR2_X1   g573(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n760));
  AND3_X1   g574(.A1(new_n753), .A2(new_n719), .A3(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT47), .ZN(new_n762));
  AOI22_X1  g576(.A1(new_n753), .A2(new_n719), .B1(KEYINPUT108), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  XOR2_X1   g579(.A(KEYINPUT110), .B(G140), .Z(new_n766));
  XNOR2_X1  g580(.A(new_n765), .B(new_n766), .ZN(G42));
  NOR2_X1   g581(.A1(new_n691), .A2(new_n695), .ZN(new_n768));
  XOR2_X1   g582(.A(new_n768), .B(KEYINPUT49), .Z(new_n769));
  INV_X1    g583(.A(new_n587), .ZN(new_n770));
  OR4_X1    g584(.A1(new_n484), .A2(new_n769), .A3(new_n770), .A4(new_n679), .ZN(new_n771));
  OR4_X1    g585(.A1(new_n243), .A2(new_n771), .A3(new_n677), .A4(new_n738), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n710), .A2(new_n599), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n740), .A2(new_n476), .A3(new_n484), .A4(new_n773), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n679), .A2(new_n714), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(KEYINPUT50), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n714), .A2(new_n678), .A3(new_n484), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n740), .A2(new_n476), .A3(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n716), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT113), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n740), .A2(new_n476), .A3(new_n773), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n691), .A2(new_n695), .A3(new_n587), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n755), .B(new_n783), .C1(new_n764), .C2(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n677), .A2(new_n475), .ZN(new_n786));
  INV_X1    g600(.A(new_n614), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n778), .A2(new_n599), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n786), .A2(new_n615), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n777), .A2(new_n782), .A3(new_n785), .A4(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT51), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n727), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n779), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT48), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n794), .B(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n615), .B1(new_n611), .B2(new_n613), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n786), .A2(new_n797), .A3(new_n788), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n796), .A2(new_n474), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n799), .B1(new_n790), .B2(new_n791), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n792), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n645), .A2(new_n657), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n681), .A2(new_n619), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n675), .A2(new_n720), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n804), .A2(new_n660), .A3(new_n688), .A4(new_n717), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT52), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n713), .B1(new_n337), .B2(new_n355), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n807), .B(new_n647), .C1(new_n659), .C2(new_n687), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n808), .A2(new_n809), .A3(new_n717), .A4(new_n804), .ZN(new_n810));
  AND4_X1   g624(.A1(new_n697), .A2(new_n700), .A3(new_n704), .A4(new_n711), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n806), .A2(new_n729), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT112), .ZN(new_n813));
  OAI21_X1  g627(.A(KEYINPUT53), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n543), .A2(new_n482), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n598), .A2(new_n815), .A3(new_n599), .A4(new_n592), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n616), .A2(new_n680), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n648), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT111), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n648), .B(KEYINPUT111), .C1(new_n816), .C2(new_n818), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n710), .A2(new_n797), .A3(new_n720), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n652), .A2(new_n592), .A3(new_n655), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n824), .B1(new_n825), .B2(new_n440), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n826), .A2(new_n645), .A3(new_n658), .A4(new_n721), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n600), .A2(new_n815), .A3(new_n797), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n823), .A2(new_n827), .A3(new_n593), .A4(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n736), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n812), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n814), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n805), .A2(KEYINPUT52), .B1(new_n724), .B2(new_n728), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n834), .A2(KEYINPUT112), .A3(new_n810), .A4(new_n811), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n834), .A2(new_n736), .A3(new_n810), .A4(new_n811), .ZN(new_n836));
  OAI211_X1 g650(.A(KEYINPUT53), .B(new_n835), .C1(new_n836), .C2(new_n829), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT54), .B1(new_n833), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n832), .A2(new_n830), .A3(KEYINPUT53), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n841), .B1(new_n836), .B2(new_n829), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n839), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n783), .A2(new_n715), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(KEYINPUT114), .ZN(new_n845));
  NOR4_X1   g659(.A1(new_n801), .A2(new_n838), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(G952), .A2(G953), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n772), .B1(new_n846), .B2(new_n847), .ZN(G75));
  NAND2_X1  g662(.A1(new_n534), .A2(new_n537), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(KEYINPUT115), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n535), .B(KEYINPUT55), .ZN(new_n851));
  XOR2_X1   g665(.A(new_n850), .B(new_n851), .Z(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  AND4_X1   g667(.A1(G210), .A2(new_n833), .A3(G902), .A4(new_n837), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n853), .B1(new_n854), .B2(KEYINPUT56), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n358), .A2(G952), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n833), .A2(new_n837), .A3(G902), .A4(new_n487), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT116), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT56), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n852), .B1(new_n858), .B2(KEYINPUT116), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n855), .B(new_n857), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(G51));
  XNOR2_X1  g678(.A(new_n583), .B(KEYINPUT57), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n833), .A2(KEYINPUT54), .A3(new_n837), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n865), .B1(new_n866), .B2(new_n838), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n694), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n833), .A2(new_n837), .A3(G902), .A4(new_n749), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT117), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n856), .B1(new_n868), .B2(new_n870), .ZN(G54));
  NAND4_X1  g685(.A1(new_n833), .A2(new_n837), .A3(KEYINPUT58), .A4(G902), .ZN(new_n872));
  INV_X1    g686(.A(G475), .ZN(new_n873));
  INV_X1    g687(.A(new_n628), .ZN(new_n874));
  OR3_X1    g688(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n874), .B1(new_n872), .B2(new_n873), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n875), .A2(new_n857), .A3(new_n876), .ZN(G60));
  XOR2_X1   g691(.A(new_n607), .B(KEYINPUT59), .Z(new_n878));
  OAI21_X1  g692(.A(new_n878), .B1(new_n838), .B2(new_n843), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n879), .A2(new_n603), .A3(new_n605), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n603), .A2(new_n605), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n881), .B(new_n878), .C1(new_n866), .C2(new_n838), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n880), .A2(new_n857), .A3(new_n882), .ZN(G63));
  NAND2_X1  g697(.A1(G217), .A2(G902), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n884), .B(KEYINPUT60), .Z(new_n885));
  XNOR2_X1  g699(.A(new_n643), .B(KEYINPUT118), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n833), .A2(new_n837), .A3(new_n885), .A4(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n887), .A2(new_n857), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n833), .A2(new_n837), .A3(new_n885), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n232), .A2(new_n234), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT61), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n888), .B(new_n891), .C1(KEYINPUT119), .C2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n887), .A2(KEYINPUT119), .A3(new_n857), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n889), .A2(new_n890), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n887), .A2(new_n857), .ZN(new_n896));
  OAI211_X1 g710(.A(KEYINPUT61), .B(new_n894), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n893), .A2(new_n897), .ZN(G66));
  AOI21_X1  g712(.A(new_n358), .B1(new_n479), .B2(new_n491), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n823), .A2(new_n828), .A3(new_n593), .A4(new_n811), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n899), .B1(new_n900), .B2(new_n358), .ZN(new_n901));
  MUX2_X1   g715(.A(new_n899), .B(new_n901), .S(KEYINPUT120), .Z(new_n902));
  INV_X1    g716(.A(G898), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n850), .B1(new_n903), .B2(G953), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n902), .B(new_n904), .ZN(G69));
  INV_X1    g719(.A(KEYINPUT123), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n808), .A2(new_n717), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n683), .A2(new_n907), .ZN(new_n908));
  XOR2_X1   g722(.A(KEYINPUT121), .B(KEYINPUT62), .Z(new_n909));
  AOI22_X1  g723(.A1(new_n908), .A2(new_n909), .B1(new_n764), .B2(new_n759), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT62), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n683), .B(new_n907), .C1(KEYINPUT121), .C2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n664), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n734), .B(new_n913), .C1(new_n797), .C2(new_n817), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT122), .B1(new_n756), .B2(new_n914), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n756), .A2(KEYINPUT122), .A3(new_n914), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n910), .B(new_n912), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n325), .B1(new_n289), .B2(new_n290), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(new_n450), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n917), .A2(new_n358), .A3(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT125), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n754), .A2(new_n921), .A3(new_n727), .A4(new_n803), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n765), .A2(new_n729), .A3(new_n756), .A4(new_n922), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n754), .A2(new_n727), .A3(new_n803), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n736), .B(new_n907), .C1(new_n924), .C2(new_n921), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n358), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n919), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n656), .A2(G953), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT124), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n926), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n906), .B1(new_n920), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(G953), .B1(new_n564), .B2(new_n656), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(G72));
  NAND2_X1  g747(.A1(G472), .A2(G902), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT63), .Z(new_n935));
  OAI21_X1  g749(.A(new_n935), .B1(new_n917), .B2(new_n900), .ZN(new_n936));
  INV_X1    g750(.A(new_n345), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n313), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n856), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n923), .A2(new_n925), .A3(new_n900), .ZN(new_n941));
  INV_X1    g755(.A(new_n935), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n312), .B(new_n345), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n840), .A2(new_n842), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n328), .A2(new_n330), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n937), .A2(new_n312), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT126), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n944), .B(new_n935), .C1(new_n946), .C2(new_n948), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n940), .A2(new_n943), .A3(new_n949), .ZN(G57));
endmodule


