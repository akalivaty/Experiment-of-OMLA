//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 0 1 1 1 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n812, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT69), .ZN(new_n188));
  OR2_X1    g002(.A1(KEYINPUT64), .A2(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT64), .A2(G146), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(G143), .A3(new_n190), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT0), .A2(G128), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  AND3_X1   g009(.A1(new_n191), .A2(new_n192), .A3(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G128), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  AND2_X1   g012(.A1(KEYINPUT64), .A2(G146), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT64), .A2(G146), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n198), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n193), .A2(G143), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n197), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n188), .B1(new_n196), .B2(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n191), .A2(new_n192), .A3(new_n195), .ZN(new_n205));
  INV_X1    g019(.A(new_n202), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n189), .A2(new_n190), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(new_n198), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n205), .B(KEYINPUT69), .C1(new_n208), .C2(new_n197), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n204), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT11), .ZN(new_n211));
  INV_X1    g025(.A(G134), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n211), .B1(new_n212), .B2(G137), .ZN(new_n213));
  INV_X1    g027(.A(G137), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(KEYINPUT11), .A3(G134), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n212), .A2(G137), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n213), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT65), .B(G131), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n217), .A2(new_n218), .A3(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n213), .A2(new_n215), .A3(new_n216), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT66), .B1(new_n222), .B2(new_n219), .ZN(new_n223));
  AOI22_X1  g037(.A1(new_n221), .A2(new_n223), .B1(G131), .B2(new_n222), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n187), .B1(new_n210), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n214), .A2(G134), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n216), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n221), .A2(new_n223), .B1(G131), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G128), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n191), .A2(new_n195), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n229), .B1(new_n191), .B2(KEYINPUT1), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(new_n208), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT2), .ZN(new_n234));
  INV_X1    g048(.A(G113), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT67), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(KEYINPUT2), .A3(G113), .ZN(new_n238));
  AOI22_X1  g052(.A1(new_n236), .A2(new_n238), .B1(new_n234), .B2(new_n235), .ZN(new_n239));
  XNOR2_X1  g053(.A(G116), .B(G119), .ZN(new_n240));
  AOI21_X1  g054(.A(KEYINPUT68), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n236), .A2(new_n238), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n234), .A2(new_n235), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n240), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n244), .A2(KEYINPUT68), .A3(new_n245), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n228), .A2(new_n233), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n222), .A2(G131), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n218), .B1(new_n217), .B2(new_n220), .ZN(new_n251));
  NOR3_X1   g065(.A1(new_n222), .A2(KEYINPUT66), .A3(new_n219), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n253), .A2(KEYINPUT70), .A3(new_n204), .A4(new_n209), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n225), .A2(new_n249), .A3(new_n254), .ZN(new_n255));
  XOR2_X1   g069(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n256));
  NOR2_X1   g070(.A1(G237), .A2(G953), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G210), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n256), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT26), .B(G101), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n259), .B(new_n260), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n261), .A2(KEYINPUT72), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n255), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n263), .A2(KEYINPUT31), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n247), .A2(new_n248), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n221), .A2(new_n223), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n227), .A2(G131), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(new_n233), .A3(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n205), .B1(new_n208), .B2(new_n197), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n268), .B1(new_n224), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n270), .A2(KEYINPUT30), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n225), .A2(new_n268), .A3(new_n254), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n271), .B1(KEYINPUT30), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n264), .B1(new_n265), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT28), .ZN(new_n275));
  INV_X1    g089(.A(new_n265), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n275), .B1(new_n255), .B2(new_n277), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n265), .B(new_n268), .C1(new_n210), .C2(new_n224), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n275), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n261), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n272), .A2(KEYINPUT30), .ZN(new_n283));
  INV_X1    g097(.A(new_n271), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n263), .B1(new_n285), .B2(new_n276), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT31), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n274), .B(new_n282), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(G472), .A2(G902), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(KEYINPUT32), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT74), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n288), .A2(new_n289), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT32), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n255), .A2(new_n277), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n281), .B1(new_n296), .B2(KEYINPUT28), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT29), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n261), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n272), .A2(new_n276), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n275), .B1(new_n300), .B2(new_n255), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT73), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n280), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n279), .A2(KEYINPUT73), .A3(new_n275), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT29), .B1(new_n301), .B2(new_n305), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n299), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G902), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n255), .B(new_n261), .C1(new_n273), .C2(new_n265), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n308), .B1(new_n309), .B2(KEYINPUT29), .ZN(new_n310));
  OAI21_X1  g124(.A(G472), .B1(new_n307), .B2(new_n310), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n288), .A2(KEYINPUT74), .A3(KEYINPUT32), .A4(new_n289), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n292), .A2(new_n295), .A3(new_n311), .A4(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT25), .ZN(new_n314));
  INV_X1    g128(.A(G140), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G125), .ZN(new_n316));
  INV_X1    g130(.A(G125), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G140), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n316), .A2(new_n318), .A3(KEYINPUT16), .ZN(new_n319));
  OR3_X1    g133(.A1(new_n317), .A2(KEYINPUT16), .A3(G140), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n193), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n319), .A2(new_n320), .A3(G146), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G119), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(KEYINPUT76), .A3(G128), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n229), .A2(G119), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(KEYINPUT76), .B1(new_n325), .B2(G128), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  XOR2_X1   g144(.A(KEYINPUT24), .B(G110), .Z(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n325), .A2(G128), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n229), .A2(KEYINPUT23), .A3(G119), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n325), .A2(G128), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n333), .B(new_n334), .C1(new_n335), .C2(KEYINPUT23), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G110), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n324), .A2(new_n332), .A3(new_n337), .ZN(new_n338));
  OAI22_X1  g152(.A1(new_n330), .A2(new_n331), .B1(new_n336), .B2(G110), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT77), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n323), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n319), .A2(new_n320), .A3(KEYINPUT77), .A4(G146), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n316), .A2(new_n318), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n199), .A2(new_n200), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n339), .A2(new_n341), .A3(new_n342), .A4(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT22), .B(G137), .ZN(new_n347));
  INV_X1    g161(.A(G953), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(G221), .A3(G234), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n347), .B(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n338), .A2(new_n346), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n350), .B1(new_n338), .B2(new_n346), .ZN(new_n353));
  NOR3_X1   g167(.A1(new_n352), .A2(new_n353), .A3(G902), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n314), .B1(new_n354), .B2(KEYINPUT78), .ZN(new_n355));
  INV_X1    g169(.A(new_n353), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(new_n308), .A3(new_n351), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT78), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n358), .A3(KEYINPUT25), .ZN(new_n359));
  XNOR2_X1  g173(.A(KEYINPUT75), .B(G217), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n361), .B1(G234), .B2(new_n308), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n355), .A2(new_n359), .A3(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n352), .A2(new_n353), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n362), .A2(G902), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n313), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G469), .ZN(new_n370));
  XNOR2_X1  g184(.A(G110), .B(G140), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n348), .A2(G227), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n371), .B(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT4), .ZN(new_n374));
  INV_X1    g188(.A(G107), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G104), .ZN(new_n376));
  OR2_X1    g190(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n377));
  NAND2_X1  g191(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G104), .ZN(new_n380));
  OAI22_X1  g194(.A1(new_n380), .A2(G107), .B1(KEYINPUT80), .B2(KEYINPUT3), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(G107), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(G101), .B1(new_n379), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n380), .A2(G107), .ZN(new_n385));
  INV_X1    g199(.A(new_n378), .ZN(new_n386));
  NOR2_X1   g200(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AND2_X1   g202(.A1(KEYINPUT81), .A2(G101), .ZN(new_n389));
  NOR2_X1   g203(.A1(KEYINPUT81), .A2(G101), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n388), .A2(new_n391), .A3(new_n382), .A4(new_n381), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n374), .B1(new_n384), .B2(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n375), .A2(G104), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n394), .B1(new_n376), .B2(new_n377), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n388), .ZN(new_n396));
  AOI21_X1  g210(.A(KEYINPUT4), .B1(new_n396), .B2(G101), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n199), .A2(new_n200), .A3(new_n198), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT1), .ZN(new_n400));
  OAI21_X1  g214(.A(G128), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n201), .A2(new_n202), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n194), .B1(new_n344), .B2(G143), .ZN(new_n403));
  AOI22_X1  g217(.A1(new_n401), .A2(new_n402), .B1(new_n403), .B2(new_n230), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT82), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n376), .A2(new_n382), .A3(new_n405), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n406), .B(G101), .C1(new_n405), .C2(new_n376), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n392), .A2(new_n407), .A3(KEYINPUT10), .ZN(new_n408));
  OAI22_X1  g222(.A1(new_n398), .A2(new_n210), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT85), .ZN(new_n410));
  OAI211_X1 g224(.A(KEYINPUT84), .B(KEYINPUT1), .C1(new_n198), .C2(G146), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G128), .ZN(new_n412));
  AOI21_X1  g226(.A(KEYINPUT84), .B1(new_n202), .B2(KEYINPUT1), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n410), .B1(new_n414), .B2(new_n403), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT1), .B1(new_n198), .B2(G146), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT84), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(G128), .A3(new_n411), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n191), .A2(new_n195), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(KEYINPUT85), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT83), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n231), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n191), .A2(KEYINPUT83), .A3(new_n195), .A4(new_n230), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n415), .A2(new_n421), .A3(new_n423), .A4(new_n424), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n392), .A2(new_n407), .ZN(new_n426));
  AOI21_X1  g240(.A(KEYINPUT10), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n409), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n373), .B1(new_n428), .B2(new_n224), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n404), .A2(new_n408), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n204), .A2(new_n209), .ZN(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT81), .B(G101), .ZN(new_n432));
  NOR3_X1   g246(.A1(new_n379), .A2(new_n383), .A3(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(G101), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n434), .B1(new_n395), .B2(new_n388), .ZN(new_n435));
  OAI21_X1  g249(.A(KEYINPUT4), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n384), .A2(new_n374), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n430), .B1(new_n431), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n421), .A2(new_n423), .A3(new_n424), .ZN(new_n440));
  AOI21_X1  g254(.A(KEYINPUT85), .B1(new_n419), .B2(new_n420), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n426), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT10), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n224), .B1(new_n439), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n429), .A2(new_n446), .ZN(new_n447));
  NOR3_X1   g261(.A1(new_n409), .A2(new_n427), .A3(new_n253), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n392), .A2(new_n407), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n404), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n442), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT12), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT86), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n452), .B1(new_n224), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(new_n253), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(KEYINPUT12), .B1(new_n253), .B2(KEYINPUT86), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n426), .A2(new_n233), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n457), .B1(new_n425), .B2(new_n426), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n456), .B1(new_n458), .B2(new_n224), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n448), .B1(new_n455), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n373), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n447), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n370), .B1(new_n462), .B2(new_n308), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n439), .A2(new_n444), .A3(new_n224), .ZN(new_n464));
  NOR3_X1   g278(.A1(new_n458), .A2(new_n224), .A3(new_n456), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n454), .B1(new_n451), .B2(new_n253), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n464), .B(new_n461), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n373), .B1(new_n448), .B2(new_n445), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(new_n370), .A3(new_n308), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT87), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(G902), .B1(new_n467), .B2(new_n468), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(KEYINPUT87), .A3(new_n370), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n463), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(G116), .B(G122), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n375), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n198), .A2(G128), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n229), .A2(G143), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n212), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n480), .A2(new_n212), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n477), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G116), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(G122), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT14), .ZN(new_n487));
  OAI21_X1  g301(.A(G107), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n488), .B1(new_n487), .B2(new_n476), .ZN(new_n489));
  OR2_X1    g303(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT9), .B(G234), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n361), .A2(G953), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT13), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT95), .B1(new_n478), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT95), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n495), .A2(new_n198), .A3(KEYINPUT13), .A4(G128), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n478), .A2(new_n493), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n494), .A2(new_n479), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G134), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT96), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n498), .A2(KEYINPUT96), .A3(G134), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(G122), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G116), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n486), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(G107), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT94), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n477), .A3(new_n508), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n486), .A2(new_n505), .A3(new_n375), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n375), .B1(new_n486), .B2(new_n505), .ZN(new_n511));
  OAI21_X1  g325(.A(KEYINPUT94), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(new_n512), .A3(new_n481), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n490), .B(new_n492), .C1(new_n503), .C2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n492), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n513), .B1(new_n501), .B2(new_n502), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n484), .A2(new_n489), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(G902), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(G478), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n520), .A2(KEYINPUT15), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  AOI211_X1 g337(.A(G902), .B(new_n521), .C1(new_n514), .C2(new_n518), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(G234), .A2(G237), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n527), .A2(G952), .A3(new_n348), .ZN(new_n528));
  XOR2_X1   g342(.A(KEYINPUT21), .B(G898), .Z(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(KEYINPUT97), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n527), .A2(G902), .A3(G953), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n526), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G475), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n345), .B1(new_n193), .B2(new_n343), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n257), .A2(G214), .ZN(new_n537));
  OR2_X1    g351(.A1(KEYINPUT91), .A2(G143), .ZN(new_n538));
  NAND2_X1  g352(.A1(KEYINPUT91), .A2(G143), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  AND2_X1   g355(.A1(KEYINPUT18), .A2(G131), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n257), .A2(G214), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n539), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n541), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n542), .B1(new_n541), .B2(new_n544), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n536), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n541), .A2(new_n220), .A3(new_n544), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n220), .B1(new_n541), .B2(new_n544), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n548), .A2(new_n549), .A3(KEYINPUT17), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n543), .B1(new_n538), .B2(new_n539), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n543), .A2(new_n539), .ZN(new_n552));
  OAI211_X1 g366(.A(KEYINPUT17), .B(new_n219), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(new_n323), .A3(new_n322), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n547), .B1(new_n550), .B2(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(G113), .B(G122), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(new_n380), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n557), .B(new_n547), .C1(new_n550), .C2(new_n554), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n535), .B1(new_n561), .B2(new_n308), .ZN(new_n562));
  NOR2_X1   g376(.A1(G475), .A2(G902), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT19), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n316), .B(new_n318), .C1(KEYINPUT92), .C2(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n565), .B(new_n344), .C1(new_n343), .C2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT93), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n566), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n316), .A2(new_n318), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n572), .A2(KEYINPUT93), .A3(new_n344), .A4(new_n565), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n341), .A2(new_n342), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n574), .B(new_n575), .C1(new_n549), .C2(new_n548), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n557), .B1(new_n576), .B2(new_n547), .ZN(new_n577));
  INV_X1    g391(.A(new_n560), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n563), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT20), .ZN(new_n580));
  INV_X1    g394(.A(new_n574), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n341), .B(new_n342), .C1(new_n548), .C2(new_n549), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n547), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n558), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n560), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT20), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n586), .A3(new_n563), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n562), .B1(new_n580), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n534), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT5), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n590), .A2(new_n325), .A3(G116), .ZN(new_n591));
  OAI211_X1 g405(.A(G113), .B(new_n591), .C1(new_n245), .C2(new_n590), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n239), .A2(new_n240), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n592), .A2(new_n593), .A3(new_n392), .A4(new_n407), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n594), .B1(new_n398), .B2(new_n265), .ZN(new_n595));
  XOR2_X1   g409(.A(G110), .B(G122), .Z(new_n596));
  INV_X1    g410(.A(KEYINPUT88), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(G110), .B(G122), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(KEYINPUT88), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n595), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n601), .B(new_n594), .C1(new_n398), .C2(new_n265), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n603), .A2(KEYINPUT6), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT6), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n595), .A2(new_n606), .A3(new_n602), .ZN(new_n607));
  OR2_X1    g421(.A1(new_n269), .A2(new_n317), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n233), .A2(new_n317), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(G224), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(G953), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n610), .B(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n605), .A2(new_n607), .A3(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT7), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n612), .B1(KEYINPUT89), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n617), .B1(KEYINPUT89), .B2(new_n616), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n608), .A2(new_n609), .A3(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT90), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n616), .B1(new_n612), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n621), .B1(new_n620), .B2(new_n612), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n608), .B2(new_n609), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT8), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n601), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n598), .A2(KEYINPUT8), .A3(new_n600), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n592), .A2(new_n593), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n449), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n627), .B1(new_n629), .B2(new_n594), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n619), .A2(new_n623), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(G902), .B1(new_n631), .B2(new_n604), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n615), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(G210), .B1(G237), .B2(G902), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n615), .A2(new_n632), .A3(new_n634), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(G214), .B1(G237), .B2(G902), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(G221), .B1(new_n491), .B2(G902), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT79), .ZN(new_n642));
  NOR4_X1   g456(.A1(new_n475), .A2(new_n589), .A3(new_n640), .A4(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n369), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(new_n432), .ZN(G3));
  NOR3_X1   g459(.A1(new_n475), .A2(new_n367), .A3(new_n642), .ZN(new_n646));
  INV_X1    g460(.A(new_n293), .ZN(new_n647));
  INV_X1    g461(.A(G472), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(new_n288), .B2(new_n308), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n533), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n638), .A2(new_n652), .A3(new_n639), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n519), .A2(new_n520), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n520), .A2(new_n308), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n514), .A2(new_n518), .ZN(new_n658));
  OAI21_X1  g472(.A(KEYINPUT33), .B1(new_n492), .B2(KEYINPUT98), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n659), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n514), .A2(new_n518), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n520), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n657), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n580), .A2(new_n587), .ZN(new_n665));
  INV_X1    g479(.A(new_n562), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT99), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(KEYINPUT99), .B1(new_n664), .B2(new_n667), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n651), .A2(new_n653), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(new_n380), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT100), .B(KEYINPUT34), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G6));
  INV_X1    g490(.A(new_n653), .ZN(new_n677));
  INV_X1    g491(.A(new_n587), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n562), .B1(new_n678), .B2(KEYINPUT101), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT101), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n580), .A2(new_n587), .A3(new_n680), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n679), .A2(new_n526), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n651), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(new_n375), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT102), .B(KEYINPUT35), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G9));
  NOR3_X1   g501(.A1(new_n475), .A2(new_n642), .A3(new_n640), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n338), .A2(new_n346), .ZN(new_n689));
  INV_X1    g503(.A(new_n350), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n690), .A2(KEYINPUT36), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n689), .B(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n365), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n363), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n534), .A2(new_n588), .A3(new_n694), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n695), .A2(new_n647), .A3(new_n649), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n688), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT37), .B(G110), .Z(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G12));
  NOR2_X1   g513(.A1(new_n475), .A2(new_n642), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n313), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(G900), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n528), .B1(new_n532), .B2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n682), .A2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n694), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n705), .A2(new_n640), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n701), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G128), .ZN(G30));
  XOR2_X1   g523(.A(new_n703), .B(KEYINPUT39), .Z(new_n710));
  NAND2_X1  g524(.A1(new_n700), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g525(.A(new_n711), .B(KEYINPUT40), .Z(new_n712));
  INV_X1    g526(.A(new_n261), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n273), .A2(new_n265), .ZN(new_n714));
  INV_X1    g528(.A(new_n255), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n715), .B1(new_n276), .B2(new_n272), .ZN(new_n717));
  AOI21_X1  g531(.A(G902), .B1(new_n717), .B2(new_n261), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n648), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n719), .B1(new_n293), .B2(new_n294), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n292), .A3(new_n312), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n638), .B(KEYINPUT38), .ZN(new_n722));
  INV_X1    g536(.A(new_n639), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n588), .A2(new_n525), .A3(new_n723), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n722), .A2(new_n706), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n712), .A2(new_n721), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G143), .ZN(G45));
  NAND3_X1  g541(.A1(new_n664), .A2(new_n667), .A3(new_n704), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n640), .A2(new_n706), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n701), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G146), .ZN(G48));
  NAND2_X1  g545(.A1(new_n313), .A2(new_n368), .ZN(new_n732));
  INV_X1    g546(.A(new_n641), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n473), .A2(new_n370), .ZN(new_n734));
  AOI211_X1 g548(.A(new_n733), .B(new_n734), .C1(new_n472), .C2(new_n474), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n668), .B(new_n669), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(new_n736), .A3(new_n677), .ZN(new_n737));
  OAI21_X1  g551(.A(KEYINPUT103), .B1(new_n732), .B2(new_n737), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n473), .A2(new_n370), .ZN(new_n739));
  AND4_X1   g553(.A1(KEYINPUT87), .A2(new_n469), .A3(new_n370), .A4(new_n308), .ZN(new_n740));
  AOI21_X1  g554(.A(KEYINPUT87), .B1(new_n473), .B2(new_n370), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n641), .B(new_n739), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n672), .A2(new_n742), .A3(new_n653), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT103), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n743), .A2(new_n744), .A3(new_n313), .A4(new_n368), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n738), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(KEYINPUT41), .B(G113), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G15));
  NOR2_X1   g562(.A1(new_n683), .A2(new_n742), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n369), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G116), .ZN(G18));
  NOR3_X1   g565(.A1(new_n742), .A2(new_n640), .A3(new_n695), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n313), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G119), .ZN(G21));
  INV_X1    g568(.A(KEYINPUT104), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n367), .B(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n289), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n255), .B(new_n262), .C1(new_n273), .C2(new_n265), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n285), .A2(new_n276), .ZN(new_n759));
  AOI22_X1  g573(.A1(new_n758), .A2(KEYINPUT31), .B1(new_n759), .B2(new_n264), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n261), .B1(new_n301), .B2(new_n305), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n757), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n756), .A2(new_n649), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n588), .A2(new_n525), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n763), .A2(new_n735), .A3(new_n677), .A4(new_n764), .ZN(new_n765));
  XOR2_X1   g579(.A(KEYINPUT105), .B(G122), .Z(new_n766));
  XNOR2_X1  g580(.A(new_n765), .B(new_n766), .ZN(G24));
  NOR3_X1   g581(.A1(new_n742), .A2(new_n640), .A3(new_n728), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n761), .B(new_n274), .C1(new_n287), .C2(new_n286), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n289), .ZN(new_n770));
  AOI21_X1  g584(.A(G902), .B1(new_n760), .B2(new_n282), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n770), .B(new_n694), .C1(new_n771), .C2(new_n648), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n768), .A2(KEYINPUT106), .A3(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT106), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n734), .B1(new_n472), .B2(new_n474), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n615), .A2(new_n632), .A3(new_n634), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n634), .B1(new_n615), .B2(new_n632), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n723), .ZN(new_n780));
  INV_X1    g594(.A(new_n728), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n776), .A2(new_n641), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n775), .B1(new_n782), .B2(new_n772), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n774), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G125), .ZN(G27));
  AND2_X1   g599(.A1(new_n295), .A2(new_n311), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n756), .B1(new_n786), .B2(new_n290), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n788));
  AOI22_X1  g602(.A1(new_n788), .A2(new_n373), .B1(new_n429), .B2(new_n446), .ZN(new_n789));
  OAI21_X1  g603(.A(G469), .B1(new_n789), .B2(G902), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n790), .B1(new_n740), .B2(new_n741), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n641), .ZN(new_n792));
  OAI21_X1  g606(.A(KEYINPUT107), .B1(new_n638), .B2(new_n723), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT107), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n779), .A2(new_n794), .A3(new_n639), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n792), .A2(new_n796), .A3(KEYINPUT108), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT108), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n472), .A2(new_n474), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n733), .B1(new_n799), .B2(new_n790), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n794), .B1(new_n779), .B2(new_n639), .ZN(new_n801));
  NOR4_X1   g615(.A1(new_n777), .A2(new_n778), .A3(KEYINPUT107), .A4(new_n723), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n798), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n781), .B(new_n787), .C1(new_n797), .C2(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(KEYINPUT108), .B1(new_n792), .B2(new_n796), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n800), .A2(new_n803), .A3(new_n798), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n732), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n728), .A2(KEYINPUT42), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n805), .A2(KEYINPUT42), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G131), .ZN(G33));
  INV_X1    g625(.A(new_n705), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n369), .B(new_n812), .C1(new_n797), .C2(new_n804), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G134), .ZN(G36));
  NOR3_X1   g628(.A1(new_n667), .A2(new_n663), .A3(new_n657), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT43), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n816), .B(new_n694), .C1(new_n647), .C2(new_n649), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT44), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n796), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n819), .B1(new_n818), .B2(new_n817), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n820), .A2(KEYINPUT110), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n789), .A2(KEYINPUT45), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n789), .A2(KEYINPUT45), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n822), .A2(G469), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(G469), .A2(G902), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n824), .A2(KEYINPUT46), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT109), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n826), .A2(new_n827), .A3(new_n799), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n827), .B1(new_n826), .B2(new_n799), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT46), .B1(new_n824), .B2(new_n825), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n831), .A2(new_n733), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n832), .A2(new_n710), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n820), .A2(KEYINPUT110), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n821), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(G137), .ZN(G39));
  NOR4_X1   g650(.A1(new_n313), .A2(new_n368), .A3(new_n796), .A4(new_n728), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n832), .A2(KEYINPUT47), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n832), .A2(KEYINPUT47), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n837), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(G140), .ZN(G42));
  INV_X1    g656(.A(new_n642), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n815), .A2(new_n843), .A3(new_n639), .ZN(new_n844));
  INV_X1    g658(.A(new_n776), .ZN(new_n845));
  AOI211_X1 g659(.A(new_n756), .B(new_n844), .C1(new_n845), .C2(KEYINPUT49), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT111), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n845), .A2(KEYINPUT49), .ZN(new_n848));
  XOR2_X1   g662(.A(new_n848), .B(KEYINPUT112), .Z(new_n849));
  OR4_X1    g663(.A1(new_n721), .A2(new_n847), .A3(new_n722), .A4(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n525), .A2(KEYINPUT113), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT113), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n853), .B1(new_n523), .B2(new_n524), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n588), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n668), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n646), .A2(new_n650), .A3(new_n677), .A4(new_n857), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n858), .A2(new_n765), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n753), .A2(new_n697), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n369), .B1(new_n643), .B2(new_n749), .ZN(new_n861));
  AND4_X1   g675(.A1(new_n746), .A2(new_n859), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n781), .B(new_n773), .C1(new_n797), .C2(new_n804), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n679), .A2(new_n681), .A3(new_n704), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n852), .A2(new_n694), .A3(new_n854), .ZN(new_n865));
  NOR4_X1   g679(.A1(new_n801), .A2(new_n802), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n866), .A2(new_n313), .A3(new_n700), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n813), .A2(new_n863), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n862), .A2(new_n810), .A3(new_n869), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n313), .B(new_n700), .C1(new_n707), .C2(new_n729), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT106), .B1(new_n768), .B2(new_n773), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n782), .A2(new_n775), .A3(new_n772), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n363), .A2(new_n693), .A3(new_n704), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n724), .A2(new_n638), .A3(new_n875), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n475), .A2(new_n733), .A3(new_n876), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n877), .A2(KEYINPUT115), .A3(new_n721), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT115), .B1(new_n877), .B2(new_n721), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT52), .B1(new_n874), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n877), .A2(new_n721), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT115), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n877), .A2(KEYINPUT115), .A3(new_n721), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT52), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n886), .A2(new_n887), .A3(new_n784), .A4(new_n871), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n881), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n851), .B1(new_n870), .B2(new_n889), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n881), .A2(new_n888), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n813), .A2(new_n863), .A3(new_n868), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT42), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n728), .B1(new_n806), .B2(new_n807), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n893), .B1(new_n894), .B2(new_n787), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n806), .A2(new_n807), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n896), .A2(new_n369), .A3(new_n809), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n892), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n891), .A2(KEYINPUT53), .A3(new_n862), .A4(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT54), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n890), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT116), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n867), .B1(new_n808), .B2(new_n812), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n805), .A2(KEYINPUT42), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n808), .A2(new_n809), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n904), .A2(new_n905), .A3(new_n906), .A4(new_n863), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n746), .A2(new_n859), .A3(new_n860), .A4(new_n861), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n909), .A2(KEYINPUT116), .A3(KEYINPUT53), .A4(new_n891), .ZN(new_n910));
  OAI21_X1  g724(.A(KEYINPUT114), .B1(new_n907), .B2(new_n908), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT114), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n862), .A2(new_n912), .A3(new_n810), .A4(new_n869), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n911), .A2(new_n913), .A3(new_n891), .ZN(new_n914));
  AOI22_X1  g728(.A1(new_n903), .A2(new_n910), .B1(new_n851), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n901), .B1(new_n915), .B2(new_n900), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT117), .ZN(new_n917));
  INV_X1    g731(.A(new_n840), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n918), .B(new_n838), .C1(new_n843), .C2(new_n845), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n816), .A2(new_n528), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n920), .A2(new_n763), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n919), .A2(new_n803), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n796), .A2(new_n742), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n920), .A2(new_n773), .A3(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n721), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n925), .A2(new_n923), .A3(new_n368), .A4(new_n528), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n926), .A2(new_n667), .A3(new_n664), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n722), .A2(new_n742), .A3(new_n639), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n928), .A2(KEYINPUT118), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(KEYINPUT118), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n921), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT50), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  AOI211_X1 g748(.A(new_n924), .B(new_n927), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n917), .B1(new_n922), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT51), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n920), .A2(new_n787), .A3(new_n923), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT48), .Z(new_n940));
  NOR2_X1   g754(.A1(new_n926), .A2(new_n672), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n742), .A2(new_n640), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n921), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n943), .A2(G952), .A3(new_n348), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n940), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n945), .B1(new_n936), .B2(new_n937), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n916), .A2(new_n938), .A3(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(G952), .A2(G953), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n850), .B1(new_n947), .B2(new_n948), .ZN(G75));
  NOR2_X1   g763(.A1(new_n348), .A2(G952), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n308), .B1(new_n890), .B2(new_n899), .ZN(new_n952));
  AOI21_X1  g766(.A(KEYINPUT56), .B1(new_n952), .B2(G210), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n605), .A2(new_n607), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(new_n614), .Z(new_n955));
  XNOR2_X1  g769(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n951), .B1(new_n953), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n959), .B1(new_n953), .B2(new_n958), .ZN(G51));
  NAND2_X1  g774(.A1(new_n890), .A2(new_n899), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(KEYINPUT54), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n901), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n825), .B(KEYINPUT57), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n469), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n952), .A2(G469), .A3(new_n823), .A4(new_n822), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n950), .B1(new_n966), .B2(new_n967), .ZN(G54));
  NAND2_X1  g782(.A1(KEYINPUT58), .A2(G475), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n585), .B1(new_n952), .B2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT120), .ZN(new_n972));
  OR2_X1    g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n971), .A2(new_n972), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n952), .A2(new_n585), .A3(new_n970), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n975), .A2(new_n951), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n973), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(KEYINPUT121), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT121), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n973), .A2(new_n979), .A3(new_n974), .A4(new_n976), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n980), .ZN(G60));
  AND2_X1   g795(.A1(new_n660), .A2(new_n662), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n655), .B(KEYINPUT59), .Z(new_n983));
  AND2_X1   g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n950), .B1(new_n963), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n982), .B1(new_n916), .B2(new_n983), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n985), .B1(new_n986), .B2(KEYINPUT122), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT122), .ZN(new_n988));
  AOI211_X1 g802(.A(new_n988), .B(new_n982), .C1(new_n916), .C2(new_n983), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n987), .A2(new_n989), .ZN(G63));
  INV_X1    g804(.A(KEYINPUT61), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n950), .B1(KEYINPUT124), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(G217), .A2(G902), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT123), .Z(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT60), .Z(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n996), .B1(new_n890), .B2(new_n899), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n992), .B1(new_n997), .B2(new_n364), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT125), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n997), .A2(new_n692), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1001), .ZN(new_n1003));
  OAI21_X1  g817(.A(KEYINPUT125), .B1(new_n1003), .B2(new_n998), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n991), .A2(KEYINPUT124), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1002), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(G66));
  XNOR2_X1  g824(.A(new_n908), .B(KEYINPUT126), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(new_n348), .ZN(new_n1012));
  OAI21_X1  g826(.A(G953), .B1(new_n531), .B2(new_n611), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n954), .B1(G898), .B2(new_n348), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n1014), .B(new_n1015), .ZN(G69));
  AOI21_X1  g830(.A(new_n348), .B1(G227), .B2(G900), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n833), .A2(new_n638), .A3(new_n724), .A4(new_n787), .ZN(new_n1018));
  INV_X1    g832(.A(new_n874), .ZN(new_n1019));
  AND3_X1   g833(.A1(new_n810), .A2(new_n813), .A3(new_n1019), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n841), .A2(new_n835), .A3(new_n1018), .A4(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n572), .A2(new_n565), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n273), .B(new_n1022), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1021), .A2(new_n348), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n726), .A2(new_n1019), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT62), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  XOR2_X1   g841(.A(new_n857), .B(KEYINPUT127), .Z(new_n1028));
  OR4_X1    g842(.A1(new_n732), .A2(new_n1028), .A3(new_n711), .A4(new_n796), .ZN(new_n1029));
  NAND4_X1  g843(.A1(new_n1027), .A2(new_n835), .A3(new_n841), .A4(new_n1029), .ZN(new_n1030));
  AND2_X1   g844(.A1(new_n1030), .A2(new_n348), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n1024), .B1(new_n1031), .B2(new_n1023), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1017), .B1(new_n1032), .B2(new_n702), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1033), .B1(new_n1017), .B2(new_n1032), .ZN(G72));
  NAND2_X1  g848(.A1(G472), .A2(G902), .ZN(new_n1035));
  XOR2_X1   g849(.A(new_n1035), .B(KEYINPUT63), .Z(new_n1036));
  NAND3_X1  g850(.A1(new_n716), .A2(new_n309), .A3(new_n1036), .ZN(new_n1037));
  NOR2_X1   g851(.A1(new_n915), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g852(.A(new_n1036), .B1(new_n1021), .B2(new_n1011), .ZN(new_n1039));
  INV_X1    g853(.A(new_n309), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1041), .A2(new_n951), .ZN(new_n1042));
  INV_X1    g856(.A(new_n716), .ZN(new_n1043));
  OAI21_X1  g857(.A(new_n1036), .B1(new_n1030), .B2(new_n1011), .ZN(new_n1044));
  AOI211_X1 g858(.A(new_n1038), .B(new_n1042), .C1(new_n1043), .C2(new_n1044), .ZN(G57));
endmodule


