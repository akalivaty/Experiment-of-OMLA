//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 1 0 0 0 0 1 1 0 0 1 1 0 1 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 0 1 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n568, new_n569, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT66), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  OR2_X1    g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n465), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  OR2_X1    g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n467), .A2(G101), .A3(G2104), .ZN(new_n473));
  OR2_X1    g048(.A1(new_n473), .A2(KEYINPUT67), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(KEYINPUT67), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n472), .A2(G137), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n468), .A2(new_n476), .ZN(G160));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G112), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n471), .A2(new_n467), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(new_n481), .B2(G124), .ZN(new_n482));
  OR3_X1    g057(.A1(new_n471), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n483));
  OAI21_X1  g058(.A(KEYINPUT68), .B1(new_n471), .B2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(G136), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n482), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  XOR2_X1   g062(.A(new_n487), .B(KEYINPUT69), .Z(G162));
  NAND2_X1  g063(.A1(new_n467), .A2(G138), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n489), .B1(new_n463), .B2(new_n464), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  OAI21_X1  g066(.A(KEYINPUT70), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT72), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(new_n469), .B2(new_n470), .ZN(new_n496));
  XNOR2_X1  g071(.A(KEYINPUT71), .B(KEYINPUT4), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n493), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n491), .A2(KEYINPUT71), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n465), .A2(new_n502), .A3(KEYINPUT72), .A4(new_n495), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n496), .A2(new_n504), .A3(KEYINPUT4), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n492), .A2(new_n498), .A3(new_n503), .A4(new_n505), .ZN(new_n506));
  OAI21_X1  g081(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n507));
  INV_X1    g082(.A(G114), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(G2105), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n509), .B1(new_n481), .B2(G126), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n515), .B1(KEYINPUT5), .B2(new_n516), .ZN(new_n517));
  NOR3_X1   g092(.A1(new_n513), .A2(KEYINPUT73), .A3(G543), .ZN(new_n518));
  OAI211_X1 g093(.A(G62), .B(new_n514), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT74), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g096(.A(KEYINPUT73), .B1(new_n513), .B2(G543), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT5), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n524), .A2(KEYINPUT74), .A3(G62), .A4(new_n514), .ZN(new_n525));
  NAND2_X1  g100(.A1(G75), .A2(G543), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n521), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT75), .ZN(new_n529));
  INV_X1    g104(.A(G651), .ZN(new_n530));
  INV_X1    g105(.A(new_n526), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n531), .B1(new_n519), .B2(new_n520), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n530), .B1(new_n532), .B2(new_n525), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT75), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g110(.A(KEYINPUT6), .B(G651), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n524), .A2(new_n514), .A3(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n538), .A2(G88), .B1(G50), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n529), .A2(new_n535), .A3(new_n541), .ZN(G303));
  INV_X1    g117(.A(G303), .ZN(G166));
  AND2_X1   g118(.A1(new_n524), .A2(new_n514), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n544), .A2(G63), .A3(G651), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT76), .B(KEYINPUT7), .Z(new_n546));
  NAND3_X1  g121(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n546), .B(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n540), .A2(G51), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n545), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n538), .A2(G89), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n550), .A2(new_n551), .ZN(G168));
  AOI22_X1  g127(.A1(new_n544), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(new_n530), .ZN(new_n554));
  INV_X1    g129(.A(G90), .ZN(new_n555));
  INV_X1    g130(.A(G52), .ZN(new_n556));
  OAI22_X1  g131(.A1(new_n537), .A2(new_n555), .B1(new_n539), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n554), .A2(new_n557), .ZN(G171));
  NAND2_X1  g133(.A1(new_n544), .A2(G56), .ZN(new_n559));
  NAND2_X1  g134(.A1(G68), .A2(G543), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n530), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n544), .A2(G81), .A3(new_n536), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n540), .A2(G43), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  NAND4_X1  g141(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND4_X1  g144(.A1(G319), .A2(G483), .A3(G661), .A4(new_n569), .ZN(G188));
  AOI22_X1  g145(.A1(new_n544), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  AND3_X1   g147(.A1(new_n540), .A2(new_n572), .A3(G53), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n572), .B1(new_n540), .B2(G53), .ZN(new_n574));
  OAI22_X1  g149(.A1(new_n571), .A2(new_n530), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n544), .A2(KEYINPUT77), .A3(new_n536), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT77), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n537), .A2(new_n577), .ZN(new_n578));
  AND3_X1   g153(.A1(new_n576), .A2(G91), .A3(new_n578), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G299));
  INV_X1    g156(.A(G171), .ZN(G301));
  INV_X1    g157(.A(G168), .ZN(G286));
  NAND3_X1  g158(.A1(new_n576), .A2(G87), .A3(new_n578), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n524), .A2(new_n514), .ZN(new_n585));
  INV_X1    g160(.A(G74), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n587), .A2(G651), .B1(G49), .B2(new_n540), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n584), .A2(new_n588), .ZN(G288));
  NAND3_X1  g164(.A1(new_n524), .A2(G61), .A3(new_n514), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n530), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n592), .A2(new_n593), .B1(new_n540), .B2(G48), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n576), .A2(G86), .A3(new_n578), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(G305));
  AOI22_X1  g172(.A1(new_n538), .A2(G85), .B1(G47), .B2(new_n540), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n544), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n530), .B2(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n576), .A2(G92), .A3(new_n578), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n602), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n585), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n607), .A2(G651), .B1(new_n540), .B2(G54), .ZN(new_n608));
  AND2_X1   g183(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n601), .B1(new_n609), .B2(G868), .ZN(G321));
  XNOR2_X1  g185(.A(G321), .B(KEYINPUT79), .ZN(G284));
  NAND2_X1  g186(.A1(G286), .A2(G868), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n580), .ZN(G297));
  OAI21_X1  g188(.A(new_n612), .B1(G868), .B2(new_n580), .ZN(G280));
  NAND2_X1  g189(.A1(new_n604), .A2(new_n608), .ZN(new_n615));
  OR2_X1    g190(.A1(new_n615), .A2(G559), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n617), .B1(G860), .B2(new_n609), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT80), .ZN(G148));
  AOI22_X1  g194(.A1(new_n544), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n563), .B(new_n562), .C1(new_n620), .C2(new_n530), .ZN(new_n621));
  INV_X1    g196(.A(G868), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(new_n617), .B2(new_n622), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n481), .A2(G123), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT81), .Z(new_n627));
  AND2_X1   g202(.A1(new_n483), .A2(new_n484), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G135), .ZN(new_n629));
  OR2_X1    g204(.A1(G99), .A2(G2105), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n630), .B(G2104), .C1(G111), .C2(new_n467), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n627), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n632), .A2(G2096), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(G2096), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2100), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n633), .A2(new_n634), .A3(new_n638), .ZN(G156));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(KEYINPUT14), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2451), .B(G2454), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n645), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT82), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n654), .A2(KEYINPUT83), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT83), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n650), .A2(new_n656), .A3(new_n653), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n650), .A2(new_n653), .ZN(new_n659));
  INV_X1    g234(.A(G14), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n658), .A2(new_n661), .ZN(G401));
  XOR2_X1   g237(.A(G2067), .B(G2678), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT84), .ZN(new_n664));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  XNOR2_X1  g240(.A(G2084), .B(G2090), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT85), .B(KEYINPUT18), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n665), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n664), .A2(new_n666), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n670), .B1(new_n671), .B2(KEYINPUT17), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n671), .A2(KEYINPUT17), .A3(new_n670), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n673), .B1(new_n664), .B2(new_n666), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n669), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT86), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2096), .B(G2100), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(G227));
  XOR2_X1   g256(.A(G1971), .B(G1976), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  XOR2_X1   g258(.A(G1956), .B(G2474), .Z(new_n684));
  XOR2_X1   g259(.A(G1961), .B(G1966), .Z(new_n685));
  AND2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT20), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n684), .A2(new_n685), .ZN(new_n689));
  NOR3_X1   g264(.A1(new_n683), .A2(new_n686), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(new_n683), .B2(new_n689), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(G1991), .B(G1996), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1981), .B(G1986), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(G229));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G33), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT25), .Z(new_n703));
  INV_X1    g278(.A(G139), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n703), .B1(new_n485), .B2(new_n704), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n705), .A2(KEYINPUT92), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(KEYINPUT92), .ZN(new_n707));
  NAND2_X1  g282(.A1(G115), .A2(G2104), .ZN(new_n708));
  INV_X1    g283(.A(G127), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n471), .B2(new_n709), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n706), .A2(new_n707), .B1(G2105), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n701), .B1(new_n711), .B2(new_n700), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT93), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT94), .ZN(new_n714));
  INV_X1    g289(.A(G2072), .ZN(new_n715));
  OR3_X1    g290(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n714), .B1(new_n713), .B2(new_n715), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n700), .A2(G32), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n628), .A2(G141), .ZN(new_n719));
  AND3_X1   g294(.A1(new_n467), .A2(G105), .A3(G2104), .ZN(new_n720));
  NAND3_X1  g295(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT26), .ZN(new_n722));
  AOI211_X1 g297(.A(new_n720), .B(new_n722), .C1(G129), .C2(new_n481), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n719), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n718), .B1(new_n724), .B2(G29), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT27), .B(G1996), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT24), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n700), .B1(new_n727), .B2(G34), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n727), .B2(G34), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G160), .B2(G29), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n725), .A2(new_n726), .B1(G2084), .B2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(new_n713), .B2(new_n715), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n716), .A2(new_n717), .A3(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT95), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n716), .A2(KEYINPUT95), .A3(new_n717), .A4(new_n733), .ZN(new_n737));
  INV_X1    g312(.A(G16), .ZN(new_n738));
  NOR2_X1   g313(.A1(G168), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n738), .B2(G21), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT96), .B(G1966), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT97), .Z(new_n743));
  NAND2_X1  g318(.A1(new_n738), .A2(G5), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G171), .B2(new_n738), .ZN(new_n745));
  INV_X1    g320(.A(G1961), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n700), .A2(G35), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G162), .B2(new_n700), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n750));
  INV_X1    g325(.A(G2090), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n749), .B(new_n752), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n743), .A2(new_n747), .A3(new_n753), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT89), .B(G16), .Z(new_n755));
  MUX2_X1   g330(.A(new_n621), .B(G19), .S(new_n755), .Z(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G1341), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n700), .A2(G26), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT28), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n628), .A2(G140), .ZN(new_n760));
  OAI21_X1  g335(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n761));
  INV_X1    g336(.A(G116), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n761), .B1(new_n762), .B2(G2105), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n481), .B2(G128), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n759), .B1(new_n765), .B2(G29), .ZN(new_n766));
  INV_X1    g341(.A(G2067), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n757), .A2(new_n768), .ZN(new_n769));
  OAI22_X1  g344(.A1(new_n740), .A2(new_n741), .B1(new_n725), .B2(new_n726), .ZN(new_n770));
  INV_X1    g345(.A(G28), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n771), .A2(KEYINPUT30), .ZN(new_n772));
  AOI21_X1  g347(.A(G29), .B1(new_n771), .B2(KEYINPUT30), .ZN(new_n773));
  OR2_X1    g348(.A1(KEYINPUT31), .A2(G11), .ZN(new_n774));
  NAND2_X1  g349(.A1(KEYINPUT31), .A2(G11), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n772), .A2(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI221_X1 g351(.A(new_n776), .B1(new_n730), .B2(G2084), .C1(new_n632), .C2(new_n700), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n770), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n755), .A2(G20), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT23), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n580), .B2(new_n738), .ZN(new_n781));
  INV_X1    g356(.A(G1956), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(G27), .A2(G29), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G164), .B2(G29), .ZN(new_n785));
  INV_X1    g360(.A(G2078), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n769), .A2(new_n778), .A3(new_n783), .A4(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(G4), .A2(G16), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT91), .Z(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n609), .B2(G16), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G1348), .ZN(new_n792));
  NOR3_X1   g367(.A1(new_n754), .A2(new_n788), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n736), .A2(new_n737), .A3(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT36), .ZN(new_n795));
  MUX2_X1   g370(.A(G6), .B(G305), .S(G16), .Z(new_n796));
  XOR2_X1   g371(.A(KEYINPUT32), .B(G1981), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n738), .A2(G23), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G288), .B2(G16), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT33), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(G1976), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n800), .A2(new_n801), .ZN(new_n804));
  AND3_X1   g379(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n803), .B1(new_n802), .B2(new_n804), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n798), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n755), .A2(G22), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G166), .B2(new_n755), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G1971), .ZN(new_n810));
  OAI21_X1  g385(.A(KEYINPUT34), .B1(new_n807), .B2(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT90), .ZN(new_n812));
  NOR3_X1   g387(.A1(new_n807), .A2(KEYINPUT34), .A3(new_n810), .ZN(new_n813));
  NOR2_X1   g388(.A1(G25), .A2(G29), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n481), .A2(G119), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n467), .A2(G107), .ZN(new_n816));
  OAI21_X1  g391(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n817));
  INV_X1    g392(.A(G131), .ZN(new_n818));
  OAI221_X1 g393(.A(new_n815), .B1(new_n816), .B2(new_n817), .C1(new_n485), .C2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT87), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n814), .B1(new_n820), .B2(G29), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT35), .B(G1991), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT88), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n821), .B(new_n823), .ZN(new_n824));
  MUX2_X1   g399(.A(G290), .B(G24), .S(new_n755), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1986), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n813), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n795), .B1(new_n812), .B2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n812), .A2(new_n827), .A3(new_n795), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n794), .B1(new_n829), .B2(new_n830), .ZN(G311));
  INV_X1    g406(.A(new_n794), .ZN(new_n832));
  INV_X1    g407(.A(new_n830), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(new_n828), .ZN(G150));
  AND2_X1   g409(.A1(new_n544), .A2(G67), .ZN(new_n835));
  AND2_X1   g410(.A1(G80), .A2(G543), .ZN(new_n836));
  OAI21_X1  g411(.A(G651), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n538), .A2(G93), .B1(G55), .B2(new_n540), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XOR2_X1   g414(.A(KEYINPUT101), .B(G860), .Z(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT37), .Z(new_n842));
  NAND2_X1  g417(.A1(new_n609), .A2(G559), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT38), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT99), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n621), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(new_n839), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT100), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(new_n565), .B2(KEYINPUT99), .ZN(new_n849));
  NOR3_X1   g424(.A1(new_n621), .A2(new_n845), .A3(KEYINPUT100), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n847), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AOI22_X1  g426(.A1(new_n621), .A2(new_n845), .B1(new_n837), .B2(new_n838), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n565), .A2(KEYINPUT99), .A3(new_n848), .ZN(new_n853));
  OAI21_X1  g428(.A(KEYINPUT100), .B1(new_n621), .B2(new_n845), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n844), .B(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(KEYINPUT39), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT102), .Z(new_n859));
  NOR2_X1   g434(.A1(new_n857), .A2(KEYINPUT39), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n860), .A2(new_n840), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n842), .B1(new_n859), .B2(new_n861), .ZN(G145));
  INV_X1    g437(.A(new_n820), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n481), .A2(G130), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n467), .A2(G118), .ZN(new_n865));
  OAI21_X1  g440(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(new_n628), .B2(G142), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(new_n636), .Z(new_n869));
  XNOR2_X1  g444(.A(new_n863), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n724), .A2(new_n765), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n719), .A2(new_n760), .A3(new_n723), .A4(new_n764), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n711), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n711), .A2(new_n873), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n511), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n711), .A2(new_n873), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n878), .A2(G164), .A3(new_n874), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n870), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(G162), .B(G160), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n632), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n869), .B(new_n820), .ZN(new_n885));
  NOR3_X1   g460(.A1(new_n875), .A2(new_n876), .A3(new_n511), .ZN(new_n886));
  AOI21_X1  g461(.A(G164), .B1(new_n878), .B2(new_n874), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(G37), .B1(new_n884), .B2(new_n888), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n870), .A2(new_n877), .A3(KEYINPUT103), .A4(new_n879), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n883), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n888), .A2(new_n892), .A3(new_n880), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n891), .A2(KEYINPUT104), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(KEYINPUT104), .B1(new_n891), .B2(new_n893), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n889), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n604), .A2(new_n580), .A3(new_n608), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n580), .B1(new_n604), .B2(new_n608), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n901), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n903), .A2(KEYINPUT105), .A3(new_n899), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n617), .A2(new_n856), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n616), .B1(new_n855), .B2(new_n851), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n902), .B(new_n904), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n905), .A2(new_n906), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT41), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(new_n900), .B2(new_n901), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n903), .A2(KEYINPUT41), .A3(new_n899), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n907), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(KEYINPUT42), .ZN(new_n914));
  XOR2_X1   g489(.A(G303), .B(G305), .Z(new_n915));
  XNOR2_X1  g490(.A(G288), .B(G290), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n915), .B(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n918), .A2(KEYINPUT106), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT42), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n907), .B(new_n920), .C1(new_n908), .C2(new_n912), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n914), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n919), .B1(new_n914), .B2(new_n921), .ZN(new_n923));
  OAI21_X1  g498(.A(G868), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n839), .A2(new_n622), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(G295));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n925), .ZN(G331));
  AND3_X1   g502(.A1(new_n851), .A2(G301), .A3(new_n855), .ZN(new_n928));
  AOI21_X1  g503(.A(G301), .B1(new_n851), .B2(new_n855), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n928), .A2(new_n929), .A3(G286), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n852), .B1(new_n854), .B2(new_n853), .ZN(new_n932));
  OAI21_X1  g507(.A(G171), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n851), .A2(G301), .A3(new_n855), .ZN(new_n934));
  AOI21_X1  g509(.A(G168), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n912), .B1(new_n930), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(G286), .B1(new_n928), .B2(new_n929), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n933), .A2(G168), .A3(new_n934), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n937), .A2(new_n938), .A3(new_n903), .A4(new_n899), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n936), .A2(new_n918), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G37), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n918), .B1(new_n936), .B2(new_n939), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT43), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n902), .A2(new_n904), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n937), .A2(new_n945), .A3(new_n938), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n936), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(new_n917), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT43), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n948), .A2(new_n949), .A3(new_n940), .A4(new_n941), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n944), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n948), .A2(new_n941), .A3(new_n940), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n955));
  INV_X1    g530(.A(new_n943), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n956), .A2(new_n949), .A3(new_n940), .A4(new_n941), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n955), .A2(KEYINPUT44), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n953), .A2(new_n958), .ZN(G397));
  INV_X1    g534(.A(G1384), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n511), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n468), .A2(G40), .A3(new_n476), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n765), .A2(G2067), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n760), .A2(new_n767), .A3(new_n764), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n965), .B1(new_n969), .B2(new_n724), .ZN(new_n970));
  INV_X1    g545(.A(new_n965), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n971), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT46), .ZN(new_n973));
  INV_X1    g548(.A(G1996), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n973), .B1(new_n965), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n970), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  XOR2_X1   g551(.A(new_n976), .B(KEYINPUT47), .Z(new_n977));
  XNOR2_X1  g552(.A(new_n724), .B(new_n974), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n968), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n979), .B1(new_n823), .B2(new_n863), .ZN(new_n980));
  OR2_X1    g555(.A1(new_n863), .A2(new_n823), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n965), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n971), .A2(G1986), .A3(G290), .ZN(new_n984));
  OR2_X1    g559(.A1(new_n984), .A2(KEYINPUT48), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n986), .B1(KEYINPUT48), .B2(new_n984), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n967), .B1(new_n981), .B2(new_n979), .ZN(new_n988));
  AOI211_X1 g563(.A(new_n977), .B(new_n987), .C1(new_n965), .C2(new_n988), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n584), .A2(new_n588), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n990), .A2(G1976), .ZN(new_n991));
  INV_X1    g566(.A(G8), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n468), .A2(G40), .A3(new_n476), .ZN(new_n993));
  AOI21_X1  g568(.A(G1384), .B1(new_n506), .B2(new_n510), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT52), .B1(new_n991), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n997), .B1(new_n990), .B2(G1976), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n995), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n998), .B(new_n995), .C1(new_n991), .C2(KEYINPUT52), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1981), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n594), .A2(new_n595), .A3(new_n596), .A4(new_n1003), .ZN(new_n1004));
  XOR2_X1   g579(.A(KEYINPUT113), .B(G86), .Z(new_n1005));
  INV_X1    g580(.A(G48), .ZN(new_n1006));
  OAI22_X1  g581(.A1(new_n537), .A2(new_n1005), .B1(new_n539), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(G1981), .B1(new_n1007), .B2(new_n592), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT114), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT49), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1004), .A2(new_n1008), .A3(new_n1011), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1012), .A2(new_n995), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1004), .A2(new_n1008), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1014), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1002), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n541), .B1(new_n533), .B2(new_n534), .ZN(new_n1018));
  AOI211_X1 g593(.A(KEYINPUT75), .B(new_n530), .C1(new_n532), .C2(new_n525), .ZN(new_n1019));
  OAI21_X1  g594(.A(G8), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT110), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT111), .ZN(new_n1023));
  NAND4_X1  g598(.A1(G303), .A2(new_n1023), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1024));
  OAI211_X1 g599(.A(KEYINPUT55), .B(G8), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT111), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n1022), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT110), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1026), .A2(new_n1024), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT109), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n961), .A2(new_n1032), .A3(new_n962), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT109), .B1(new_n994), .B2(KEYINPUT45), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n964), .B1(new_n994), .B2(KEYINPUT45), .ZN(new_n1036));
  AOI21_X1  g611(.A(G1971), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n961), .A2(KEYINPUT50), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n994), .A2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1038), .A2(new_n751), .A3(new_n993), .A4(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(G8), .B1(new_n1037), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1017), .B1(new_n1031), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1032), .B1(new_n961), .B2(new_n962), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n994), .A2(KEYINPUT109), .A3(KEYINPUT45), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1036), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G1971), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n992), .B1(new_n1049), .B2(new_n1041), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n511), .A2(KEYINPUT45), .A3(new_n960), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n993), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n994), .A2(KEYINPUT45), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n741), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G2084), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1038), .A2(new_n1056), .A3(new_n993), .A4(new_n1040), .ZN(new_n1057));
  AOI211_X1 g632(.A(new_n992), .B(G286), .C1(new_n1055), .C2(new_n1057), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1044), .A2(KEYINPUT63), .A3(new_n1051), .A4(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1026), .A2(new_n1024), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1022), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1043), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n1000), .A2(new_n1001), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1051), .A2(new_n1064), .A3(new_n1065), .A4(new_n1058), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT63), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1059), .A2(new_n1068), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1051), .A2(new_n1065), .A3(new_n1064), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1055), .A2(G168), .A3(new_n1057), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(G8), .ZN(new_n1072));
  AOI21_X1  g647(.A(G168), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT51), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1071), .A2(new_n1075), .A3(G8), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT62), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n786), .B(new_n1036), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1040), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n993), .B1(new_n994), .B2(new_n1039), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT118), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1038), .A2(new_n1085), .A3(new_n993), .A4(new_n1040), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1084), .A2(new_n746), .A3(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n963), .A2(new_n1036), .A3(KEYINPUT53), .A4(new_n786), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1081), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(G171), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT62), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1074), .A2(new_n1092), .A3(new_n1076), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1070), .A2(new_n1078), .A3(new_n1091), .A4(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n995), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1016), .A2(new_n803), .A3(new_n990), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(new_n1004), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT115), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1095), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1096), .A2(KEYINPUT115), .A3(new_n1004), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1051), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1099), .A2(new_n1100), .B1(new_n1101), .B2(new_n1065), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1069), .A2(new_n1094), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n1104));
  OR2_X1    g679(.A1(new_n786), .A2(KEYINPUT123), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n786), .A2(KEYINPUT123), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1080), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n963), .A2(new_n1036), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT124), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n963), .A2(new_n1036), .A3(KEYINPUT124), .A4(new_n1107), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1112), .A2(new_n1081), .A3(new_n1087), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1104), .B1(new_n1113), .B2(G171), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1081), .A2(new_n1087), .A3(G301), .A4(new_n1088), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1114), .A2(KEYINPUT126), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT126), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1077), .B(new_n1070), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1112), .A2(new_n1081), .A3(new_n1087), .A4(G301), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1090), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT125), .B1(new_n1120), .B2(new_n1104), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT125), .ZN(new_n1122));
  AOI211_X1 g697(.A(new_n1122), .B(KEYINPUT54), .C1(new_n1090), .C2(new_n1119), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1118), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT60), .ZN(new_n1126));
  INV_X1    g701(.A(G1348), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1084), .A2(new_n1127), .A3(new_n1086), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n993), .A2(new_n994), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1128), .B1(G2067), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n609), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1128), .B(new_n615), .C1(G2067), .C2(new_n1129), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1126), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n565), .A2(KEYINPUT121), .ZN(new_n1134));
  XNOR2_X1  g709(.A(KEYINPUT120), .B(G1996), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1036), .B(new_n1136), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1137));
  XOR2_X1   g712(.A(KEYINPUT58), .B(G1341), .Z(new_n1138));
  NAND2_X1  g713(.A1(new_n1129), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1134), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT59), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI211_X1 g717(.A(KEYINPUT59), .B(new_n1134), .C1(new_n1137), .C2(new_n1139), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n609), .A2(new_n1126), .ZN(new_n1144));
  OAI22_X1  g719(.A1(new_n1142), .A2(new_n1143), .B1(new_n1130), .B2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1133), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1053), .B1(new_n1034), .B2(new_n1033), .ZN(new_n1147));
  XNOR2_X1  g722(.A(KEYINPUT56), .B(G2072), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1147), .A2(KEYINPUT117), .A3(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1036), .B(new_n1148), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT117), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1038), .A2(new_n993), .A3(new_n1040), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(new_n782), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1149), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT116), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n580), .A2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1157), .B(KEYINPUT57), .ZN(new_n1158));
  OR2_X1    g733(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1154), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1160));
  AOI21_X1  g735(.A(KEYINPUT117), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1158), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1159), .A2(KEYINPUT61), .A3(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1162), .A2(KEYINPUT122), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT122), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1155), .A2(new_n1166), .A3(new_n1158), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1164), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1146), .B(new_n1163), .C1(new_n1168), .C2(KEYINPUT61), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1131), .A2(new_n1162), .ZN(new_n1170));
  AND3_X1   g745(.A1(new_n1159), .A2(new_n1170), .A3(KEYINPUT119), .ZN(new_n1171));
  AOI21_X1  g746(.A(KEYINPUT119), .B1(new_n1159), .B2(new_n1170), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1169), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1103), .B1(new_n1125), .B2(new_n1174), .ZN(new_n1175));
  AND3_X1   g750(.A1(new_n965), .A2(G1986), .A3(G290), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n984), .A2(new_n1176), .ZN(new_n1177));
  XOR2_X1   g752(.A(new_n1177), .B(KEYINPUT108), .Z(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(new_n983), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n989), .B1(new_n1175), .B2(new_n1179), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g755(.A1(new_n679), .A2(G319), .A3(new_n680), .ZN(new_n1182));
  NOR3_X1   g756(.A1(G401), .A2(KEYINPUT127), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g757(.A(KEYINPUT127), .ZN(new_n1184));
  INV_X1    g758(.A(new_n1182), .ZN(new_n1185));
  NAND2_X1  g759(.A1(new_n658), .A2(new_n661), .ZN(new_n1186));
  AOI21_X1  g760(.A(new_n1184), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NOR3_X1   g761(.A1(new_n1183), .A2(new_n1187), .A3(G229), .ZN(new_n1188));
  AND3_X1   g762(.A1(new_n1188), .A2(new_n951), .A3(new_n896), .ZN(G308));
  NAND3_X1  g763(.A1(new_n1188), .A2(new_n951), .A3(new_n896), .ZN(G225));
endmodule


