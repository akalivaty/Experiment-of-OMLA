//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 1 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT28), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT11), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G137), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT11), .A3(G134), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n190), .A2(G137), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G131), .ZN(new_n196));
  INV_X1    g010(.A(G131), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n191), .A2(new_n193), .A3(new_n197), .A4(new_n194), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT66), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT64), .B(G146), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G143), .ZN(new_n205));
  AND2_X1   g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  NOR2_X1   g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n202), .A2(G143), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n209), .B1(new_n204), .B2(G143), .ZN(new_n210));
  AOI22_X1  g024(.A1(new_n205), .A2(new_n208), .B1(new_n210), .B2(new_n206), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n196), .A2(KEYINPUT66), .A3(new_n198), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n201), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n202), .A2(KEYINPUT64), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G146), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n214), .A2(new_n216), .A3(G143), .ZN(new_n217));
  INV_X1    g031(.A(new_n209), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n217), .A2(G128), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G128), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT65), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n221), .B1(new_n217), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n203), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n214), .A2(new_n216), .ZN(new_n229));
  INV_X1    g043(.A(G143), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n220), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n194), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n190), .A2(G137), .ZN(new_n234));
  OAI21_X1  g048(.A(G131), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n235), .A2(new_n198), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n232), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n213), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT2), .B(G113), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(G116), .B(G119), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n241), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n239), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n238), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n245), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n213), .A2(new_n247), .A3(new_n237), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n188), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n248), .A2(new_n188), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(G237), .A2(G953), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G210), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n253), .B(KEYINPUT27), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT26), .B(G101), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n254), .B(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT29), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(G902), .B1(new_n251), .B2(new_n259), .ZN(new_n260));
  XOR2_X1   g074(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n261));
  AND3_X1   g075(.A1(new_n213), .A2(new_n247), .A3(new_n237), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n211), .A2(new_n199), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n247), .B1(new_n263), .B2(new_n237), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n261), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT69), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n248), .A2(new_n188), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n265), .A2(new_n266), .A3(new_n256), .A4(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT30), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n232), .A2(new_n236), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n217), .A2(new_n206), .A3(new_n218), .ZN(new_n271));
  AOI21_X1  g085(.A(G143), .B1(new_n214), .B2(new_n216), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n208), .B1(new_n272), .B2(new_n228), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n199), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n269), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n213), .A2(KEYINPUT30), .A3(new_n237), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(new_n276), .A3(new_n245), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n248), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n257), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n268), .A2(new_n279), .A3(new_n258), .ZN(new_n280));
  INV_X1    g094(.A(new_n261), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n245), .B1(new_n270), .B2(new_n274), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n281), .B1(new_n282), .B2(new_n248), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(new_n250), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n266), .B1(new_n284), .B2(new_n256), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n260), .B1(new_n280), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n187), .B1(new_n286), .B2(G472), .ZN(new_n287));
  INV_X1    g101(.A(G472), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n265), .A2(new_n256), .A3(new_n267), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT69), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT29), .B1(new_n278), .B2(new_n257), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(new_n268), .A3(new_n291), .ZN(new_n292));
  AOI211_X1 g106(.A(KEYINPUT70), .B(new_n288), .C1(new_n292), .C2(new_n260), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n257), .B1(new_n283), .B2(new_n250), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT31), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n277), .A2(new_n295), .A3(new_n256), .A4(new_n248), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n277), .A2(new_n256), .A3(new_n248), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT31), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT67), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n298), .A2(KEYINPUT67), .A3(KEYINPUT31), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n297), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(G472), .A2(G902), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NOR3_X1   g119(.A1(new_n303), .A2(KEYINPUT32), .A3(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT32), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n294), .A2(new_n296), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n298), .A2(KEYINPUT67), .A3(KEYINPUT31), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT67), .B1(new_n298), .B2(KEYINPUT31), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n307), .B1(new_n311), .B2(new_n304), .ZN(new_n312));
  OAI22_X1  g126(.A1(new_n287), .A2(new_n293), .B1(new_n306), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G469), .ZN(new_n314));
  INV_X1    g128(.A(G902), .ZN(new_n315));
  INV_X1    g129(.A(G104), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT3), .B1(new_n316), .B2(G107), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT3), .ZN(new_n318));
  INV_X1    g132(.A(G107), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(new_n319), .A3(G104), .ZN(new_n320));
  INV_X1    g134(.A(G101), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n316), .A2(G107), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n317), .A2(new_n320), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n319), .A2(G104), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n316), .A2(G107), .ZN(new_n325));
  OAI21_X1  g139(.A(G101), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n220), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n203), .A2(KEYINPUT1), .ZN(new_n330));
  AOI22_X1  g144(.A1(new_n217), .A2(new_n218), .B1(new_n330), .B2(G128), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n328), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n327), .B(new_n220), .C1(new_n227), .C2(new_n231), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n212), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT66), .B1(new_n196), .B2(new_n198), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT12), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n339), .B1(new_n196), .B2(new_n198), .ZN(new_n340));
  AOI22_X1  g154(.A1(new_n338), .A2(new_n339), .B1(new_n334), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT10), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n332), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n327), .A2(KEYINPUT79), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n323), .A2(new_n326), .A3(new_n345), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n232), .A2(KEYINPUT10), .A3(new_n344), .A4(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n317), .A2(new_n320), .A3(new_n322), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G101), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(KEYINPUT4), .A3(new_n323), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT4), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n348), .A2(new_n351), .A3(G101), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n211), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n201), .A2(new_n212), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n343), .A2(new_n347), .A3(new_n353), .A4(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(G110), .B(G140), .ZN(new_n356));
  INV_X1    g170(.A(G953), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n357), .A2(G227), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n356), .B(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n341), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n217), .A2(new_n218), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n330), .A2(G128), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n327), .B1(new_n365), .B2(new_n220), .ZN(new_n366));
  INV_X1    g180(.A(new_n350), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n273), .A2(new_n352), .A3(new_n271), .ZN(new_n368));
  OAI22_X1  g182(.A1(new_n366), .A2(KEYINPUT10), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  AND4_X1   g183(.A1(KEYINPUT10), .A2(new_n232), .A3(new_n344), .A4(new_n346), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n337), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n360), .B1(new_n371), .B2(new_n355), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n314), .B(new_n315), .C1(new_n362), .C2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n355), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n359), .B1(new_n341), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n371), .A2(new_n360), .A3(new_n355), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n376), .A3(G469), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n314), .A2(new_n315), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n373), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G221), .ZN(new_n381));
  XNOR2_X1  g195(.A(KEYINPUT9), .B(G234), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(KEYINPUT78), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n381), .B1(new_n383), .B2(new_n315), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT80), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(G214), .B1(G237), .B2(G902), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(G210), .B1(G237), .B2(G902), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G125), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n393), .B(new_n220), .C1(new_n227), .C2(new_n231), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n394), .B1(new_n211), .B2(new_n393), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT81), .B(G224), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(G953), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT82), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(KEYINPUT7), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G113), .ZN(new_n404));
  INV_X1    g218(.A(G119), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G116), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT5), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n404), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n241), .A2(KEYINPUT5), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n409), .A2(new_n410), .B1(new_n240), .B2(new_n241), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n344), .A2(new_n411), .A3(new_n346), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n350), .A2(new_n245), .A3(new_n352), .ZN(new_n413));
  XNOR2_X1  g227(.A(G110), .B(G122), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  OR2_X1    g229(.A1(new_n411), .A2(new_n327), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n411), .A2(new_n327), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n414), .B(KEYINPUT8), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n395), .A2(new_n399), .A3(new_n401), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n403), .A2(new_n415), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT83), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n421), .A2(new_n422), .A3(new_n315), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n412), .A2(new_n413), .ZN(new_n424));
  INV_X1    g238(.A(new_n414), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n426), .A2(KEYINPUT6), .A3(new_n415), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n395), .B(new_n397), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT6), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n424), .A2(new_n429), .A3(new_n425), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n427), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n423), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n422), .B1(new_n421), .B2(new_n315), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n392), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n421), .A2(new_n315), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT83), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n436), .A2(new_n391), .A3(new_n431), .A4(new_n423), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n390), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n380), .A2(KEYINPUT80), .A3(new_n385), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n388), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT74), .ZN(new_n441));
  INV_X1    g255(.A(G140), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G125), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n393), .A2(G140), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n443), .A2(new_n444), .A3(KEYINPUT16), .ZN(new_n445));
  OR3_X1    g259(.A1(new_n393), .A2(KEYINPUT16), .A3(G140), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n441), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NOR3_X1   g261(.A1(new_n393), .A2(KEYINPUT16), .A3(G140), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n448), .A2(KEYINPUT74), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n202), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n446), .A2(new_n441), .ZN(new_n451));
  XNOR2_X1  g265(.A(G125), .B(G140), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n448), .B1(new_n452), .B2(KEYINPUT16), .ZN(new_n453));
  OAI211_X1 g267(.A(G146), .B(new_n451), .C1(new_n453), .C2(new_n441), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n450), .A2(new_n454), .A3(KEYINPUT75), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT75), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n456), .B(new_n202), .C1(new_n447), .C2(new_n449), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n221), .A2(G119), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n405), .A2(G128), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT24), .B(G110), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G110), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT23), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n464), .B1(new_n405), .B2(G128), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT72), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(new_n405), .B2(G128), .ZN(new_n467));
  NOR2_X1   g281(.A1(KEYINPUT72), .A2(KEYINPUT23), .ZN(new_n468));
  OAI22_X1  g282(.A1(new_n465), .A2(new_n467), .B1(new_n458), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT73), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n463), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT23), .B1(new_n221), .B2(G119), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT72), .B1(new_n221), .B2(G119), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n405), .A2(G128), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n466), .A2(new_n464), .ZN(new_n475));
  AOI22_X1  g289(.A1(new_n472), .A2(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT73), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n462), .B1(new_n471), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n455), .A2(new_n457), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n204), .A2(new_n452), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n476), .A2(new_n463), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT76), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n460), .A2(new_n461), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n482), .B1(new_n481), .B2(new_n483), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n454), .B(new_n480), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n479), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT22), .B(G137), .ZN(new_n488));
  INV_X1    g302(.A(G234), .ZN(new_n489));
  NOR3_X1   g303(.A1(new_n381), .A2(new_n489), .A3(G953), .ZN(new_n490));
  XOR2_X1   g304(.A(new_n488), .B(new_n490), .Z(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n479), .A2(new_n486), .A3(new_n491), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(G217), .B1(new_n489), .B2(G902), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n315), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n496), .B(KEYINPUT71), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n493), .A2(new_n315), .A3(new_n494), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT25), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT77), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n499), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n500), .A2(new_n501), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n493), .A2(KEYINPUT25), .A3(new_n315), .A4(new_n494), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(KEYINPUT77), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n498), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(G113), .B(G122), .ZN(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT86), .B(G104), .ZN(new_n510));
  XOR2_X1   g324(.A(new_n509), .B(new_n510), .Z(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(G237), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(new_n357), .A3(G214), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n514), .A2(new_n230), .ZN(new_n515));
  AOI21_X1  g329(.A(G143), .B1(new_n252), .B2(G214), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT18), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n517), .B1(new_n518), .B2(new_n197), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n480), .B1(new_n202), .B2(new_n452), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n514), .B(new_n230), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n518), .A2(new_n197), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n524), .A2(KEYINPUT84), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(KEYINPUT84), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n521), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n452), .A2(KEYINPUT85), .ZN(new_n529));
  XOR2_X1   g343(.A(new_n529), .B(KEYINPUT19), .Z(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n204), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n522), .A2(G131), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n517), .A2(new_n197), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n531), .A2(new_n534), .A3(new_n454), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n512), .B1(new_n528), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n522), .A2(KEYINPUT17), .A3(G131), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n537), .B1(new_n534), .B2(KEYINPUT17), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n455), .A2(new_n457), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n538), .B1(new_n539), .B2(KEYINPUT87), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT87), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n455), .A2(new_n541), .A3(new_n457), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n527), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n536), .B1(new_n543), .B2(new_n512), .ZN(new_n544));
  NOR2_X1   g358(.A1(G475), .A2(G902), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(KEYINPUT88), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT20), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n536), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n539), .A2(KEYINPUT87), .ZN(new_n549));
  INV_X1    g363(.A(new_n538), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(new_n542), .A3(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n551), .A2(new_n528), .A3(new_n512), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT20), .ZN(new_n554));
  INV_X1    g368(.A(new_n546), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AOI211_X1 g370(.A(new_n527), .B(new_n511), .C1(new_n540), .C2(new_n542), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n512), .B1(new_n551), .B2(new_n528), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n315), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n547), .A2(new_n556), .B1(new_n559), .B2(G475), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n357), .A2(G952), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n561), .B1(G234), .B2(G237), .ZN(new_n562));
  OAI211_X1 g376(.A(G902), .B(G953), .C1(new_n489), .C2(new_n513), .ZN(new_n563));
  XOR2_X1   g377(.A(new_n563), .B(KEYINPUT92), .Z(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT21), .B(G898), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n562), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(G478), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(KEYINPUT15), .ZN(new_n569));
  INV_X1    g383(.A(G116), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(G122), .ZN(new_n571));
  OR2_X1    g385(.A1(new_n571), .A2(KEYINPUT14), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(KEYINPUT14), .ZN(new_n573));
  INV_X1    g387(.A(G122), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(G116), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n572), .A2(new_n573), .A3(KEYINPUT90), .A4(new_n575), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n576), .B(G107), .C1(KEYINPUT90), .C2(new_n572), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n230), .A2(G128), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n221), .A2(G143), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(new_n190), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n575), .A2(new_n571), .A3(new_n319), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n577), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n575), .A2(new_n571), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(G107), .ZN(new_n585));
  AOI22_X1  g399(.A1(new_n585), .A2(new_n582), .B1(new_n580), .B2(new_n190), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT13), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n579), .B1(new_n578), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT13), .B1(new_n230), .B2(G128), .ZN(new_n589));
  OAI21_X1  g403(.A(G134), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT89), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n590), .A2(new_n591), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n586), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n383), .A2(G217), .A3(new_n357), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n583), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n595), .B1(new_n583), .B2(new_n594), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n315), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n569), .B1(new_n598), .B2(KEYINPUT91), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(KEYINPUT91), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT91), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n601), .B(new_n315), .C1(new_n596), .C2(new_n597), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n599), .B1(new_n603), .B2(new_n569), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n560), .A2(new_n567), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n313), .A2(new_n440), .A3(new_n508), .A4(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G101), .ZN(G3));
  AND3_X1   g422(.A1(new_n388), .A2(new_n508), .A3(new_n439), .ZN(new_n609));
  OAI21_X1  g423(.A(G472), .B1(new_n303), .B2(G902), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n311), .A2(new_n304), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(new_n613), .B(KEYINPUT93), .Z(new_n614));
  NAND2_X1  g428(.A1(new_n434), .A2(new_n437), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n615), .A2(new_n389), .A3(new_n567), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n559), .A2(G475), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n554), .B1(new_n553), .B2(new_n555), .ZN(new_n618));
  AOI211_X1 g432(.A(KEYINPUT20), .B(new_n546), .C1(new_n548), .C2(new_n552), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n598), .A2(G478), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n568), .A2(new_n315), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OR3_X1    g437(.A1(new_n596), .A2(new_n597), .A3(KEYINPUT33), .ZN(new_n624));
  OAI21_X1  g438(.A(KEYINPUT33), .B1(new_n596), .B2(new_n597), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(G478), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n620), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n616), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n614), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT94), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT34), .B(G104), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  INV_X1    g448(.A(new_n604), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n560), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n616), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n614), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT35), .B(G107), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  NOR2_X1   g454(.A1(new_n492), .A2(KEYINPUT36), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n487), .B(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n642), .A2(new_n315), .A3(new_n496), .ZN(new_n643));
  INV_X1    g457(.A(new_n507), .ZN(new_n644));
  INV_X1    g458(.A(new_n499), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n645), .B1(new_n505), .B2(KEYINPUT77), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n643), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT95), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI211_X1 g463(.A(KEYINPUT95), .B(new_n643), .C1(new_n644), .C2(new_n646), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n440), .A2(new_n651), .A3(new_n606), .A4(new_n612), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT96), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT37), .B(G110), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G12));
  INV_X1    g469(.A(new_n562), .ZN(new_n656));
  INV_X1    g470(.A(G900), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n564), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n656), .B1(new_n658), .B2(KEYINPUT97), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n659), .B1(KEYINPUT97), .B2(new_n658), .ZN(new_n660));
  XOR2_X1   g474(.A(new_n660), .B(KEYINPUT98), .Z(new_n661));
  NOR2_X1   g475(.A1(new_n636), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n313), .A2(new_n440), .A3(new_n651), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  XNOR2_X1  g478(.A(KEYINPUT100), .B(KEYINPUT39), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n661), .B(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n388), .A2(new_n439), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT101), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  OR2_X1    g483(.A1(new_n669), .A2(KEYINPUT40), .ZN(new_n670));
  INV_X1    g484(.A(new_n651), .ZN(new_n671));
  OAI21_X1  g485(.A(KEYINPUT32), .B1(new_n303), .B2(new_n305), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n311), .A2(new_n307), .A3(new_n304), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n246), .A2(new_n257), .A3(new_n248), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n315), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n257), .B1(new_n277), .B2(new_n248), .ZN(new_n677));
  OAI21_X1  g491(.A(G472), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(new_n678), .B(KEYINPUT99), .Z(new_n679));
  NAND2_X1  g493(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n615), .B(KEYINPUT38), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n560), .A2(new_n390), .A3(new_n604), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n671), .A2(new_n680), .A3(new_n681), .A4(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n683), .B1(new_n669), .B2(KEYINPUT40), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n670), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G143), .ZN(G45));
  NOR3_X1   g500(.A1(new_n560), .A2(new_n627), .A3(new_n661), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n313), .A2(new_n440), .A3(new_n651), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n315), .B1(new_n362), .B2(new_n372), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(G469), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n373), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n690), .B1(new_n693), .B2(new_n384), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n692), .A2(KEYINPUT102), .A3(new_n385), .A4(new_n373), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n694), .A2(new_n508), .A3(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n313), .A2(new_n630), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT41), .B(G113), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G15));
  NAND3_X1  g513(.A1(new_n313), .A2(new_n696), .A3(new_n637), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT103), .B(G116), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G18));
  AND3_X1   g516(.A1(new_n694), .A2(new_n438), .A3(new_n695), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n313), .A2(new_n703), .A3(new_n651), .A4(new_n606), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G119), .ZN(G21));
  OAI211_X1 g519(.A(new_n299), .B(new_n296), .C1(new_n251), .C2(new_n256), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n304), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n610), .A2(new_n508), .A3(new_n707), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n694), .A2(new_n695), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n438), .A2(new_n620), .A3(new_n635), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n708), .A2(new_n709), .A3(new_n710), .A4(new_n567), .ZN(new_n711));
  XOR2_X1   g525(.A(KEYINPUT104), .B(G122), .Z(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G24));
  AND2_X1   g527(.A1(new_n610), .A2(new_n707), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n703), .A2(new_n651), .A3(new_n687), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G125), .ZN(G27));
  NAND3_X1  g530(.A1(new_n434), .A2(new_n389), .A3(new_n437), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n386), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n434), .A2(new_n437), .A3(KEYINPUT105), .A4(new_n389), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n722), .A2(new_n313), .A3(new_n508), .A4(new_n687), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT42), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n508), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n286), .A2(G472), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(KEYINPUT70), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n286), .A2(new_n187), .A3(G472), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n726), .B1(new_n730), .B2(new_n674), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n731), .A2(KEYINPUT42), .A3(new_n687), .A4(new_n722), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n725), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G131), .ZN(G33));
  NAND4_X1  g548(.A1(new_n722), .A2(new_n313), .A3(new_n508), .A4(new_n662), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G134), .ZN(G36));
  NOR2_X1   g550(.A1(new_n671), .A2(new_n612), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n620), .A2(new_n627), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT43), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n739), .A2(KEYINPUT106), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n739), .A2(KEYINPUT106), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n738), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n742), .B1(new_n738), .B2(new_n741), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n737), .A2(new_n743), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n744), .A2(KEYINPUT44), .ZN(new_n745));
  INV_X1    g559(.A(new_n373), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n375), .A2(new_n376), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n747), .A2(KEYINPUT45), .ZN(new_n748));
  OAI21_X1  g562(.A(G469), .B1(new_n747), .B2(KEYINPUT45), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(new_n378), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT46), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n746), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n751), .A2(KEYINPUT46), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n384), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n666), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n719), .A2(new_n721), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n744), .A2(KEYINPUT44), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n745), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G137), .ZN(G39));
  XNOR2_X1  g577(.A(new_n756), .B(KEYINPUT47), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n547), .A2(new_n556), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n627), .B1(new_n765), .B2(new_n617), .ZN(new_n766));
  INV_X1    g580(.A(new_n661), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR4_X1   g582(.A1(new_n759), .A2(new_n313), .A3(new_n508), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n764), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G140), .ZN(G42));
  NAND2_X1  g585(.A1(new_n743), .A2(new_n562), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n681), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n774), .A2(new_n709), .A3(new_n390), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n773), .A2(new_n708), .A3(new_n775), .ZN(new_n776));
  XOR2_X1   g590(.A(new_n776), .B(KEYINPUT50), .Z(new_n777));
  AND3_X1   g591(.A1(new_n773), .A2(new_n708), .A3(new_n758), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n693), .A2(new_n385), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n778), .B1(new_n764), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n758), .A2(new_n709), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n772), .A2(new_n781), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n651), .A2(new_n714), .ZN(new_n783));
  NOR4_X1   g597(.A1(new_n781), .A2(new_n726), .A3(new_n656), .A4(new_n680), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n620), .A2(new_n628), .ZN(new_n785));
  AOI22_X1  g599(.A1(new_n782), .A2(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n777), .A2(new_n780), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(KEYINPUT51), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT51), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n777), .A2(new_n780), .A3(new_n789), .A4(new_n786), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n773), .A2(new_n703), .A3(new_n708), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(KEYINPUT111), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n561), .B1(new_n784), .B2(new_n766), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n782), .A2(KEYINPUT48), .A3(new_n731), .ZN(new_n797));
  INV_X1    g611(.A(new_n731), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n772), .A2(new_n798), .A3(new_n781), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n799), .A2(KEYINPUT48), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n796), .A2(new_n797), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n794), .B1(new_n793), .B2(new_n795), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n791), .A2(new_n803), .A3(KEYINPUT113), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT113), .B1(new_n791), .B2(new_n803), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n620), .A2(KEYINPUT108), .A3(new_n604), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT108), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n807), .B1(new_n560), .B2(new_n635), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n616), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n809), .A2(new_n810), .A3(new_n612), .A4(new_n609), .ZN(new_n811));
  OAI21_X1  g625(.A(KEYINPUT107), .B1(new_n616), .B2(new_n629), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT107), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n766), .A2(new_n813), .A3(new_n438), .A4(new_n567), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n812), .A2(new_n609), .A3(new_n612), .A4(new_n814), .ZN(new_n815));
  AND4_X1   g629(.A1(new_n607), .A2(new_n811), .A3(new_n704), .A4(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n439), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n617), .B(new_n604), .C1(new_n618), .C2(new_n619), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT80), .B1(new_n380), .B2(new_n385), .ZN(new_n819));
  NOR4_X1   g633(.A1(new_n817), .A2(new_n818), .A3(new_n819), .A4(new_n661), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n820), .A2(new_n313), .A3(new_n651), .A4(new_n758), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n722), .A2(new_n651), .A3(new_n687), .A4(new_n714), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n821), .A2(new_n735), .A3(new_n822), .ZN(new_n823));
  AND4_X1   g637(.A1(new_n652), .A2(new_n697), .A3(new_n700), .A4(new_n711), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n816), .A2(new_n823), .A3(new_n733), .A4(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n647), .A2(new_n386), .A3(new_n661), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n680), .A2(new_n710), .A3(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n663), .A2(new_n688), .A3(new_n715), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT52), .ZN(new_n831));
  AOI22_X1  g645(.A1(new_n730), .A2(new_n674), .B1(new_n649), .B2(new_n650), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n388), .A2(new_n438), .A3(new_n439), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n833), .A2(new_n636), .A3(new_n661), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n768), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n832), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n836), .A2(new_n837), .A3(new_n715), .A4(new_n829), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n831), .A2(KEYINPUT110), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT110), .B1(new_n831), .B2(new_n838), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n827), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n831), .A2(new_n838), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT109), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n825), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n821), .A2(new_n735), .A3(new_n822), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n848), .B1(new_n725), .B2(new_n732), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n811), .A2(new_n815), .A3(new_n607), .A4(new_n704), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n652), .A2(new_n697), .A3(new_n700), .A4(new_n711), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n849), .A2(KEYINPUT109), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n845), .B1(new_n847), .B2(new_n853), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n843), .B(new_n844), .C1(new_n854), .C2(KEYINPUT53), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n825), .A2(new_n846), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT109), .B1(new_n849), .B2(new_n852), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n826), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n840), .A2(new_n842), .ZN(new_n859));
  OAI22_X1  g673(.A1(new_n858), .A2(new_n859), .B1(new_n854), .B2(new_n826), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n855), .B1(new_n860), .B2(new_n844), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n804), .A2(new_n805), .A3(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(G952), .A2(G953), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n693), .A2(KEYINPUT49), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n693), .A2(KEYINPUT49), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n385), .A2(new_n389), .ZN(new_n866));
  NOR4_X1   g680(.A1(new_n726), .A2(new_n864), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n867), .A2(new_n774), .A3(new_n738), .ZN(new_n868));
  OAI22_X1  g682(.A1(new_n862), .A2(new_n863), .B1(new_n680), .B2(new_n868), .ZN(G75));
  OAI21_X1  g683(.A(new_n843), .B1(new_n854), .B2(KEYINPUT53), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n870), .A2(G210), .A3(G902), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT56), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n427), .A2(new_n430), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(new_n428), .ZN(new_n875));
  XOR2_X1   g689(.A(KEYINPUT114), .B(KEYINPUT55), .Z(new_n876));
  XNOR2_X1  g690(.A(new_n875), .B(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n357), .A2(G952), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT116), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT117), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  XOR2_X1   g696(.A(KEYINPUT115), .B(KEYINPUT56), .Z(new_n883));
  NOR2_X1   g697(.A1(new_n877), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n882), .B1(new_n871), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n878), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT118), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n886), .B(new_n887), .ZN(G51));
  NAND2_X1  g702(.A1(new_n870), .A2(KEYINPUT54), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n855), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n378), .B(KEYINPUT57), .Z(new_n892));
  OAI22_X1  g706(.A1(new_n891), .A2(new_n892), .B1(new_n372), .B2(new_n362), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n849), .A2(KEYINPUT53), .A3(new_n852), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n894), .A2(new_n839), .A3(new_n841), .ZN(new_n895));
  INV_X1    g709(.A(new_n845), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n896), .B1(new_n856), .B2(new_n857), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n895), .B1(new_n897), .B2(new_n826), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n898), .A2(new_n315), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n750), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n880), .B1(new_n893), .B2(new_n900), .ZN(G54));
  NAND4_X1  g715(.A1(new_n899), .A2(KEYINPUT58), .A3(G475), .A4(new_n553), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT119), .ZN(new_n903));
  OR2_X1    g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n902), .A2(new_n903), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n899), .A2(KEYINPUT58), .A3(G475), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n880), .B1(new_n906), .B2(new_n544), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n904), .A2(new_n905), .A3(new_n907), .ZN(G60));
  NAND2_X1  g722(.A1(new_n624), .A2(new_n625), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT120), .Z(new_n910));
  XOR2_X1   g724(.A(new_n622), .B(KEYINPUT59), .Z(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n882), .B1(new_n890), .B2(new_n913), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n861), .A2(new_n911), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n914), .B1(new_n915), .B2(new_n910), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(KEYINPUT121), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT121), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n918), .B(new_n914), .C1(new_n915), .C2(new_n910), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n917), .A2(new_n919), .ZN(G63));
  INV_X1    g734(.A(KEYINPUT123), .ZN(new_n921));
  XNOR2_X1  g735(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n922));
  NAND2_X1  g736(.A1(G217), .A2(G902), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n922), .B(new_n923), .Z(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n921), .B1(new_n898), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n870), .A2(KEYINPUT123), .A3(new_n924), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n926), .A2(new_n495), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n926), .A2(new_n927), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n882), .B1(new_n929), .B2(new_n642), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT124), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n931), .B1(new_n929), .B2(new_n642), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n928), .B(new_n930), .C1(new_n932), .C2(KEYINPUT61), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n870), .A2(KEYINPUT123), .A3(new_n924), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT123), .B1(new_n870), .B2(new_n924), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n642), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT61), .B1(new_n936), .B2(KEYINPUT124), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n936), .A2(new_n881), .A3(new_n928), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n933), .A2(new_n939), .ZN(G66));
  OAI21_X1  g754(.A(G953), .B1(new_n396), .B2(new_n565), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n941), .B1(new_n852), .B2(G953), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n874), .B1(G898), .B2(new_n357), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(G69));
  NAND2_X1  g758(.A1(new_n836), .A2(new_n715), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n945), .B1(new_n670), .B2(new_n684), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT62), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n762), .A2(new_n770), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n668), .B1(new_n766), .B2(new_n809), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n950), .A2(new_n798), .A3(new_n759), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n948), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n946), .A2(new_n947), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n357), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n275), .A2(new_n276), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(new_n530), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT125), .ZN(new_n960));
  INV_X1    g774(.A(new_n949), .ZN(new_n961));
  INV_X1    g775(.A(new_n710), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n757), .A2(new_n798), .A3(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n735), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n963), .A2(new_n945), .A3(new_n964), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n961), .A2(KEYINPUT126), .A3(new_n733), .A4(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT126), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n965), .A2(new_n733), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n967), .B1(new_n968), .B2(new_n949), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n966), .A2(new_n969), .A3(new_n357), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n958), .B1(G900), .B2(G953), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n959), .A2(new_n960), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n357), .B1(G227), .B2(G900), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(G72));
  NAND3_X1  g789(.A1(new_n966), .A2(new_n969), .A3(new_n852), .ZN(new_n976));
  NAND2_X1  g790(.A1(G472), .A2(G902), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT63), .Z(new_n978));
  AOI211_X1 g792(.A(new_n256), .B(new_n278), .C1(new_n976), .C2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n978), .ZN(new_n980));
  INV_X1    g794(.A(new_n298), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n981), .A2(KEYINPUT127), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(new_n279), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n860), .A2(new_n980), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n278), .A2(new_n256), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n952), .A2(new_n852), .A3(new_n954), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n985), .B1(new_n986), .B2(new_n978), .ZN(new_n987));
  NOR4_X1   g801(.A1(new_n979), .A2(new_n880), .A3(new_n984), .A4(new_n987), .ZN(G57));
endmodule


