//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 1 1 0 0 0 1 1 1 1 1 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1250, new_n1251,
    new_n1252;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n207));
  INV_X1    g0007(.A(G58), .ZN(new_n208));
  INV_X1    g0008(.A(G232), .ZN(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n206), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n206), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT0), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(G50), .B1(G58), .B2(G68), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(new_n219), .A2(new_n220), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n226), .B1(new_n220), .B2(new_n219), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n217), .A2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G226), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n234), .B(new_n235), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  INV_X1    g0037(.A(G107), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n238), .A2(G97), .ZN(new_n239));
  INV_X1    g0039(.A(G97), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G107), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n202), .A2(G68), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n210), .A2(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n244), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(KEYINPUT18), .ZN(new_n251));
  INV_X1    g0051(.A(G13), .ZN(new_n252));
  NOR3_X1   g0052(.A1(new_n252), .A2(new_n222), .A3(G1), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n221), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n258), .B1(new_n259), .B2(G20), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n256), .B1(new_n260), .B2(new_n255), .ZN(new_n261));
  XOR2_X1   g0061(.A(new_n261), .B(KEYINPUT74), .Z(new_n262));
  XOR2_X1   g0062(.A(KEYINPUT71), .B(KEYINPUT16), .Z(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT3), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G33), .ZN(new_n268));
  AOI21_X1  g0068(.A(G20), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(KEYINPUT72), .B1(new_n269), .B2(KEYINPUT7), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT72), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT7), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT3), .B(G33), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n271), .B(new_n272), .C1(new_n273), .C2(G20), .ZN(new_n274));
  OR3_X1    g0074(.A1(new_n267), .A2(KEYINPUT73), .A3(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n266), .A2(KEYINPUT73), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(new_n276), .A3(new_n268), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n272), .A2(G20), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n270), .A2(new_n274), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(new_n210), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n208), .A2(new_n210), .ZN(new_n281));
  OAI21_X1  g0081(.A(G20), .B1(new_n281), .B2(new_n201), .ZN(new_n282));
  INV_X1    g0082(.A(G159), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G20), .A2(G33), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n282), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n264), .B1(new_n280), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n258), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n272), .B1(new_n273), .B2(G20), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n266), .A2(new_n268), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(KEYINPUT7), .A3(new_n222), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n286), .B1(new_n292), .B2(G68), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n288), .B1(new_n293), .B2(KEYINPUT16), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n262), .B1(new_n287), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n259), .B1(G41), .B2(G45), .ZN(new_n296));
  INV_X1    g0096(.A(G274), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(G33), .A2(G41), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n300), .A2(G1), .A3(G13), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n296), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n299), .B1(new_n302), .B2(new_n209), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n273), .A2(G226), .A3(G1698), .ZN(new_n304));
  INV_X1    g0104(.A(G87), .ZN(new_n305));
  INV_X1    g0105(.A(G1698), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n273), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G223), .ZN(new_n308));
  OAI221_X1 g0108(.A(new_n304), .B1(new_n265), .B2(new_n305), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n301), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n303), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n311), .A2(G179), .ZN(new_n312));
  INV_X1    g0112(.A(G169), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n251), .B1(new_n295), .B2(new_n315), .ZN(new_n316));
  NOR3_X1   g0116(.A1(new_n295), .A2(new_n315), .A3(new_n251), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n316), .B1(new_n317), .B2(KEYINPUT75), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT75), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n319), .B(new_n251), .C1(new_n295), .C2(new_n315), .ZN(new_n320));
  INV_X1    g0120(.A(G200), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n311), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n322), .B1(G190), .B2(new_n311), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n295), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT17), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT17), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n295), .A2(new_n323), .A3(new_n326), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n318), .A2(new_n320), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  XOR2_X1   g0128(.A(KEYINPUT8), .B(G58), .Z(new_n329));
  NOR2_X1   g0129(.A1(new_n265), .A2(G20), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n329), .A2(new_n330), .B1(G150), .B2(new_n284), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n203), .A2(G20), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n288), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n253), .A2(new_n202), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n288), .B1(G1), .B2(new_n222), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n334), .B1(new_n335), .B2(new_n202), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  OR2_X1    g0137(.A1(new_n337), .A2(KEYINPUT9), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(KEYINPUT9), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT10), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n338), .B(new_n339), .C1(KEYINPUT66), .C2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n273), .A2(G222), .A3(new_n306), .ZN(new_n342));
  INV_X1    g0142(.A(G77), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n273), .A2(G1698), .ZN(new_n344));
  OAI221_X1 g0144(.A(new_n342), .B1(new_n343), .B2(new_n273), .C1(new_n344), .C2(new_n308), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n310), .ZN(new_n346));
  INV_X1    g0146(.A(new_n302), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n298), .B1(new_n347), .B2(G226), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G200), .ZN(new_n350));
  INV_X1    g0150(.A(G190), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n350), .B1(new_n351), .B2(new_n349), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n341), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT66), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n353), .B1(new_n354), .B2(KEYINPUT10), .ZN(new_n355));
  OAI211_X1 g0155(.A(KEYINPUT66), .B(new_n340), .C1(new_n341), .C2(new_n352), .ZN(new_n356));
  INV_X1    g0156(.A(new_n337), .ZN(new_n357));
  INV_X1    g0157(.A(new_n349), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n357), .B1(new_n358), .B2(G169), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n349), .A2(G179), .ZN(new_n360));
  OR2_X1    g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n355), .A2(new_n356), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n253), .A2(new_n343), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n335), .B2(new_n343), .ZN(new_n365));
  OAI22_X1  g0165(.A1(new_n255), .A2(new_n285), .B1(new_n222), .B2(new_n343), .ZN(new_n366));
  XOR2_X1   g0166(.A(KEYINPUT15), .B(G87), .Z(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n330), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n366), .B1(KEYINPUT65), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(KEYINPUT65), .B2(new_n368), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n365), .B1(new_n370), .B2(new_n258), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n290), .A2(G107), .ZN(new_n372));
  OAI221_X1 g0172(.A(new_n372), .B1(new_n344), .B2(new_n211), .C1(new_n209), .C2(new_n307), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n310), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n298), .B1(new_n347), .B2(G244), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n371), .B1(new_n313), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G179), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n374), .A2(new_n378), .A3(new_n375), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n376), .A2(G200), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n381), .B(new_n371), .C1(new_n351), .C2(new_n376), .ZN(new_n382));
  AND4_X1   g0182(.A1(new_n328), .A2(new_n363), .A3(new_n380), .A4(new_n382), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n266), .A2(new_n268), .A3(G232), .A4(G1698), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n266), .A2(new_n268), .A3(G226), .A4(new_n306), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n265), .A2(new_n240), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n310), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT67), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n302), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n301), .A2(KEYINPUT67), .A3(new_n296), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n391), .A2(G238), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n389), .A2(new_n393), .A3(new_n299), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT13), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT13), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n389), .A2(new_n393), .A3(new_n396), .A4(new_n299), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT68), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT68), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n399), .B1(new_n394), .B2(KEYINPUT13), .ZN(new_n400));
  OAI21_X1  g0200(.A(G169), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT14), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT14), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n403), .B(G169), .C1(new_n398), .C2(new_n400), .ZN(new_n404));
  AND3_X1   g0204(.A1(new_n395), .A2(G179), .A3(new_n397), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n402), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT70), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n405), .B1(new_n401), .B2(KEYINPUT14), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT70), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(new_n410), .A3(new_n404), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT69), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n285), .B2(new_n202), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n284), .A2(KEYINPUT69), .A3(G50), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n330), .A2(G77), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n210), .A2(G20), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n414), .A2(new_n415), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n418), .A2(new_n258), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT11), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT12), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n421), .B1(new_n253), .B2(new_n210), .ZN(new_n422));
  NOR3_X1   g0222(.A1(new_n254), .A2(KEYINPUT12), .A3(G68), .ZN(new_n423));
  OAI221_X1 g0223(.A(new_n420), .B1(new_n210), .B2(new_n335), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n419), .A2(KEYINPUT11), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(G200), .B1(new_n398), .B2(new_n400), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n395), .A2(new_n397), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n427), .B1(G190), .B2(new_n429), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n412), .A2(new_n427), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n383), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n273), .A2(G257), .A3(new_n306), .ZN(new_n433));
  INV_X1    g0233(.A(G303), .ZN(new_n434));
  INV_X1    g0234(.A(G264), .ZN(new_n435));
  OAI221_X1 g0235(.A(new_n433), .B1(new_n434), .B2(new_n273), .C1(new_n344), .C2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n310), .ZN(new_n437));
  INV_X1    g0237(.A(G41), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n259), .B(G45), .C1(new_n438), .C2(KEYINPUT5), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n438), .A2(KEYINPUT5), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n441), .A2(new_n310), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n442), .A2(G270), .B1(G274), .B2(new_n441), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n313), .B1(new_n437), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n254), .A2(G116), .ZN(new_n445));
  AOI211_X1 g0245(.A(new_n258), .B(new_n253), .C1(new_n259), .C2(G33), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n445), .B1(new_n446), .B2(G116), .ZN(new_n447));
  NAND2_X1  g0247(.A1(G33), .A2(G283), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n448), .B(new_n222), .C1(G33), .C2(new_n240), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n449), .B(new_n258), .C1(new_n222), .C2(G116), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT20), .ZN(new_n451));
  XNOR2_X1  g0251(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n447), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n444), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT21), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n444), .A2(KEYINPUT21), .A3(new_n453), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n453), .A2(G179), .A3(new_n437), .A4(new_n443), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(KEYINPUT25), .B1(new_n253), .B2(new_n238), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n253), .A2(KEYINPUT25), .A3(new_n238), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n446), .A2(G107), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g0263(.A1(KEYINPUT81), .A2(G87), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n266), .A2(new_n268), .A3(new_n464), .A4(new_n222), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT22), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n273), .A2(KEYINPUT22), .A3(new_n222), .A4(new_n464), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT23), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n469), .B1(new_n222), .B2(G107), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n238), .A2(KEYINPUT23), .A3(G20), .ZN(new_n471));
  AND2_X1   g0271(.A1(G33), .A2(G116), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n470), .A2(new_n471), .B1(new_n222), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n467), .A2(new_n468), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT24), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT82), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n474), .A2(KEYINPUT82), .A3(KEYINPUT24), .ZN(new_n478));
  OR2_X1    g0278(.A1(new_n474), .A2(KEYINPUT24), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n480), .A2(KEYINPUT83), .A3(new_n258), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT83), .B1(new_n480), .B2(new_n258), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n463), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n273), .A2(G250), .A3(new_n306), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n273), .A2(G257), .A3(G1698), .ZN(new_n485));
  INV_X1    g0285(.A(G294), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n484), .B(new_n485), .C1(new_n265), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n310), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n442), .A2(G264), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n441), .A2(G274), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(new_n378), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n492), .B1(G169), .B2(new_n491), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n459), .B1(new_n483), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n463), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT83), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n474), .A2(KEYINPUT82), .A3(KEYINPUT24), .ZN(new_n498));
  AOI21_X1  g0298(.A(KEYINPUT82), .B1(new_n474), .B2(KEYINPUT24), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n474), .A2(KEYINPUT24), .ZN(new_n500));
  NOR3_X1   g0300(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n497), .B1(new_n501), .B2(new_n288), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n480), .A2(KEYINPUT83), .A3(new_n258), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n496), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n491), .A2(new_n351), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n505), .B1(G200), .B2(new_n491), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n254), .A2(G97), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n508), .B1(new_n446), .B2(G97), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n240), .A2(G107), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT6), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT76), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT76), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n511), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  XNOR2_X1  g0316(.A(KEYINPUT76), .B(KEYINPUT6), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n516), .B1(new_n242), .B2(new_n517), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n518), .A2(G20), .B1(G77), .B2(new_n284), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(new_n279), .B2(new_n238), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n510), .B1(new_n258), .B2(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(G257), .B(new_n301), .C1(new_n439), .C2(new_n440), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n490), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n266), .A2(new_n268), .A3(G244), .A4(new_n306), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT4), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n273), .A2(KEYINPUT4), .A3(G244), .A4(new_n306), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n273), .A2(G250), .A3(G1698), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n526), .A2(new_n527), .A3(new_n448), .A4(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n523), .B1(new_n529), .B2(new_n310), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G190), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n310), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n532), .A2(new_n490), .A3(new_n522), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n533), .A2(KEYINPUT77), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT77), .ZN(new_n535));
  OAI21_X1  g0335(.A(G200), .B1(new_n530), .B2(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n521), .B(new_n531), .C1(new_n534), .C2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n518), .A2(G20), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n284), .A2(G77), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n270), .A2(new_n274), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n277), .A2(new_n278), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n540), .B1(new_n543), .B2(G107), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n509), .B1(new_n544), .B2(new_n288), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT78), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n533), .B2(G179), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n530), .A2(G169), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n530), .A2(KEYINPUT78), .A3(new_n378), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n545), .A2(new_n547), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n266), .A2(new_n268), .A3(G244), .A4(G1698), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n266), .A2(new_n268), .A3(G238), .A4(new_n306), .ZN(new_n553));
  INV_X1    g0353(.A(G116), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n552), .B(new_n553), .C1(new_n265), .C2(new_n554), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n555), .A2(new_n310), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n259), .A2(G45), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n557), .A2(new_n297), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n301), .A2(G250), .A3(new_n557), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n558), .B1(new_n559), .B2(KEYINPUT79), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT79), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n301), .A2(new_n561), .A3(G250), .A4(new_n557), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(G200), .B1(new_n556), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n273), .A2(new_n222), .A3(G68), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n330), .A2(G97), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT19), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT80), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT80), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(KEYINPUT19), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g0372(.A(KEYINPUT80), .B(KEYINPUT19), .ZN(new_n573));
  AOI21_X1  g0373(.A(G20), .B1(new_n573), .B2(new_n386), .ZN(new_n574));
  NOR3_X1   g0374(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n565), .B(new_n572), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n367), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n576), .A2(new_n258), .B1(new_n253), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n555), .A2(new_n310), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n579), .A2(G190), .A3(new_n562), .A4(new_n560), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n446), .A2(G87), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n564), .A2(new_n578), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n313), .B1(new_n556), .B2(new_n563), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n446), .A2(new_n367), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n565), .A2(new_n572), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n386), .A2(new_n568), .A3(new_n570), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n575), .B1(new_n586), .B2(new_n222), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n258), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n577), .A2(new_n253), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n584), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n579), .A2(new_n378), .A3(new_n562), .A4(new_n560), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n583), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n582), .A2(new_n592), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n537), .A2(new_n551), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n437), .A2(new_n443), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n453), .B1(new_n595), .B2(G200), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n351), .B2(new_n595), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n495), .A2(new_n507), .A3(new_n594), .A4(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n432), .A2(new_n598), .ZN(G372));
  INV_X1    g0399(.A(new_n361), .ZN(new_n600));
  INV_X1    g0400(.A(new_n317), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n316), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n426), .B1(new_n408), .B2(new_n411), .ZN(new_n603));
  INV_X1    g0403(.A(new_n380), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n430), .A2(new_n428), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n325), .A2(new_n327), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n602), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n355), .A2(new_n356), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n600), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT26), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n582), .A2(new_n592), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n612), .B1(new_n551), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n521), .A2(new_n548), .ZN(new_n615));
  INV_X1    g0415(.A(new_n550), .ZN(new_n616));
  AOI21_X1  g0416(.A(KEYINPUT78), .B1(new_n530), .B2(new_n378), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n593), .A2(new_n615), .A3(KEYINPUT26), .A4(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(KEYINPUT85), .B1(new_n620), .B2(new_n592), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT85), .ZN(new_n622));
  INV_X1    g0422(.A(new_n592), .ZN(new_n623));
  AOI211_X1 g0423(.A(new_n622), .B(new_n623), .C1(new_n614), .C2(new_n619), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n457), .A2(new_n458), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT21), .B1(new_n444), .B2(new_n453), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n628), .B1(new_n504), .B2(new_n493), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT84), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n537), .A2(new_n551), .A3(new_n593), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n504), .B2(new_n506), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n483), .A2(new_n494), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT84), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(new_n634), .A3(new_n628), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n630), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n625), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n611), .B1(new_n432), .B2(new_n637), .ZN(G369));
  NOR2_X1   g0438(.A1(new_n252), .A2(G20), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n259), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n640), .A2(KEYINPUT27), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(KEYINPUT27), .ZN(new_n642));
  INV_X1    g0442(.A(G213), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(G343), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n453), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n628), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n597), .ZN(new_n649));
  INV_X1    g0449(.A(G330), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n633), .A2(new_n507), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n504), .A2(new_n645), .ZN(new_n653));
  OAI22_X1  g0453(.A1(new_n652), .A2(new_n653), .B1(new_n633), .B2(new_n645), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n633), .ZN(new_n656));
  XOR2_X1   g0456(.A(new_n645), .B(KEYINPUT86), .Z(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n459), .A2(new_n645), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n661), .A2(new_n507), .A3(new_n633), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n655), .A2(new_n659), .A3(new_n662), .ZN(G399));
  INV_X1    g0463(.A(KEYINPUT29), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n623), .B1(new_n614), .B2(new_n619), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n594), .A2(new_n507), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n665), .B1(new_n666), .B2(new_n495), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n664), .B1(new_n667), .B2(new_n645), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n665), .B(KEYINPUT85), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n630), .A2(new_n632), .A3(new_n635), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n657), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n668), .B1(new_n671), .B2(new_n664), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n595), .A2(new_n378), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n488), .A2(new_n489), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n556), .A2(new_n563), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n673), .A2(new_n674), .A3(new_n530), .A4(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT30), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n674), .A2(new_n675), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n679), .A2(KEYINPUT30), .A3(new_n530), .A4(new_n673), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n595), .A2(new_n378), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(new_n675), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n682), .A2(new_n491), .A3(new_n533), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n678), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n684), .A2(KEYINPUT31), .A3(new_n657), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n646), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT31), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI211_X1 g0488(.A(new_n685), .B(new_n688), .C1(new_n598), .C2(new_n657), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G330), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n672), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n259), .ZN(new_n692));
  INV_X1    g0492(.A(new_n218), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(G41), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n575), .A2(new_n554), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n694), .A2(new_n695), .A3(new_n259), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n696), .B1(new_n225), .B2(new_n694), .ZN(new_n697));
  XOR2_X1   g0497(.A(new_n697), .B(KEYINPUT28), .Z(new_n698));
  NAND2_X1  g0498(.A1(new_n692), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT87), .Z(G364));
  AOI21_X1  g0500(.A(new_n222), .B1(KEYINPUT89), .B2(new_n313), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n313), .A2(KEYINPUT89), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n221), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n222), .A2(new_n351), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n378), .A2(G200), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(G322), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n290), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n321), .A2(G179), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n704), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n222), .A2(G190), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n705), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  AOI22_X1  g0514(.A1(G303), .A2(new_n711), .B1(new_n714), .B2(G311), .ZN(new_n715));
  INV_X1    g0515(.A(G283), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n712), .A2(new_n709), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n378), .A2(new_n321), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n712), .ZN(new_n719));
  XOR2_X1   g0519(.A(KEYINPUT33), .B(G317), .Z(new_n720));
  OAI221_X1 g0520(.A(new_n715), .B1(new_n716), .B2(new_n717), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n378), .A2(new_n321), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT90), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n712), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  AOI211_X1 g0525(.A(new_n708), .B(new_n721), .C1(G329), .C2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n704), .A2(new_n718), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G326), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n723), .A2(G190), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G20), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n729), .B1(new_n732), .B2(new_n486), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n733), .A2(KEYINPUT92), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(KEYINPUT92), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n726), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT93), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n719), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n731), .A2(G97), .B1(G68), .B2(new_n739), .ZN(new_n740));
  XOR2_X1   g0540(.A(new_n740), .B(KEYINPUT91), .Z(new_n741));
  OAI21_X1  g0541(.A(new_n273), .B1(new_n717), .B2(new_n238), .ZN(new_n742));
  AOI22_X1  g0542(.A1(new_n728), .A2(G50), .B1(new_n714), .B2(G77), .ZN(new_n743));
  OAI221_X1 g0543(.A(new_n743), .B1(new_n208), .B2(new_n706), .C1(new_n305), .C2(new_n710), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n725), .A2(G159), .ZN(new_n745));
  AOI211_X1 g0545(.A(new_n742), .B(new_n744), .C1(KEYINPUT32), .C2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(KEYINPUT32), .B2(new_n745), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n738), .B1(new_n741), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n736), .A2(new_n737), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n703), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n259), .B1(new_n639), .B2(G45), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n694), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n273), .A2(G355), .A3(new_n218), .ZN(new_n755));
  INV_X1    g0555(.A(G45), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n249), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n693), .A2(new_n273), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(G45), .B2(new_n224), .ZN(new_n759));
  OAI221_X1 g0559(.A(new_n755), .B1(G116), .B2(new_n218), .C1(new_n757), .C2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G13), .A2(G33), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n703), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n754), .B1(new_n760), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n649), .ZN(new_n766));
  INV_X1    g0566(.A(new_n763), .ZN(new_n767));
  OAI211_X1 g0567(.A(new_n750), .B(new_n765), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n651), .A2(KEYINPUT88), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n766), .A2(G330), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n753), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n770), .A2(new_n772), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n768), .B1(new_n774), .B2(new_n775), .ZN(G396));
  NOR2_X1   g0576(.A1(new_n380), .A2(new_n646), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n371), .A2(new_n645), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n382), .A2(new_n778), .B1(new_n377), .B2(new_n379), .ZN(new_n779));
  OR3_X1    g0579(.A1(new_n777), .A2(new_n779), .A3(KEYINPUT97), .ZN(new_n780));
  OAI21_X1  g0580(.A(KEYINPUT97), .B1(new_n777), .B2(new_n779), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n671), .B(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n690), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n753), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(new_n785), .B2(new_n784), .ZN(new_n787));
  INV_X1    g0587(.A(new_n703), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n762), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT94), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n753), .B1(new_n790), .B2(G77), .ZN(new_n791));
  INV_X1    g0591(.A(new_n717), .ZN(new_n792));
  AOI22_X1  g0592(.A1(G87), .A2(new_n792), .B1(new_n714), .B2(G116), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n793), .B1(new_n238), .B2(new_n710), .C1(new_n434), .C2(new_n727), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n290), .B1(new_n719), .B2(new_n716), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n732), .A2(new_n240), .B1(new_n486), .B2(new_n706), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT95), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G311), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n796), .B(new_n799), .C1(new_n800), .C2(new_n724), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n797), .A2(new_n798), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n273), .B1(new_n717), .B2(new_n210), .C1(new_n202), .C2(new_n710), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(new_n725), .B2(G132), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n208), .B2(new_n732), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n728), .A2(G137), .B1(new_n714), .B2(G159), .ZN(new_n806));
  INV_X1    g0606(.A(G143), .ZN(new_n807));
  INV_X1    g0607(.A(G150), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n806), .B1(new_n807), .B2(new_n706), .C1(new_n808), .C2(new_n719), .ZN(new_n809));
  XNOR2_X1  g0609(.A(KEYINPUT96), .B(KEYINPUT34), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n809), .B(new_n810), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n801), .A2(new_n802), .B1(new_n805), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n791), .B1(new_n812), .B2(new_n703), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n782), .B2(new_n762), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n787), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(G384));
  AND4_X1   g0616(.A1(new_n410), .A2(new_n402), .A3(new_n404), .A4(new_n406), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n410), .B1(new_n409), .B2(new_n404), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n427), .B(new_n646), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(KEYINPUT99), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT99), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n412), .A2(new_n821), .A3(new_n427), .A4(new_n646), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n427), .A2(new_n646), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n431), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n658), .B(new_n782), .C1(new_n625), .C2(new_n636), .ZN(new_n827));
  INV_X1    g0627(.A(new_n777), .ZN(new_n828));
  AND3_X1   g0628(.A1(new_n827), .A2(KEYINPUT98), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(KEYINPUT98), .B1(new_n827), .B2(new_n828), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n826), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT100), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n827), .A2(new_n828), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT98), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n827), .A2(KEYINPUT98), .A3(new_n828), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n838), .A2(KEYINPUT100), .A3(new_n826), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n294), .B1(new_n263), .B2(new_n293), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT101), .ZN(new_n841));
  AND3_X1   g0641(.A1(new_n840), .A2(new_n841), .A3(new_n261), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n841), .B1(new_n840), .B2(new_n261), .ZN(new_n843));
  NOR3_X1   g0643(.A1(new_n312), .A2(new_n314), .A3(new_n644), .ZN(new_n844));
  NOR3_X1   g0644(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n324), .ZN(new_n846));
  OAI21_X1  g0646(.A(KEYINPUT37), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OR2_X1    g0647(.A1(new_n844), .A2(new_n295), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT37), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n848), .A2(new_n849), .A3(new_n324), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n842), .A2(new_n843), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n644), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n851), .B1(new_n328), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT38), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n851), .B(KEYINPUT38), .C1(new_n328), .C2(new_n853), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n833), .A2(new_n839), .A3(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n602), .A2(new_n644), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n858), .A2(KEYINPUT39), .ZN(new_n861));
  INV_X1    g0661(.A(new_n850), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n849), .B1(new_n848), .B2(new_n324), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n295), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n644), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n602), .B2(new_n607), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n855), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n857), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n861), .B1(KEYINPUT39), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n603), .A2(new_n645), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n860), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n859), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n672), .A2(new_n432), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n609), .A2(new_n610), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n361), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  XOR2_X1   g0678(.A(new_n874), .B(new_n878), .Z(new_n879));
  NAND3_X1  g0679(.A1(new_n684), .A2(KEYINPUT31), .A3(new_n646), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n688), .B(new_n880), .C1(new_n598), .C2(new_n657), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n383), .A2(G330), .A3(new_n431), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n782), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n883), .B1(new_n825), .B2(new_n823), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n869), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT40), .B1(new_n856), .B2(new_n857), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n885), .A2(KEYINPUT40), .B1(new_n886), .B2(new_n884), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n882), .B1(new_n887), .B2(new_n650), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n383), .A2(new_n431), .A3(new_n881), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n888), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  OAI22_X1  g0690(.A1(new_n879), .A2(new_n890), .B1(new_n259), .B2(new_n639), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n890), .B2(new_n879), .ZN(new_n892));
  OAI211_X1 g0692(.A(G116), .B(new_n223), .C1(new_n518), .C2(KEYINPUT35), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(KEYINPUT35), .B2(new_n518), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT36), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n225), .B(G77), .C1(new_n208), .C2(new_n210), .ZN(new_n896));
  AOI211_X1 g0696(.A(new_n259), .B(G13), .C1(new_n896), .C2(new_n245), .ZN(new_n897));
  OR3_X1    g0697(.A1(new_n892), .A2(new_n895), .A3(new_n897), .ZN(G367));
  AND2_X1   g0698(.A1(new_n656), .A2(new_n537), .ZN(new_n899));
  INV_X1    g0699(.A(new_n551), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n658), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n537), .B(new_n551), .C1(new_n658), .C2(new_n521), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n551), .B2(new_n658), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  OR2_X1    g0704(.A1(new_n904), .A2(new_n662), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT42), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n901), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT102), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n909), .B1(new_n907), .B2(new_n906), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n578), .A2(new_n581), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n646), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n593), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n592), .B2(new_n912), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n910), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(KEYINPUT103), .B(KEYINPUT104), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n920));
  OR3_X1    g0720(.A1(new_n910), .A2(new_n915), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n655), .B2(new_n904), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n662), .B1(new_n654), .B2(new_n661), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n650), .B2(new_n649), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n655), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n691), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n659), .A2(new_n662), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n904), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT44), .Z(new_n930));
  NOR2_X1   g0730(.A1(new_n928), .A2(new_n904), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT45), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n927), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n934), .A2(new_n691), .ZN(new_n935));
  XOR2_X1   g0735(.A(KEYINPUT105), .B(KEYINPUT41), .Z(new_n936));
  XNOR2_X1  g0736(.A(new_n694), .B(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n751), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n655), .A2(new_n904), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n918), .A2(new_n939), .A3(new_n919), .A4(new_n921), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n923), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n273), .B1(new_n714), .B2(G283), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n711), .A2(KEYINPUT46), .A3(G116), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT46), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n710), .B2(new_n554), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n942), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  AOI22_X1  g0746(.A1(G311), .A2(new_n728), .B1(new_n739), .B2(G294), .ZN(new_n947));
  OAI221_X1 g0747(.A(new_n947), .B1(new_n240), .B2(new_n717), .C1(new_n434), .C2(new_n706), .ZN(new_n948));
  AOI211_X1 g0748(.A(new_n946), .B(new_n948), .C1(G317), .C2(new_n725), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n238), .B2(new_n732), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT106), .Z(new_n951));
  OAI22_X1  g0751(.A1(new_n808), .A2(new_n706), .B1(new_n719), .B2(new_n283), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n727), .A2(new_n807), .B1(new_n717), .B2(new_n343), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n273), .B1(new_n713), .B2(new_n202), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n710), .A2(new_n208), .ZN(new_n955));
  NOR4_X1   g0755(.A1(new_n952), .A2(new_n953), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(G137), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n956), .B1(new_n957), .B2(new_n724), .C1(new_n210), .C2(new_n732), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n951), .A2(new_n958), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n959), .A2(KEYINPUT47), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(KEYINPUT47), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n960), .A2(new_n703), .A3(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n758), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n236), .A2(new_n963), .ZN(new_n964));
  AOI211_X1 g0764(.A(new_n763), .B(new_n703), .C1(new_n693), .C2(new_n367), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n754), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n962), .B(new_n966), .C1(new_n767), .C2(new_n914), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n941), .A2(new_n967), .ZN(G387));
  INV_X1    g0768(.A(new_n926), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n752), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT107), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n654), .A2(new_n767), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n728), .A2(G322), .B1(new_n714), .B2(G303), .ZN(new_n973));
  INV_X1    g0773(.A(G317), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n973), .B1(new_n800), .B2(new_n719), .C1(new_n974), .C2(new_n706), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT48), .Z(new_n976));
  OAI22_X1  g0776(.A1(new_n732), .A2(new_n716), .B1(new_n486), .B2(new_n710), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n977), .A2(KEYINPUT109), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n977), .A2(KEYINPUT109), .ZN(new_n979));
  NOR3_X1   g0779(.A1(new_n976), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n980), .A2(KEYINPUT49), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(KEYINPUT49), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n290), .B1(new_n717), .B2(new_n554), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(new_n725), .B2(G326), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n981), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n727), .A2(new_n283), .B1(new_n706), .B2(new_n202), .ZN(new_n986));
  AOI211_X1 g0786(.A(new_n290), .B(new_n986), .C1(G97), .C2(new_n792), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n731), .A2(new_n367), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n725), .A2(G150), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n719), .A2(new_n255), .B1(new_n713), .B2(new_n210), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n710), .A2(new_n343), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n987), .A2(new_n988), .A3(new_n989), .A4(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n788), .B1(new_n985), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n233), .A2(new_n756), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n329), .A2(new_n202), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT50), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  AOI211_X1 g0798(.A(G45), .B(new_n695), .C1(G68), .C2(G77), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n963), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n995), .B1(new_n1001), .B2(KEYINPUT108), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(KEYINPUT108), .B2(new_n1001), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n695), .A2(new_n218), .A3(new_n273), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1003), .B(new_n1004), .C1(G107), .C2(new_n218), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n754), .B(new_n994), .C1(new_n764), .C2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n971), .B1(new_n972), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n969), .B1(new_n690), .B2(new_n672), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n694), .ZN(new_n1009));
  OR3_X1    g0809(.A1(new_n1008), .A2(new_n927), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1007), .A2(new_n1010), .ZN(G393));
  INV_X1    g0811(.A(new_n655), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n933), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT110), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n655), .B1(new_n930), .B2(new_n932), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n691), .B2(new_n926), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n934), .A2(new_n1009), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n904), .A2(new_n763), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n244), .A2(new_n963), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n764), .B1(new_n240), .B2(new_n218), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n753), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n727), .A2(new_n974), .B1(new_n706), .B2(new_n800), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT113), .Z(new_n1025));
  NOR2_X1   g0825(.A1(new_n1025), .A2(KEYINPUT52), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT114), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n725), .A2(G322), .B1(G283), .B2(new_n711), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1025), .A2(KEYINPUT52), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n719), .A2(new_n434), .B1(new_n713), .B2(new_n486), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n273), .B(new_n1032), .C1(G107), .C2(new_n792), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1033), .B1(new_n732), .B2(new_n554), .C1(new_n1028), .C2(new_n1027), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n731), .A2(G77), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n202), .B2(new_n719), .C1(new_n255), .C2(new_n713), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT112), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n727), .A2(new_n808), .B1(new_n706), .B2(new_n283), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT51), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n273), .B1(new_n717), .B2(new_n305), .C1(new_n210), .C2(new_n710), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n725), .B2(G143), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1038), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n1031), .A2(new_n1034), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1023), .B1(new_n1045), .B2(new_n703), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n1018), .A2(new_n1019), .B1(new_n1020), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT111), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n751), .B1(new_n1017), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n1048), .B2(new_n1017), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1047), .A2(new_n1050), .ZN(G390));
  INV_X1    g0851(.A(KEYINPUT117), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n820), .A2(new_n822), .B1(new_n431), .B2(new_n824), .ZN(new_n1053));
  NOR3_X1   g0853(.A1(new_n1053), .A2(new_n650), .A3(new_n883), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n870), .B1(new_n831), .B2(new_n871), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT115), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n782), .A2(new_n667), .A3(new_n645), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n823), .A2(new_n825), .B1(new_n1057), .B2(new_n828), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n869), .A2(new_n871), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1056), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n872), .B1(new_n857), .B2(new_n868), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1057), .A2(new_n828), .ZN(new_n1062));
  OAI211_X1 g0862(.A(KEYINPUT115), .B(new_n1061), .C1(new_n1062), .C2(new_n1053), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1054), .B1(new_n1055), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n689), .A2(G330), .A3(new_n782), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n826), .A2(new_n1067), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n872), .B1(new_n838), .B2(new_n826), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1068), .B(new_n1069), .C1(new_n1070), .C2(new_n870), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n1065), .A2(new_n1071), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n823), .B(new_n825), .C1(new_n883), .C2(new_n650), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1068), .A2(new_n1062), .A3(new_n1073), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n829), .A2(new_n830), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n884), .A2(G330), .B1(new_n1053), .B2(new_n1066), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n611), .B(new_n882), .C1(new_n672), .C2(new_n432), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT116), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1077), .A2(KEYINPUT116), .A3(new_n1079), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1052), .B1(new_n1072), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1009), .B1(new_n1072), .B2(new_n1084), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n826), .A2(new_n1067), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n1054), .A2(new_n1087), .B1(new_n829), .B2(new_n830), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1081), .B(new_n1078), .C1(new_n1088), .C2(new_n1074), .ZN(new_n1089));
  AOI21_X1  g0889(.A(KEYINPUT116), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1065), .A2(new_n1071), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1091), .A2(new_n1092), .A3(KEYINPUT117), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1085), .A2(new_n1086), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1072), .A2(new_n752), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n753), .B1(new_n790), .B2(new_n329), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n706), .A2(new_n554), .B1(new_n717), .B2(new_n210), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n273), .B(new_n1097), .C1(G87), .C2(new_n711), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n725), .A2(G294), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n727), .A2(new_n716), .B1(new_n719), .B2(new_n238), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(G97), .B2(new_n714), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1098), .A2(new_n1035), .A3(new_n1099), .A4(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n290), .B1(new_n792), .B2(G50), .ZN(new_n1103));
  INV_X1    g0903(.A(G128), .ZN(new_n1104));
  INV_X1    g0904(.A(G132), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1103), .B1(new_n1104), .B2(new_n727), .C1(new_n1105), .C2(new_n706), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n710), .A2(new_n808), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT119), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1108), .A2(KEYINPUT53), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1106), .B(new_n1109), .C1(G125), .C2(new_n725), .ZN(new_n1110));
  XOR2_X1   g0910(.A(KEYINPUT54), .B(G143), .Z(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n1112), .A2(new_n713), .B1(new_n957), .B2(new_n719), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n731), .B2(G159), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(KEYINPUT118), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1108), .A2(KEYINPUT53), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1110), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1115), .A2(KEYINPUT118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1102), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1096), .B1(new_n1120), .B2(new_n703), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n870), .B2(new_n762), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1095), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1094), .A2(new_n1124), .ZN(G378));
  INV_X1    g0925(.A(KEYINPUT57), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1078), .B1(new_n1072), .B2(new_n1084), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n357), .A2(new_n644), .ZN(new_n1128));
  XOR2_X1   g0928(.A(new_n362), .B(new_n1128), .Z(new_n1129));
  XNOR2_X1  g0929(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(KEYINPUT122), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n887), .B2(new_n650), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT40), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n884), .B2(new_n869), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n884), .A2(new_n886), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1135), .B(G330), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n859), .A2(new_n1137), .A3(new_n873), .A4(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n859), .A2(new_n873), .B1(new_n1137), .B2(new_n1141), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1126), .B1(new_n1127), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1079), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1137), .A2(new_n1141), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n874), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n1142), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1147), .A2(KEYINPUT57), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1146), .A2(new_n694), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n792), .A2(G58), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n1153), .B1(new_n238), .B2(new_n706), .C1(new_n577), .C2(new_n713), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n290), .A2(new_n438), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n727), .A2(new_n554), .B1(new_n719), .B2(new_n240), .ZN(new_n1156));
  NOR4_X1   g0956(.A1(new_n1154), .A2(new_n991), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1157), .B1(new_n210), .B2(new_n732), .C1(new_n716), .C2(new_n724), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT58), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1155), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(G132), .A2(new_n739), .B1(new_n711), .B2(new_n1111), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n706), .A2(new_n1104), .B1(new_n713), .B2(new_n957), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(G125), .B2(new_n728), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1164), .B(new_n1166), .C1(new_n732), .C2(new_n808), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT120), .Z(new_n1168));
  OR2_X1    g0968(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1169));
  AOI211_X1 g0969(.A(G33), .B(G41), .C1(new_n792), .C2(G159), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT121), .B(G124), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1170), .B1(new_n724), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n1168), .B2(KEYINPUT59), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1160), .B(new_n1163), .C1(new_n1169), .C2(new_n1173), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n753), .B1(G50), .B2(new_n790), .C1(new_n1174), .C2(new_n788), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n1134), .B2(new_n761), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n1150), .B2(new_n752), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1152), .A2(new_n1177), .ZN(G375));
  NOR2_X1   g0978(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1091), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n937), .B(KEYINPUT123), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT124), .Z(new_n1185));
  NAND2_X1  g0985(.A1(new_n1053), .A2(new_n761), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n753), .B1(new_n790), .B2(G68), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1153), .A2(new_n273), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n1112), .A2(new_n719), .B1(new_n957), .B2(new_n706), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n710), .A2(new_n283), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n727), .A2(new_n1105), .B1(new_n713), .B2(new_n808), .ZN(new_n1191));
  NOR4_X1   g0991(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1192), .B1(new_n202), .B2(new_n732), .C1(new_n1104), .C2(new_n724), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n706), .A2(new_n716), .B1(new_n713), .B2(new_n238), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n273), .B(new_n1194), .C1(G77), .C2(new_n792), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n725), .A2(G303), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n727), .A2(new_n486), .B1(new_n710), .B2(new_n240), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G116), .B2(new_n739), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1195), .A2(new_n988), .A3(new_n1196), .A4(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1193), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1187), .B1(new_n1200), .B2(new_n703), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1077), .A2(new_n752), .B1(new_n1186), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1185), .A2(new_n1202), .ZN(G381));
  OR4_X1    g1003(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n694), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1205));
  AOI21_X1  g1005(.A(KEYINPUT117), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1123), .B1(new_n1207), .B2(new_n1093), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1152), .A2(new_n1208), .A3(new_n1177), .ZN(new_n1209));
  OR4_X1    g1009(.A1(G387), .A2(G381), .A3(new_n1204), .A4(new_n1209), .ZN(G407));
  OAI211_X1 g1010(.A(G407), .B(G213), .C1(G343), .C2(new_n1209), .ZN(G409));
  XNOR2_X1  g1011(.A(G387), .B(G390), .ZN(new_n1212));
  XOR2_X1   g1012(.A(G393), .B(G396), .Z(new_n1213));
  XNOR2_X1  g1013(.A(new_n1212), .B(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT61), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n694), .B1(new_n1179), .B2(KEYINPUT60), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n1181), .B2(KEYINPUT60), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1218), .A2(G384), .A3(new_n1202), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1202), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n815), .B1(new_n1217), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(G2897), .ZN(new_n1223));
  NOR3_X1   g1023(.A1(new_n643), .A2(new_n1223), .A3(G343), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1222), .B(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1208), .B1(new_n1152), .B2(new_n1177), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1147), .A2(new_n1150), .A3(new_n1183), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n1177), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(G378), .A2(new_n1228), .B1(new_n643), .B2(G343), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1226), .A2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1215), .B1(new_n1225), .B2(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1214), .A2(new_n1231), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1226), .A2(new_n1229), .A3(new_n1222), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(KEYINPUT63), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1222), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT125), .B1(new_n1230), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT125), .ZN(new_n1237));
  NOR4_X1   g1037(.A1(new_n1226), .A2(new_n1229), .A3(new_n1222), .A4(new_n1237), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1236), .A2(new_n1238), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1232), .B(new_n1234), .C1(KEYINPUT63), .C2(new_n1239), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1233), .A2(KEYINPUT62), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT62), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1242), .B1(new_n1236), .B2(new_n1238), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1241), .B1(new_n1243), .B2(KEYINPUT126), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT126), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1245), .B(new_n1242), .C1(new_n1236), .C2(new_n1238), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1231), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1214), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1240), .B1(new_n1247), .B2(new_n1248), .ZN(G405));
  INV_X1    g1049(.A(new_n1226), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n1209), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(new_n1222), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1252), .B(new_n1214), .ZN(G402));
endmodule


