//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 1 0 0 0 0 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 1 0 1 1 0 1 0 1 1 1 1 0 1 1 0 1 1 0 0 0 1 0 1 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1250, new_n1251, new_n1252, new_n1253, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT0), .Z(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n209), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n214), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT64), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n225), .A2(new_n226), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n211), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(KEYINPUT1), .ZN(new_n233));
  OR2_X1    g0033(.A1(new_n232), .A2(KEYINPUT1), .ZN(new_n234));
  NAND3_X1  g0034(.A1(new_n219), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(KEYINPUT65), .Z(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  INV_X1    g0037(.A(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT66), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n247), .B(new_n248), .Z(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G1), .A3(G13), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  AND2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(G1698), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G222), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n267), .A2(G223), .A3(G1698), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n268), .B1(new_n223), .B2(new_n267), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n256), .B1(new_n262), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n255), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G41), .ZN(new_n274));
  INV_X1    g0074(.A(G45), .ZN(new_n275));
  AOI21_X1  g0075(.A(G1), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G274), .ZN(new_n277));
  AND2_X1   g0077(.A1(G1), .A2(G13), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n277), .B1(new_n278), .B2(new_n254), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n273), .A2(G226), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n270), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G169), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n203), .A2(G20), .ZN(new_n284));
  INV_X1    g0084(.A(G150), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G20), .A2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT8), .B(G58), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n209), .A2(G33), .ZN(new_n289));
  OAI221_X1 g0089(.A(new_n284), .B1(new_n285), .B2(new_n287), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT67), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT67), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n293), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n292), .A2(new_n215), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n290), .A2(new_n295), .B1(new_n202), .B2(new_n297), .ZN(new_n298));
  AND3_X1   g0098(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n278), .B1(new_n299), .B2(new_n293), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n300), .A2(KEYINPUT68), .A3(new_n296), .A4(new_n292), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n292), .A2(new_n294), .A3(new_n215), .A4(new_n296), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT68), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OR3_X1    g0104(.A1(new_n209), .A2(KEYINPUT69), .A3(G1), .ZN(new_n305));
  OAI21_X1  g0105(.A(KEYINPUT69), .B1(new_n209), .B2(G1), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n301), .A2(new_n304), .A3(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n298), .B1(new_n202), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G179), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n270), .A2(new_n310), .A3(new_n280), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n283), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G190), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n281), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(G200), .B2(new_n281), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n309), .B(KEYINPUT9), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT10), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT10), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n315), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n312), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n238), .A2(G1698), .ZN(new_n322));
  OAI221_X1 g0122(.A(new_n322), .B1(G226), .B2(G1698), .C1(new_n257), .C2(new_n258), .ZN(new_n323));
  NAND2_X1  g0123(.A1(G33), .A2(G97), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n255), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n276), .A2(new_n255), .A3(G274), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(new_n222), .B2(new_n272), .ZN(new_n327));
  OR3_X1    g0127(.A1(new_n325), .A2(new_n327), .A3(KEYINPUT13), .ZN(new_n328));
  OAI21_X1  g0128(.A(KEYINPUT13), .B1(new_n325), .B2(new_n327), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(KEYINPUT71), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT71), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n331), .B(KEYINPUT13), .C1(new_n325), .C2(new_n327), .ZN(new_n332));
  AND3_X1   g0132(.A1(new_n330), .A2(G200), .A3(new_n332), .ZN(new_n333));
  AND3_X1   g0133(.A1(new_n328), .A2(G190), .A3(new_n329), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n286), .A2(G50), .ZN(new_n335));
  XNOR2_X1  g0135(.A(new_n335), .B(KEYINPUT72), .ZN(new_n336));
  OAI22_X1  g0136(.A1(new_n289), .A2(new_n223), .B1(new_n209), .B2(G68), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n295), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT11), .ZN(new_n339));
  OR2_X1    g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n296), .A2(G68), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n341), .B(KEYINPUT12), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n342), .B1(new_n338), .B2(new_n339), .ZN(new_n343));
  INV_X1    g0143(.A(new_n302), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n344), .A2(G68), .A3(new_n307), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n340), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  NOR3_X1   g0146(.A1(new_n333), .A2(new_n334), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n330), .A2(G169), .A3(new_n332), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT14), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT14), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n330), .A2(new_n350), .A3(G169), .A4(new_n332), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n328), .A2(G179), .A3(new_n329), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n349), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n347), .B1(new_n346), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n344), .A2(G77), .A3(new_n307), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n288), .A2(new_n287), .B1(new_n209), .B2(new_n223), .ZN(new_n356));
  XNOR2_X1  g0156(.A(KEYINPUT15), .B(G87), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(new_n289), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n295), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n297), .A2(new_n223), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n355), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n326), .B1(new_n224), .B2(new_n272), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n260), .A2(G232), .ZN(new_n363));
  XNOR2_X1  g0163(.A(new_n363), .B(KEYINPUT70), .ZN(new_n364));
  INV_X1    g0164(.A(G1698), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n259), .A2(new_n365), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n366), .A2(G238), .B1(G107), .B2(new_n259), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n362), .B1(new_n368), .B2(new_n256), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n361), .B1(new_n369), .B2(G190), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n255), .B1(new_n364), .B2(new_n367), .ZN(new_n371));
  OAI21_X1  g0171(.A(G200), .B1(new_n371), .B2(new_n362), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n369), .A2(new_n310), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n282), .B1(new_n371), .B2(new_n362), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n374), .A2(new_n361), .A3(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n321), .A2(new_n354), .A3(new_n373), .A4(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n288), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n308), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT75), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n378), .A2(new_n297), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n379), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n302), .A2(new_n303), .B1(new_n305), .B2(new_n306), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n288), .B1(new_n384), .B2(new_n301), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT75), .B1(new_n385), .B2(new_n381), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n295), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT74), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n265), .A2(new_n209), .A3(new_n266), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT7), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT73), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n265), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n266), .ZN(new_n394));
  AND3_X1   g0194(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n393), .A2(KEYINPUT7), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n390), .A2(new_n391), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(G68), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n389), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT7), .B1(new_n259), .B2(new_n209), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n221), .B1(new_n400), .B2(new_n396), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(KEYINPUT74), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(G58), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n405), .A2(new_n221), .ZN(new_n406));
  OAI21_X1  g0206(.A(G20), .B1(new_n406), .B2(new_n201), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n286), .A2(G159), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT16), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n388), .B1(new_n404), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n221), .B1(new_n392), .B2(new_n394), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n410), .B1(new_n413), .B2(new_n409), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n387), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT76), .ZN(new_n416));
  OR2_X1    g0216(.A1(G223), .A2(G1698), .ZN(new_n417));
  INV_X1    g0217(.A(G226), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(G1698), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n417), .B(new_n419), .C1(new_n257), .C2(new_n258), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G33), .A2(G87), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n256), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n255), .A2(G232), .A3(new_n271), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n326), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n416), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n255), .B1(new_n420), .B2(new_n421), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n428), .A2(new_n425), .A3(KEYINPUT76), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n282), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n428), .A2(new_n425), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n310), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT18), .B1(new_n415), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(G200), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(new_n427), .B2(new_n429), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n431), .A2(new_n313), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n415), .A2(KEYINPUT17), .A3(new_n438), .ZN(new_n439));
  AND4_X1   g0239(.A1(KEYINPUT74), .A2(new_n402), .A3(G68), .A4(new_n397), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT74), .B1(new_n401), .B2(new_n402), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n411), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n442), .A2(new_n295), .A3(new_n414), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n380), .B1(new_n379), .B2(new_n382), .ZN(new_n444));
  AOI211_X1 g0244(.A(KEYINPUT75), .B(new_n381), .C1(new_n308), .C2(new_n378), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT18), .ZN(new_n448));
  INV_X1    g0248(.A(new_n433), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n443), .A2(new_n446), .A3(new_n438), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT17), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n434), .A2(new_n439), .A3(new_n450), .A4(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n377), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n267), .A2(G244), .A3(G1698), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G116), .ZN(new_n457));
  OAI211_X1 g0257(.A(G238), .B(new_n365), .C1(new_n257), .C2(new_n258), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n256), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n275), .A2(G1), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n279), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n208), .A2(G45), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n255), .A2(G250), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n460), .A2(G190), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT79), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n460), .A2(new_n466), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G200), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n465), .B1(new_n459), .B2(new_n256), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT79), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n471), .A2(new_n472), .A3(G190), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n267), .A2(new_n209), .A3(G68), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT19), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n209), .B1(new_n324), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n476), .B1(G87), .B2(new_n206), .ZN(new_n477));
  INV_X1    g0277(.A(G97), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n475), .B1(new_n289), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n474), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n295), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n357), .A2(new_n297), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n208), .A2(G33), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n344), .A2(G87), .A3(new_n483), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n468), .A2(new_n470), .A3(new_n473), .A4(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n344), .A2(new_n483), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n481), .B(new_n482), .C1(new_n487), .C2(new_n357), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n471), .A2(new_n310), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n488), .B(new_n489), .C1(G169), .C2(new_n471), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n486), .A2(KEYINPUT80), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n394), .ZN(new_n493));
  OAI21_X1  g0293(.A(G107), .B1(new_n400), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT6), .ZN(new_n495));
  AND2_X1   g0295(.A1(G97), .A2(G107), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n495), .B1(new_n496), .B2(new_n205), .ZN(new_n497));
  INV_X1    g0297(.A(G107), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(KEYINPUT6), .A3(G97), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n500), .A2(G20), .B1(G77), .B2(new_n286), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n388), .B1(new_n494), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n344), .A2(G97), .A3(new_n483), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n296), .A2(G97), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n502), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(G250), .A2(G1698), .ZN(new_n507));
  NAND2_X1  g0307(.A1(KEYINPUT4), .A2(G244), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(G1698), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n267), .A2(new_n509), .B1(G33), .B2(G283), .ZN(new_n510));
  OAI211_X1 g0310(.A(G244), .B(new_n365), .C1(new_n257), .C2(new_n258), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT4), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n256), .ZN(new_n515));
  NAND2_X1  g0315(.A1(KEYINPUT5), .A2(G41), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(KEYINPUT5), .A2(G41), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n461), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n519), .A2(G257), .A3(new_n255), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT5), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n274), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n463), .B1(new_n522), .B2(new_n516), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n279), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n515), .A2(new_n526), .A3(new_n310), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n255), .B1(new_n510), .B2(new_n513), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n282), .B1(new_n528), .B2(new_n525), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(KEYINPUT78), .B1(new_n506), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n515), .A2(new_n526), .A3(KEYINPUT77), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT77), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n528), .B2(new_n525), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n534), .A3(G200), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n528), .A2(new_n525), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G190), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n506), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n500), .A2(G20), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n286), .A2(G77), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n498), .B1(new_n392), .B2(new_n394), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n295), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n505), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n543), .A2(new_n503), .A3(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT78), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n545), .A2(new_n546), .A3(new_n527), .A4(new_n529), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n531), .A2(new_n538), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(KEYINPUT80), .B1(new_n486), .B2(new_n490), .ZN(new_n549));
  NOR3_X1   g0349(.A1(new_n492), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n487), .A2(new_n498), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n297), .A2(new_n498), .ZN(new_n552));
  XNOR2_X1  g0352(.A(new_n552), .B(KEYINPUT25), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT22), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n556), .A2(KEYINPUT81), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n209), .B(G87), .C1(new_n257), .C2(new_n258), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(KEYINPUT81), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n559), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n267), .A2(new_n209), .A3(G87), .A4(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT23), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n209), .B2(G107), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n498), .A2(KEYINPUT23), .A3(G20), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(G116), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n567), .B1(new_n568), .B2(new_n289), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n563), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT82), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n569), .B1(new_n560), .B2(new_n562), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(KEYINPUT82), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n573), .A2(KEYINPUT24), .A3(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n574), .A2(KEYINPUT82), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT24), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n388), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n555), .B1(new_n576), .B2(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(G257), .B(G1698), .C1(new_n257), .C2(new_n258), .ZN(new_n581));
  OAI211_X1 g0381(.A(G250), .B(new_n365), .C1(new_n257), .C2(new_n258), .ZN(new_n582));
  INV_X1    g0382(.A(G294), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n581), .B(new_n582), .C1(new_n264), .C2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n256), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT83), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n584), .A2(KEYINPUT83), .A3(new_n256), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n523), .A2(new_n256), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n589), .A2(G264), .B1(new_n279), .B2(new_n523), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n587), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(G264), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n585), .A2(new_n524), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n591), .A2(G169), .B1(new_n594), .B2(G179), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n580), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n571), .A2(new_n572), .A3(new_n578), .ZN(new_n597));
  OAI21_X1  g0397(.A(KEYINPUT24), .B1(new_n574), .B2(KEYINPUT82), .ZN(new_n598));
  AOI211_X1 g0398(.A(new_n572), .B(new_n569), .C1(new_n562), .C2(new_n560), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n597), .B(new_n295), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n587), .A2(new_n313), .A3(new_n588), .A4(new_n590), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n593), .A2(new_n435), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n600), .A2(new_n554), .A3(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n344), .A2(G116), .A3(new_n483), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n297), .A2(new_n568), .ZN(new_n607));
  AOI21_X1  g0407(.A(G20), .B1(G33), .B2(G283), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n264), .A2(G97), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n608), .A2(new_n609), .B1(G20), .B2(new_n568), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n295), .A2(KEYINPUT20), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(KEYINPUT20), .B1(new_n295), .B2(new_n610), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n606), .B(new_n607), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n589), .A2(G270), .B1(new_n279), .B2(new_n523), .ZN(new_n615));
  OAI211_X1 g0415(.A(G264), .B(G1698), .C1(new_n257), .C2(new_n258), .ZN(new_n616));
  OAI211_X1 g0416(.A(G257), .B(new_n365), .C1(new_n257), .C2(new_n258), .ZN(new_n617));
  INV_X1    g0417(.A(G303), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n616), .B(new_n617), .C1(new_n618), .C2(new_n267), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n256), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(G200), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n614), .B(new_n622), .C1(new_n313), .C2(new_n621), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n613), .A2(G169), .A3(new_n621), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT21), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n615), .A2(G179), .A3(new_n620), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n613), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n613), .A2(new_n621), .A3(KEYINPUT21), .A4(G169), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n623), .A2(new_n626), .A3(new_n628), .A4(new_n629), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n596), .A2(new_n605), .A3(new_n630), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n455), .A2(new_n550), .A3(new_n631), .ZN(G372));
  INV_X1    g0432(.A(new_n490), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n470), .A2(new_n485), .A3(new_n467), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n604), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(new_n548), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n628), .A2(new_n629), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n637), .B(new_n626), .C1(new_n580), .C2(new_n595), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n633), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n486), .A2(new_n490), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT80), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n531), .A2(new_n547), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n642), .A2(KEYINPUT26), .A3(new_n491), .A4(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n490), .A2(new_n634), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n545), .A2(new_n527), .A3(new_n529), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n639), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n455), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n353), .A2(new_n346), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n347), .B2(new_n376), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n439), .A2(new_n453), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n448), .B1(new_n447), .B2(new_n449), .ZN(new_n656));
  AOI211_X1 g0456(.A(KEYINPUT18), .B(new_n433), .C1(new_n443), .C2(new_n446), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n318), .A2(new_n320), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n312), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n651), .A2(new_n661), .ZN(G369));
  NAND2_X1  g0462(.A1(new_n637), .A2(new_n626), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n664), .B(KEYINPUT84), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT27), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT85), .ZN(new_n668));
  INV_X1    g0468(.A(G213), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n669), .B1(new_n665), .B2(new_n666), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n668), .A2(G343), .A3(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(new_n614), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n663), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n630), .B2(new_n672), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  INV_X1    g0475(.A(new_n596), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n604), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n580), .A2(new_n671), .ZN(new_n678));
  OAI22_X1  g0478(.A1(new_n677), .A2(new_n678), .B1(new_n676), .B2(new_n671), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n671), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n681), .B1(new_n637), .B2(new_n626), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n676), .A2(new_n604), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n596), .A2(new_n671), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n680), .A2(new_n686), .ZN(G399));
  INV_X1    g0487(.A(new_n212), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G41), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(G1), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n217), .B2(new_n690), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT28), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n531), .A2(new_n538), .A3(new_n547), .ZN(new_n695));
  INV_X1    g0495(.A(new_n634), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n696), .B1(new_n580), .B2(new_n603), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n638), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n490), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n642), .A2(new_n645), .A3(new_n491), .A4(new_n643), .ZN(new_n700));
  OAI21_X1  g0500(.A(KEYINPUT26), .B1(new_n646), .B2(new_n647), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n671), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(KEYINPUT29), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n681), .B1(new_n639), .B2(new_n649), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT29), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n550), .A2(new_n631), .A3(new_n671), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT30), .ZN(new_n710));
  AOI22_X1  g0510(.A1(new_n584), .A2(new_n256), .B1(new_n589), .B2(G264), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n536), .A2(new_n471), .A3(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n615), .A2(G179), .A3(new_n620), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n710), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n471), .A2(new_n711), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n715), .A2(new_n627), .A3(new_n536), .A4(KEYINPUT30), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n471), .A2(G179), .ZN(new_n717));
  INV_X1    g0517(.A(new_n536), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n717), .A2(new_n718), .A3(new_n621), .A4(new_n593), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n714), .A2(new_n716), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n681), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT31), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n720), .A2(KEYINPUT31), .A3(new_n681), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n709), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n725), .A2(G330), .ZN(new_n726));
  OR3_X1    g0526(.A1(new_n708), .A2(new_n726), .A3(KEYINPUT86), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT86), .B1(new_n708), .B2(new_n726), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n694), .B1(new_n729), .B2(G1), .ZN(G364));
  INV_X1    g0530(.A(G13), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G20), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n208), .B1(new_n732), .B2(G45), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n689), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n212), .A2(new_n267), .ZN(new_n736));
  INV_X1    g0536(.A(G355), .ZN(new_n737));
  OAI22_X1  g0537(.A1(new_n736), .A2(new_n737), .B1(G116), .B2(new_n212), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n249), .A2(new_n275), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n212), .A2(new_n259), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n740), .B1(new_n275), .B2(new_n218), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n738), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G13), .A2(G33), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n215), .B1(G20), .B2(new_n282), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT87), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n735), .B1(new_n742), .B2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT89), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n209), .A2(G190), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n310), .A2(new_n435), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n750), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n751), .A2(KEYINPUT89), .A3(new_n310), .A4(new_n435), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  XOR2_X1   g0557(.A(KEYINPUT90), .B(G159), .Z(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(G20), .B1(new_n753), .B2(new_n313), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT91), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI22_X1  g0565(.A1(KEYINPUT32), .A2(new_n759), .B1(new_n765), .B2(G97), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n209), .A2(new_n310), .A3(new_n435), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT88), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(G190), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n766), .B1(KEYINPUT32), .B2(new_n759), .C1(new_n221), .C2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n768), .A2(new_n313), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n202), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n310), .A2(G200), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(new_n751), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n775), .A2(G20), .A3(G190), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n267), .B1(new_n776), .B2(new_n223), .C1(new_n405), .C2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n209), .A2(G179), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n779), .A2(new_n313), .A3(G200), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n779), .A2(G190), .A3(G200), .ZN(new_n781));
  INV_X1    g0581(.A(G87), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n780), .A2(new_n498), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR4_X1   g0583(.A1(new_n771), .A2(new_n774), .A3(new_n778), .A4(new_n783), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT92), .ZN(new_n785));
  XOR2_X1   g0585(.A(KEYINPUT33), .B(G317), .Z(new_n786));
  INV_X1    g0586(.A(G322), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n770), .A2(new_n786), .B1(new_n787), .B2(new_n777), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n788), .B(KEYINPUT94), .Z(new_n789));
  AOI22_X1  g0589(.A1(G294), .A2(new_n765), .B1(new_n772), .B2(G326), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n791), .A2(KEYINPUT93), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(KEYINPUT93), .ZN(new_n793));
  INV_X1    g0593(.A(new_n776), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n267), .B1(new_n794), .B2(G311), .ZN(new_n795));
  INV_X1    g0595(.A(G283), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n795), .B1(new_n796), .B2(new_n780), .C1(new_n618), .C2(new_n781), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(G329), .B2(new_n757), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n792), .A2(new_n793), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n785), .B1(new_n789), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n749), .B1(new_n800), .B2(new_n746), .ZN(new_n801));
  INV_X1    g0601(.A(new_n745), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n674), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n675), .A2(new_n735), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(G330), .B2(new_n674), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(G396));
  NAND4_X1  g0607(.A1(new_n374), .A2(new_n361), .A3(new_n375), .A4(new_n671), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n361), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n671), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n373), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n809), .B1(new_n813), .B2(new_n376), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n705), .A2(new_n814), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n644), .A2(new_n648), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n671), .B(new_n814), .C1(new_n816), .C2(new_n699), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n726), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(new_n735), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n726), .A2(new_n815), .A3(new_n817), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n746), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n744), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n735), .B1(G77), .B2(new_n823), .ZN(new_n824));
  AOI22_X1  g0624(.A1(G97), .A2(new_n765), .B1(new_n769), .B2(G283), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n757), .A2(G311), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n259), .B1(new_n777), .B2(new_n583), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n780), .A2(new_n782), .B1(new_n781), .B2(new_n498), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n827), .B(new_n828), .C1(G116), .C2(new_n794), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n772), .A2(G303), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n825), .A2(new_n826), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n777), .ZN(new_n832));
  XOR2_X1   g0632(.A(KEYINPUT95), .B(G143), .Z(new_n833));
  AOI22_X1  g0633(.A1(new_n832), .A2(new_n833), .B1(new_n794), .B2(new_n758), .ZN(new_n834));
  INV_X1    g0634(.A(G137), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n834), .B1(new_n770), .B2(new_n285), .C1(new_n835), .C2(new_n773), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT34), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n780), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(G68), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n202), .B2(new_n781), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT96), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n259), .B1(new_n757), .B2(G132), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n405), .B2(new_n764), .ZN(new_n844));
  OR3_X1    g0644(.A1(new_n838), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n836), .A2(new_n837), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n831), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n824), .B1(new_n847), .B2(new_n746), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n814), .B2(new_n744), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n821), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(G384));
  NOR2_X1   g0651(.A1(new_n732), .A2(new_n208), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT37), .ZN(new_n853));
  INV_X1    g0653(.A(new_n409), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n440), .B2(new_n441), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n410), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n387), .B1(new_n856), .B2(new_n412), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n857), .A2(new_n433), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n668), .A2(new_n670), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n442), .A2(new_n295), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT16), .B1(new_n404), .B2(new_n854), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n446), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n861), .A2(new_n864), .B1(new_n415), .B2(new_n438), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n853), .B1(new_n859), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT97), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n857), .A2(new_n860), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n866), .A2(new_n867), .B1(new_n454), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n451), .B1(new_n857), .B2(new_n860), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT37), .B1(new_n870), .B2(new_n858), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n447), .A2(new_n449), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n447), .A2(new_n861), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n872), .A2(new_n873), .A3(new_n853), .A4(new_n451), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n871), .A2(KEYINPUT97), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT38), .B1(new_n869), .B2(new_n875), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n867), .B(KEYINPUT37), .C1(new_n870), .C2(new_n858), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n454), .A2(new_n868), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n875), .A2(KEYINPUT38), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT98), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(new_n721), .B2(new_n722), .ZN(new_n883));
  AOI211_X1 g0683(.A(KEYINPUT98), .B(KEYINPUT31), .C1(new_n720), .C2(new_n681), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n709), .A2(new_n885), .A3(new_n724), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n811), .B1(new_n370), .B2(new_n372), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n374), .A2(new_n361), .A3(new_n375), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n808), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n347), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n681), .A2(new_n346), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n652), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n346), .B(new_n681), .C1(new_n353), .C2(new_n347), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n889), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT40), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n886), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n886), .A2(new_n894), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT38), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n451), .B1(new_n415), .B2(new_n433), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n415), .A2(new_n860), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT37), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n901), .A2(new_n874), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n873), .B1(new_n654), .B2(new_n658), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n898), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n897), .B1(new_n879), .B2(new_n904), .ZN(new_n905));
  OAI22_X1  g0705(.A1(new_n881), .A2(new_n896), .B1(new_n905), .B2(new_n895), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n906), .A2(new_n455), .A3(new_n886), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(G330), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n906), .B1(new_n455), .B2(new_n886), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT39), .B1(new_n904), .B2(new_n879), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n875), .A2(new_n877), .A3(new_n878), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n898), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(KEYINPUT39), .A3(new_n879), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n652), .A2(new_n681), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n912), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n658), .A2(new_n861), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n914), .A2(new_n879), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n892), .A2(new_n893), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n817), .B2(new_n808), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n918), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n917), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n708), .A2(new_n455), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n925), .A2(new_n661), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n924), .B(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n852), .B1(new_n910), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n927), .B2(new_n910), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n500), .A2(KEYINPUT35), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n500), .A2(KEYINPUT35), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n930), .A2(G116), .A3(new_n216), .A4(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT36), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n406), .A2(new_n217), .A3(new_n223), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n221), .A2(G50), .ZN(new_n935));
  OAI211_X1 g0735(.A(G1), .B(new_n731), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n929), .A2(new_n933), .A3(new_n936), .ZN(G367));
  INV_X1    g0737(.A(KEYINPUT46), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n781), .B2(new_n568), .ZN(new_n939));
  INV_X1    g0739(.A(new_n781), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n940), .A2(KEYINPUT46), .A3(G116), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n939), .B(new_n941), .C1(new_n770), .C2(new_n583), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n942), .A2(KEYINPUT109), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(KEYINPUT109), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n780), .A2(new_n478), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n267), .B1(new_n794), .B2(G283), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n618), .B2(new_n777), .ZN(new_n947));
  AOI211_X1 g0747(.A(new_n945), .B(new_n947), .C1(G317), .C2(new_n757), .ZN(new_n948));
  AOI22_X1  g0748(.A1(G107), .A2(new_n765), .B1(new_n772), .B2(G311), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n943), .A2(new_n944), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT110), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n756), .A2(new_n835), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n832), .A2(G150), .B1(new_n794), .B2(G50), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n405), .B2(new_n781), .ZN(new_n954));
  AOI211_X1 g0754(.A(new_n952), .B(new_n954), .C1(new_n769), .C2(new_n758), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT111), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n780), .A2(new_n223), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n956), .B1(new_n957), .B2(new_n259), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n765), .A2(G68), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n772), .A2(new_n833), .ZN(new_n960));
  OAI211_X1 g0760(.A(KEYINPUT111), .B(new_n267), .C1(new_n780), .C2(new_n223), .ZN(new_n961));
  AND4_X1   g0761(.A1(new_n958), .A2(new_n959), .A3(new_n960), .A4(new_n961), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n950), .A2(new_n951), .B1(new_n955), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n951), .B2(new_n950), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT47), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n746), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n671), .A2(new_n485), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n967), .A2(new_n490), .A3(new_n634), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT99), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n969), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n970), .B(new_n971), .C1(new_n490), .C2(new_n967), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n972), .A2(new_n802), .ZN(new_n973));
  INV_X1    g0773(.A(new_n748), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n974), .B1(new_n212), .B2(new_n357), .C1(new_n245), .C2(new_n740), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n975), .A2(KEYINPUT108), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(KEYINPUT108), .ZN(new_n977));
  AND3_X1   g0777(.A1(new_n976), .A2(new_n735), .A3(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n966), .A2(new_n973), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n683), .B1(new_n679), .B2(new_n682), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(new_n675), .Z(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(new_n727), .B2(new_n728), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT107), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n681), .A2(new_n545), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n695), .A2(new_n984), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n647), .A2(new_n671), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI211_X1 g0787(.A(KEYINPUT106), .B(KEYINPUT44), .C1(new_n686), .C2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n987), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT106), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT44), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n990), .A2(new_n991), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n989), .A2(new_n685), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  AND2_X1   g0795(.A1(new_n988), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n686), .A2(KEYINPUT45), .A3(new_n987), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT45), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n989), .B2(new_n685), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n680), .B1(new_n996), .B2(new_n1000), .ZN(new_n1001));
  AND4_X1   g0801(.A1(new_n680), .A2(new_n1000), .A3(new_n988), .A4(new_n995), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n982), .A2(new_n983), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n983), .B1(new_n982), .B2(new_n1003), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n729), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n689), .B(KEYINPUT41), .Z(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n734), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n987), .B(KEYINPUT101), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1011), .A2(new_n680), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT104), .Z(new_n1013));
  INV_X1    g0813(.A(KEYINPUT105), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n987), .A2(new_n676), .A3(new_n604), .A4(new_n682), .ZN(new_n1016));
  OR3_X1    g0816(.A1(new_n1016), .A2(KEYINPUT102), .A3(KEYINPUT42), .ZN(new_n1017));
  OAI21_X1  g0817(.A(KEYINPUT102), .B1(new_n1016), .B2(KEYINPUT42), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n1017), .A2(new_n1018), .B1(KEYINPUT42), .B2(new_n1016), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1011), .A2(new_n676), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n671), .B1(new_n1020), .B2(new_n643), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n972), .A2(KEYINPUT100), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n972), .A2(KEYINPUT100), .ZN(new_n1023));
  NOR3_X1   g0823(.A1(new_n1022), .A2(new_n1023), .A3(KEYINPUT43), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1019), .A2(new_n1021), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT103), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1024), .B1(KEYINPUT43), .B2(new_n972), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n1014), .A2(new_n1013), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1015), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1027), .A2(new_n1030), .A3(new_n1015), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n979), .B1(new_n1010), .B2(new_n1034), .ZN(G387));
  OR3_X1    g0835(.A1(new_n982), .A2(KEYINPUT113), .A3(new_n690), .ZN(new_n1036));
  OAI21_X1  g0836(.A(KEYINPUT113), .B1(new_n982), .B2(new_n690), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n981), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1036), .B(new_n1037), .C1(new_n729), .C2(new_n1038), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n679), .A2(new_n802), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n736), .A2(new_n691), .B1(G107), .B2(new_n212), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n241), .A2(new_n275), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n691), .ZN(new_n1043));
  AOI211_X1 g0843(.A(G45), .B(new_n1043), .C1(G68), .C2(G77), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n288), .A2(G50), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT50), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n740), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1041), .B1(new_n1042), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n735), .B1(new_n1048), .B2(new_n748), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n756), .A2(new_n285), .B1(new_n223), .B2(new_n781), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT112), .Z(new_n1051));
  OAI221_X1 g0851(.A(new_n267), .B1(new_n776), .B2(new_n221), .C1(new_n202), .C2(new_n777), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n945), .B(new_n1052), .C1(new_n772), .C2(G159), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n769), .A2(new_n378), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n357), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n765), .A2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1051), .A2(new_n1053), .A3(new_n1054), .A4(new_n1056), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n764), .A2(new_n796), .B1(new_n583), .B2(new_n781), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n769), .A2(G311), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n832), .A2(G317), .B1(new_n794), .B2(G303), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1059), .B(new_n1060), .C1(new_n773), .C2(new_n787), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT48), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1058), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n1062), .B2(new_n1061), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT49), .Z(new_n1065));
  INV_X1    g0865(.A(G326), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n259), .B1(new_n568), .B2(new_n780), .C1(new_n756), .C2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1057), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1049), .B1(new_n1068), .B2(new_n746), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1038), .A2(new_n734), .B1(new_n1040), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1039), .A2(new_n1070), .ZN(G393));
  NAND2_X1  g0871(.A1(new_n1003), .A2(new_n734), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n974), .B1(new_n478), .B2(new_n212), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n252), .A2(new_n740), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n735), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n1075), .B(KEYINPUT114), .Z(new_n1076));
  AOI22_X1  g0876(.A1(new_n772), .A2(G317), .B1(G311), .B2(new_n832), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT52), .Z(new_n1078));
  AOI21_X1  g0878(.A(new_n267), .B1(new_n794), .B2(G294), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1079), .B1(new_n498), .B2(new_n780), .C1(new_n796), .C2(new_n781), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(G322), .B2(new_n757), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G116), .A2(new_n765), .B1(new_n769), .B2(G303), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1078), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n772), .A2(G150), .B1(G159), .B2(new_n832), .ZN(new_n1084));
  XOR2_X1   g0884(.A(KEYINPUT115), .B(KEYINPUT51), .Z(new_n1085));
  NOR2_X1   g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n259), .B1(new_n794), .B2(new_n378), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1088), .B1(new_n221), .B2(new_n781), .C1(new_n782), .C2(new_n780), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n757), .B2(new_n833), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G77), .A2(new_n765), .B1(new_n769), .B2(G50), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1087), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1083), .B1(new_n1086), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1076), .B1(new_n1093), .B2(new_n746), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1011), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1094), .B1(new_n1095), .B2(new_n802), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1072), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n729), .A2(new_n1038), .ZN(new_n1098));
  OR2_X1    g0898(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1099));
  OAI21_X1  g0899(.A(KEYINPUT107), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n1004), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n690), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1097), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(G390));
  AND3_X1   g0904(.A1(new_n914), .A2(KEYINPUT39), .A3(new_n879), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n743), .B1(new_n1105), .B2(new_n911), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n735), .B1(new_n378), .B2(new_n823), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n259), .B1(new_n781), .B2(new_n782), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n769), .A2(G107), .B1(KEYINPUT117), .B2(new_n1108), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n1109), .B1(KEYINPUT117), .B2(new_n1108), .C1(new_n796), .C2(new_n773), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n777), .A2(new_n568), .B1(new_n776), .B2(new_n478), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(G68), .B2(new_n839), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n1112), .B1(new_n583), .B2(new_n756), .C1(new_n223), .C2(new_n764), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(G128), .A2(new_n772), .B1(new_n769), .B2(G137), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n781), .A2(new_n285), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT53), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n765), .A2(G159), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1114), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(KEYINPUT54), .B(G143), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n267), .B1(new_n776), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(G132), .B2(new_n832), .ZN(new_n1121));
  INV_X1    g0921(.A(G125), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1121), .B1(new_n202), .B2(new_n780), .C1(new_n1122), .C2(new_n756), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n1110), .A2(new_n1113), .B1(new_n1118), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1107), .B1(new_n1124), .B2(new_n746), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1106), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT116), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n916), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n809), .B1(new_n705), .B2(new_n814), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1127), .B(new_n1128), .C1(new_n1129), .C2(new_n921), .ZN(new_n1130));
  OAI21_X1  g0930(.A(KEYINPUT116), .B1(new_n922), .B2(new_n916), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1130), .B(new_n1131), .C1(new_n1105), .C2(new_n911), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n887), .A2(new_n888), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n703), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n920), .B1(new_n1134), .B2(new_n809), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n904), .A2(new_n879), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1135), .A2(new_n1128), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n726), .A2(new_n814), .A3(new_n920), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1132), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1137), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1128), .B1(new_n1129), .B2(new_n921), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n912), .A2(new_n915), .B1(new_n1141), .B2(KEYINPUT116), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1140), .B1(new_n1142), .B2(new_n1130), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n886), .A2(G330), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n894), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1139), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1126), .B1(new_n1146), .B2(new_n733), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1144), .A2(new_n455), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n925), .A2(new_n661), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1129), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1145), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n920), .B1(new_n726), .B2(new_n814), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1150), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1134), .A2(new_n809), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n886), .A2(G330), .A3(new_n814), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n921), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1138), .A2(new_n1154), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1149), .B1(new_n1153), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n690), .B1(new_n1146), .B2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1139), .B(new_n1158), .C1(new_n1143), .C2(new_n1145), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1147), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(G378));
  INV_X1    g0963(.A(new_n1149), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n917), .A2(new_n923), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n861), .A2(new_n309), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n321), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n321), .A2(new_n1167), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  OR3_X1    g0971(.A1(new_n1168), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1171), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n906), .B2(G330), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n897), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n895), .B1(new_n1136), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n896), .B1(new_n914), .B2(new_n879), .ZN(new_n1178));
  OAI211_X1 g0978(.A(G330), .B(new_n1174), .C1(new_n1177), .C2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1166), .B1(new_n1175), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(G330), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1174), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n924), .A2(new_n1184), .A3(new_n1179), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1181), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1165), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT57), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(KEYINPUT122), .A3(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT122), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1161), .A2(new_n1164), .B1(new_n1181), .B2(new_n1185), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1190), .B1(new_n1191), .B2(KEYINPUT57), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n690), .B1(new_n1191), .B2(KEYINPUT57), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1189), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1183), .A2(new_n743), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n735), .B1(G50), .B2(new_n823), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n478), .A2(new_n770), .B1(new_n773), .B2(new_n568), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n757), .A2(G283), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n780), .A2(new_n405), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n832), .A2(G107), .B1(new_n794), .B2(new_n1055), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n959), .A2(new_n1198), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n274), .B(new_n259), .C1(new_n781), .C2(new_n223), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT118), .Z(new_n1204));
  NOR3_X1   g1004(.A1(new_n1197), .A2(new_n1202), .A3(new_n1204), .ZN(new_n1205));
  XOR2_X1   g1005(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n1206));
  XNOR2_X1  g1006(.A(new_n1205), .B(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(G50), .B1(new_n264), .B2(new_n274), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n267), .B2(G41), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n832), .A2(G128), .B1(new_n794), .B2(G137), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n781), .B2(new_n1119), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n773), .A2(new_n1122), .B1(new_n285), .B2(new_n764), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT120), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1211), .B(new_n1213), .C1(G132), .C2(new_n769), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT59), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n757), .A2(G124), .ZN(new_n1218));
  AOI211_X1 g1018(.A(G33), .B(G41), .C1(new_n839), .C2(new_n758), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(new_n1214), .C2(new_n1215), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1207), .B(new_n1209), .C1(new_n1217), .C2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT121), .ZN(new_n1222));
  OR2_X1    g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n822), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1196), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1186), .A2(new_n734), .B1(new_n1195), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1194), .A2(new_n1226), .ZN(G375));
  NAND3_X1  g1027(.A1(new_n1153), .A2(new_n1149), .A3(new_n1157), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1159), .A2(new_n1009), .A3(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1153), .A2(new_n1157), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n921), .A2(new_n743), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n735), .B1(G68), .B2(new_n823), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n267), .B1(new_n776), .B2(new_n285), .C1(new_n835), .C2(new_n777), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1199), .B(new_n1233), .C1(G159), .C2(new_n940), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1119), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(G50), .A2(new_n765), .B1(new_n769), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n757), .A2(G128), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n772), .A2(G132), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1234), .A2(new_n1236), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(G116), .A2(new_n769), .B1(new_n772), .B2(G294), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n259), .B1(new_n776), .B2(new_n498), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n957), .B(new_n1241), .C1(G283), .C2(new_n832), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1240), .A2(new_n1056), .A3(new_n1242), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n756), .A2(new_n618), .B1(new_n478), .B2(new_n781), .ZN(new_n1244));
  XOR2_X1   g1044(.A(new_n1244), .B(KEYINPUT123), .Z(new_n1245));
  OAI21_X1  g1045(.A(new_n1239), .B1(new_n1243), .B2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1232), .B1(new_n1246), .B2(new_n746), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1230), .A2(new_n734), .B1(new_n1231), .B2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1229), .A2(new_n1248), .ZN(G381));
  NAND3_X1  g1049(.A1(new_n1194), .A2(new_n1162), .A3(new_n1226), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1039), .A2(new_n806), .A3(new_n1070), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(G381), .A2(G384), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1251), .A2(new_n1103), .A3(new_n1252), .ZN(new_n1253));
  OR3_X1    g1053(.A1(new_n1250), .A2(G387), .A3(new_n1253), .ZN(G407));
  OAI211_X1 g1054(.A(G407), .B(G213), .C1(G343), .C2(new_n1250), .ZN(G409));
  NAND3_X1  g1055(.A1(new_n1194), .A2(G378), .A3(new_n1226), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1226), .B1(new_n1187), .B2(new_n1008), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n1162), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1256), .A2(new_n1258), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n669), .A2(G343), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT60), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n690), .B(new_n1158), .C1(new_n1263), .C2(new_n1228), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1228), .ZN(new_n1265));
  AOI21_X1  g1065(.A(KEYINPUT124), .B1(new_n1265), .B2(KEYINPUT60), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1265), .A2(KEYINPUT124), .A3(KEYINPUT60), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1264), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1268), .A2(G384), .A3(new_n1248), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(G384), .B1(new_n1268), .B2(new_n1248), .ZN(new_n1271));
  OAI211_X1 g1071(.A(G2897), .B(new_n1260), .C1(new_n1270), .C2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1271), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1260), .A2(G2897), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1273), .A2(new_n1269), .A3(new_n1274), .ZN(new_n1275));
  AND2_X1   g1075(.A1(new_n1272), .A2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT61), .B1(new_n1262), .B2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT63), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1273), .A2(new_n1269), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1278), .B1(new_n1262), .B2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n806), .B1(new_n1039), .B2(new_n1070), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1251), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(G387), .A2(new_n1103), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(new_n1100), .A2(new_n1004), .B1(new_n727), .B2(new_n728), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n733), .B1(new_n1285), .B2(new_n1008), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1033), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1287), .A2(new_n1031), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1289), .A2(new_n979), .A3(G390), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1284), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT125), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1283), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  AOI211_X1 g1093(.A(KEYINPUT125), .B(new_n1282), .C1(new_n1284), .C2(new_n1290), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1260), .B1(new_n1256), .B2(new_n1258), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1279), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1296), .A2(KEYINPUT63), .A3(new_n1297), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1277), .A2(new_n1280), .A3(new_n1295), .A4(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT62), .ZN(new_n1300));
  AND3_X1   g1100(.A1(new_n1296), .A2(new_n1300), .A3(new_n1297), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT61), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1272), .A2(new_n1275), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1302), .B1(new_n1296), .B2(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1300), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1305));
  NOR3_X1   g1105(.A1(new_n1301), .A2(new_n1304), .A3(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(KEYINPUT126), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1307));
  AOI21_X1  g1107(.A(G390), .B1(new_n1289), .B2(new_n979), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n979), .ZN(new_n1309));
  AOI211_X1 g1109(.A(new_n1309), .B(new_n1103), .C1(new_n1286), .C2(new_n1288), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1292), .B1(new_n1308), .B2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n1282), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT126), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1291), .A2(new_n1292), .A3(new_n1283), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1312), .A2(new_n1313), .A3(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1307), .A2(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1299), .B1(new_n1306), .B2(new_n1316), .ZN(G405));
  INV_X1    g1117(.A(KEYINPUT127), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1279), .A2(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1319), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1279), .A2(new_n1318), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(G375), .A2(G378), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1321), .A2(new_n1322), .A3(new_n1250), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1297), .A2(KEYINPUT127), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1312), .A2(new_n1325), .A3(new_n1314), .ZN(new_n1326));
  AND3_X1   g1126(.A1(new_n1320), .A2(new_n1324), .A3(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1324), .B1(new_n1320), .B2(new_n1326), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1327), .A2(new_n1328), .ZN(G402));
endmodule


