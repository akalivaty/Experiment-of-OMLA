

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U561 ( .A(n644), .B(KEYINPUT30), .ZN(n646) );
  AND2_X1 U562 ( .A1(n713), .A2(n712), .ZN(n716) );
  XNOR2_X1 U563 ( .A(n714), .B(KEYINPUT98), .ZN(n715) );
  NOR2_X1 U564 ( .A1(n690), .A2(n726), .ZN(n742) );
  XNOR2_X1 U565 ( .A(KEYINPUT91), .B(n732), .ZN(n527) );
  OR2_X1 U566 ( .A1(n680), .A2(n679), .ZN(n685) );
  INV_X1 U567 ( .A(G168), .ZN(n645) );
  AND2_X1 U568 ( .A1(n646), .A2(n645), .ZN(n650) );
  NOR2_X1 U569 ( .A1(G1966), .A2(n705), .ZN(n721) );
  AND2_X1 U570 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U571 ( .A1(n733), .A2(n527), .ZN(n734) );
  INV_X1 U572 ( .A(G2105), .ZN(n543) );
  OR2_X1 U573 ( .A1(n737), .A2(n736), .ZN(n758) );
  XOR2_X1 U574 ( .A(KEYINPUT1), .B(n528), .Z(n802) );
  NOR2_X1 U575 ( .A1(n670), .A2(n669), .ZN(n672) );
  NAND2_X1 U576 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U577 ( .A(n672), .B(n671), .ZN(n1012) );
  XOR2_X1 U578 ( .A(G543), .B(KEYINPUT0), .Z(n608) );
  NOR2_X1 U579 ( .A1(G651), .A2(n608), .ZN(n801) );
  NAND2_X1 U580 ( .A1(n801), .A2(G47), .ZN(n530) );
  XOR2_X1 U581 ( .A(KEYINPUT70), .B(G651), .Z(n532) );
  NOR2_X1 U582 ( .A1(G543), .A2(n532), .ZN(n528) );
  NAND2_X1 U583 ( .A1(G60), .A2(n802), .ZN(n529) );
  NAND2_X1 U584 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U585 ( .A(n531), .B(KEYINPUT71), .ZN(n534) );
  NOR2_X1 U586 ( .A1(n608), .A2(n532), .ZN(n798) );
  NAND2_X1 U587 ( .A1(G72), .A2(n798), .ZN(n533) );
  NAND2_X1 U588 ( .A1(n534), .A2(n533), .ZN(n537) );
  NOR2_X1 U589 ( .A1(G651), .A2(G543), .ZN(n797) );
  NAND2_X1 U590 ( .A1(G85), .A2(n797), .ZN(n535) );
  XNOR2_X1 U591 ( .A(KEYINPUT69), .B(n535), .ZN(n536) );
  NOR2_X1 U592 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U593 ( .A(KEYINPUT72), .B(n538), .Z(G290) );
  NOR2_X1 U594 ( .A1(G2105), .A2(G2104), .ZN(n539) );
  XOR2_X2 U595 ( .A(KEYINPUT17), .B(n539), .Z(n902) );
  NAND2_X1 U596 ( .A1(G138), .A2(n902), .ZN(n542) );
  NAND2_X1 U597 ( .A1(n543), .A2(G2104), .ZN(n540) );
  XNOR2_X1 U598 ( .A(n540), .B(KEYINPUT67), .ZN(n903) );
  NAND2_X1 U599 ( .A1(G102), .A2(n903), .ZN(n541) );
  NAND2_X1 U600 ( .A1(n542), .A2(n541), .ZN(n548) );
  AND2_X1 U601 ( .A1(G2105), .A2(G2104), .ZN(n897) );
  NAND2_X1 U602 ( .A1(n897), .A2(G114), .ZN(n546) );
  NOR2_X1 U603 ( .A1(n543), .A2(G2104), .ZN(n544) );
  XNOR2_X1 U604 ( .A(n544), .B(KEYINPUT66), .ZN(n898) );
  NAND2_X1 U605 ( .A1(G126), .A2(n898), .ZN(n545) );
  NAND2_X1 U606 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U607 ( .A1(n548), .A2(n547), .ZN(G164) );
  NAND2_X1 U608 ( .A1(G101), .A2(n903), .ZN(n549) );
  XOR2_X1 U609 ( .A(KEYINPUT23), .B(n549), .Z(n557) );
  NAND2_X1 U610 ( .A1(G113), .A2(n897), .ZN(n551) );
  NAND2_X1 U611 ( .A1(G137), .A2(n902), .ZN(n550) );
  NAND2_X1 U612 ( .A1(n551), .A2(n550), .ZN(n553) );
  INV_X1 U613 ( .A(KEYINPUT68), .ZN(n552) );
  XNOR2_X1 U614 ( .A(n553), .B(n552), .ZN(n555) );
  NAND2_X1 U615 ( .A1(G125), .A2(n898), .ZN(n554) );
  AND2_X1 U616 ( .A1(n555), .A2(n554), .ZN(n556) );
  AND2_X1 U617 ( .A1(n557), .A2(n556), .ZN(G160) );
  NAND2_X1 U618 ( .A1(n801), .A2(G51), .ZN(n558) );
  XOR2_X1 U619 ( .A(KEYINPUT79), .B(n558), .Z(n560) );
  NAND2_X1 U620 ( .A1(G63), .A2(n802), .ZN(n559) );
  NAND2_X1 U621 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U622 ( .A(KEYINPUT6), .B(n561), .ZN(n568) );
  NAND2_X1 U623 ( .A1(n797), .A2(G89), .ZN(n562) );
  XNOR2_X1 U624 ( .A(n562), .B(KEYINPUT4), .ZN(n564) );
  NAND2_X1 U625 ( .A1(G76), .A2(n798), .ZN(n563) );
  NAND2_X1 U626 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U627 ( .A(KEYINPUT78), .B(n565), .Z(n566) );
  XNOR2_X1 U628 ( .A(KEYINPUT5), .B(n566), .ZN(n567) );
  NOR2_X1 U629 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U630 ( .A(n569), .B(KEYINPUT7), .Z(n570) );
  XNOR2_X1 U631 ( .A(KEYINPUT80), .B(n570), .ZN(G168) );
  NAND2_X1 U632 ( .A1(G90), .A2(n797), .ZN(n572) );
  NAND2_X1 U633 ( .A1(G77), .A2(n798), .ZN(n571) );
  NAND2_X1 U634 ( .A1(n572), .A2(n571), .ZN(n574) );
  XOR2_X1 U635 ( .A(KEYINPUT73), .B(KEYINPUT9), .Z(n573) );
  XNOR2_X1 U636 ( .A(n574), .B(n573), .ZN(n578) );
  NAND2_X1 U637 ( .A1(n802), .A2(G64), .ZN(n576) );
  NAND2_X1 U638 ( .A1(n801), .A2(G52), .ZN(n575) );
  AND2_X1 U639 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U640 ( .A1(n578), .A2(n577), .ZN(G301) );
  NAND2_X1 U641 ( .A1(G65), .A2(n802), .ZN(n585) );
  NAND2_X1 U642 ( .A1(G91), .A2(n797), .ZN(n580) );
  NAND2_X1 U643 ( .A1(G78), .A2(n798), .ZN(n579) );
  NAND2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U645 ( .A1(n801), .A2(G53), .ZN(n581) );
  XOR2_X1 U646 ( .A(KEYINPUT74), .B(n581), .Z(n582) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U648 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U649 ( .A(KEYINPUT75), .B(n586), .Z(G299) );
  XNOR2_X1 U650 ( .A(KEYINPUT81), .B(KEYINPUT8), .ZN(n587) );
  XNOR2_X1 U651 ( .A(n587), .B(G168), .ZN(G286) );
  NAND2_X1 U652 ( .A1(G88), .A2(n797), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(KEYINPUT86), .ZN(n591) );
  NAND2_X1 U654 ( .A1(G50), .A2(n801), .ZN(n589) );
  XOR2_X1 U655 ( .A(KEYINPUT85), .B(n589), .Z(n590) );
  NAND2_X1 U656 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U657 ( .A1(G62), .A2(n802), .ZN(n593) );
  NAND2_X1 U658 ( .A1(G75), .A2(n798), .ZN(n592) );
  NAND2_X1 U659 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U660 ( .A1(n595), .A2(n594), .ZN(G166) );
  INV_X1 U661 ( .A(G166), .ZN(G303) );
  XOR2_X1 U662 ( .A(KEYINPUT84), .B(KEYINPUT2), .Z(n597) );
  NAND2_X1 U663 ( .A1(G73), .A2(n798), .ZN(n596) );
  XNOR2_X1 U664 ( .A(n597), .B(n596), .ZN(n601) );
  NAND2_X1 U665 ( .A1(G86), .A2(n797), .ZN(n599) );
  NAND2_X1 U666 ( .A1(G48), .A2(n801), .ZN(n598) );
  NAND2_X1 U667 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U668 ( .A1(n601), .A2(n600), .ZN(n603) );
  NAND2_X1 U669 ( .A1(G61), .A2(n802), .ZN(n602) );
  NAND2_X1 U670 ( .A1(n603), .A2(n602), .ZN(G305) );
  NAND2_X1 U671 ( .A1(G49), .A2(n801), .ZN(n605) );
  NAND2_X1 U672 ( .A1(G74), .A2(G651), .ZN(n604) );
  NAND2_X1 U673 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U674 ( .A1(n802), .A2(n606), .ZN(n607) );
  XOR2_X1 U675 ( .A(KEYINPUT83), .B(n607), .Z(n610) );
  NAND2_X1 U676 ( .A1(n608), .A2(G87), .ZN(n609) );
  NAND2_X1 U677 ( .A1(n610), .A2(n609), .ZN(G288) );
  XOR2_X1 U678 ( .A(KEYINPUT38), .B(KEYINPUT88), .Z(n612) );
  NAND2_X1 U679 ( .A1(G105), .A2(n903), .ZN(n611) );
  XNOR2_X1 U680 ( .A(n612), .B(n611), .ZN(n616) );
  NAND2_X1 U681 ( .A1(G117), .A2(n897), .ZN(n614) );
  NAND2_X1 U682 ( .A1(G141), .A2(n902), .ZN(n613) );
  NAND2_X1 U683 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U684 ( .A1(n616), .A2(n615), .ZN(n618) );
  NAND2_X1 U685 ( .A1(G129), .A2(n898), .ZN(n617) );
  NAND2_X1 U686 ( .A1(n618), .A2(n617), .ZN(n882) );
  NOR2_X1 U687 ( .A1(G1996), .A2(n882), .ZN(n982) );
  NAND2_X1 U688 ( .A1(G1996), .A2(n882), .ZN(n619) );
  XNOR2_X1 U689 ( .A(n619), .B(KEYINPUT89), .ZN(n627) );
  NAND2_X1 U690 ( .A1(G131), .A2(n902), .ZN(n621) );
  NAND2_X1 U691 ( .A1(G95), .A2(n903), .ZN(n620) );
  NAND2_X1 U692 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U693 ( .A1(n897), .A2(G107), .ZN(n623) );
  NAND2_X1 U694 ( .A1(G119), .A2(n898), .ZN(n622) );
  NAND2_X1 U695 ( .A1(n623), .A2(n622), .ZN(n624) );
  OR2_X1 U696 ( .A1(n625), .A2(n624), .ZN(n883) );
  AND2_X1 U697 ( .A1(G1991), .A2(n883), .ZN(n626) );
  NOR2_X1 U698 ( .A1(n627), .A2(n626), .ZN(n988) );
  INV_X1 U699 ( .A(n988), .ZN(n631) );
  NOR2_X1 U700 ( .A1(G1991), .A2(n883), .ZN(n977) );
  NOR2_X1 U701 ( .A1(G1986), .A2(G290), .ZN(n628) );
  XNOR2_X1 U702 ( .A(KEYINPUT102), .B(n628), .ZN(n629) );
  NOR2_X1 U703 ( .A1(n977), .A2(n629), .ZN(n630) );
  NOR2_X1 U704 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U705 ( .A1(n982), .A2(n632), .ZN(n633) );
  XNOR2_X1 U706 ( .A(KEYINPUT39), .B(n633), .ZN(n635) );
  NOR2_X1 U707 ( .A1(G164), .A2(G1384), .ZN(n640) );
  NAND2_X1 U708 ( .A1(G160), .A2(G40), .ZN(n634) );
  NOR2_X1 U709 ( .A1(n640), .A2(n634), .ZN(n771) );
  NAND2_X1 U710 ( .A1(n635), .A2(n771), .ZN(n733) );
  INV_X1 U711 ( .A(n733), .ZN(n639) );
  XNOR2_X1 U712 ( .A(KEYINPUT87), .B(G1986), .ZN(n636) );
  XNOR2_X1 U713 ( .A(n636), .B(G290), .ZN(n1018) );
  NAND2_X1 U714 ( .A1(n1018), .A2(n988), .ZN(n637) );
  NAND2_X1 U715 ( .A1(n637), .A2(n771), .ZN(n638) );
  OR2_X1 U716 ( .A1(n639), .A2(n638), .ZN(n754) );
  INV_X1 U717 ( .A(n754), .ZN(n737) );
  AND2_X1 U718 ( .A1(n640), .A2(G40), .ZN(n641) );
  NAND2_X1 U719 ( .A1(G160), .A2(n641), .ZN(n707) );
  INV_X1 U720 ( .A(n707), .ZN(n690) );
  INV_X1 U721 ( .A(G8), .ZN(n726) );
  INV_X1 U722 ( .A(n742), .ZN(n705) );
  NOR2_X1 U723 ( .A1(G2084), .A2(n707), .ZN(n642) );
  XNOR2_X1 U724 ( .A(KEYINPUT92), .B(n642), .ZN(n717) );
  OR2_X1 U725 ( .A1(n726), .A2(n717), .ZN(n643) );
  NOR2_X1 U726 ( .A1(n721), .A2(n643), .ZN(n644) );
  XOR2_X1 U727 ( .A(G2078), .B(KEYINPUT25), .Z(n937) );
  NOR2_X1 U728 ( .A1(n937), .A2(n707), .ZN(n648) );
  NOR2_X1 U729 ( .A1(n690), .A2(G1961), .ZN(n647) );
  NOR2_X1 U730 ( .A1(n648), .A2(n647), .ZN(n653) );
  AND2_X1 U731 ( .A1(G301), .A2(n653), .ZN(n649) );
  NOR2_X1 U732 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U733 ( .A(n651), .B(KEYINPUT31), .Z(n652) );
  XNOR2_X1 U734 ( .A(n652), .B(KEYINPUT96), .ZN(n704) );
  NOR2_X1 U735 ( .A1(n653), .A2(G301), .ZN(n654) );
  XNOR2_X1 U736 ( .A(n654), .B(KEYINPUT93), .ZN(n702) );
  NAND2_X1 U737 ( .A1(G92), .A2(n797), .ZN(n656) );
  NAND2_X1 U738 ( .A1(G79), .A2(n798), .ZN(n655) );
  NAND2_X1 U739 ( .A1(n656), .A2(n655), .ZN(n660) );
  NAND2_X1 U740 ( .A1(n801), .A2(G54), .ZN(n658) );
  NAND2_X1 U741 ( .A1(G66), .A2(n802), .ZN(n657) );
  NAND2_X1 U742 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U743 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U744 ( .A(KEYINPUT15), .B(n661), .Z(n1009) );
  INV_X1 U745 ( .A(n1009), .ZN(n680) );
  NAND2_X1 U746 ( .A1(n802), .A2(G56), .ZN(n662) );
  XOR2_X1 U747 ( .A(KEYINPUT14), .B(n662), .Z(n670) );
  NAND2_X1 U748 ( .A1(n797), .A2(G81), .ZN(n663) );
  XNOR2_X1 U749 ( .A(n663), .B(KEYINPUT12), .ZN(n665) );
  NAND2_X1 U750 ( .A1(G68), .A2(n798), .ZN(n664) );
  NAND2_X1 U751 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U752 ( .A(n666), .B(KEYINPUT13), .ZN(n668) );
  NAND2_X1 U753 ( .A1(G43), .A2(n801), .ZN(n667) );
  NAND2_X1 U754 ( .A1(n668), .A2(n667), .ZN(n669) );
  INV_X1 U755 ( .A(KEYINPUT76), .ZN(n671) );
  INV_X1 U756 ( .A(G1996), .ZN(n934) );
  NOR2_X1 U757 ( .A1(n707), .A2(n934), .ZN(n674) );
  XOR2_X1 U758 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n673) );
  XNOR2_X1 U759 ( .A(n674), .B(n673), .ZN(n676) );
  NAND2_X1 U760 ( .A1(n707), .A2(G1341), .ZN(n675) );
  NAND2_X1 U761 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U762 ( .A1(n1012), .A2(n677), .ZN(n678) );
  XNOR2_X1 U763 ( .A(KEYINPUT65), .B(n678), .ZN(n679) );
  NAND2_X1 U764 ( .A1(n680), .A2(n679), .ZN(n687) );
  INV_X1 U765 ( .A(G1348), .ZN(n1010) );
  NOR2_X1 U766 ( .A1(n690), .A2(n1010), .ZN(n681) );
  XNOR2_X1 U767 ( .A(n681), .B(KEYINPUT95), .ZN(n683) );
  NAND2_X1 U768 ( .A1(n690), .A2(G2067), .ZN(n682) );
  NAND2_X1 U769 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U770 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U771 ( .A1(n687), .A2(n686), .ZN(n694) );
  INV_X1 U772 ( .A(G299), .ZN(n1025) );
  NAND2_X1 U773 ( .A1(G2072), .A2(n690), .ZN(n688) );
  XNOR2_X1 U774 ( .A(n688), .B(KEYINPUT94), .ZN(n689) );
  XNOR2_X1 U775 ( .A(KEYINPUT27), .B(n689), .ZN(n692) );
  INV_X1 U776 ( .A(G1956), .ZN(n950) );
  NOR2_X1 U777 ( .A1(n690), .A2(n950), .ZN(n691) );
  NOR2_X1 U778 ( .A1(n692), .A2(n691), .ZN(n695) );
  NAND2_X1 U779 ( .A1(n1025), .A2(n695), .ZN(n693) );
  NAND2_X1 U780 ( .A1(n694), .A2(n693), .ZN(n699) );
  NOR2_X1 U781 ( .A1(n1025), .A2(n695), .ZN(n697) );
  INV_X1 U782 ( .A(KEYINPUT28), .ZN(n696) );
  XNOR2_X1 U783 ( .A(n697), .B(n696), .ZN(n698) );
  NAND2_X1 U784 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U785 ( .A(KEYINPUT29), .B(n700), .Z(n701) );
  NAND2_X1 U786 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U787 ( .A1(n704), .A2(n703), .ZN(n719) );
  NAND2_X1 U788 ( .A1(n719), .A2(G286), .ZN(n713) );
  NOR2_X1 U789 ( .A1(G1971), .A2(n705), .ZN(n706) );
  XNOR2_X1 U790 ( .A(KEYINPUT97), .B(n706), .ZN(n710) );
  NOR2_X1 U791 ( .A1(G2090), .A2(n707), .ZN(n708) );
  NOR2_X1 U792 ( .A1(G166), .A2(n708), .ZN(n709) );
  NAND2_X1 U793 ( .A1(n710), .A2(n709), .ZN(n711) );
  OR2_X1 U794 ( .A1(n726), .A2(n711), .ZN(n712) );
  XNOR2_X1 U795 ( .A(KEYINPUT32), .B(KEYINPUT99), .ZN(n714) );
  XNOR2_X1 U796 ( .A(n716), .B(n715), .ZN(n723) );
  NAND2_X1 U797 ( .A1(G8), .A2(n717), .ZN(n718) );
  NAND2_X1 U798 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U799 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U800 ( .A1(n723), .A2(n722), .ZN(n738) );
  NOR2_X1 U801 ( .A1(G2090), .A2(G303), .ZN(n724) );
  XNOR2_X1 U802 ( .A(n724), .B(KEYINPUT101), .ZN(n725) );
  NOR2_X1 U803 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U804 ( .A1(n738), .A2(n727), .ZN(n728) );
  NOR2_X1 U805 ( .A1(n742), .A2(n728), .ZN(n735) );
  NOR2_X1 U806 ( .A1(G1981), .A2(G305), .ZN(n729) );
  XOR2_X1 U807 ( .A(n729), .B(KEYINPUT90), .Z(n730) );
  XNOR2_X1 U808 ( .A(KEYINPUT24), .B(n730), .ZN(n731) );
  NOR2_X1 U809 ( .A1(n705), .A2(n731), .ZN(n732) );
  NOR2_X1 U810 ( .A1(n735), .A2(n734), .ZN(n736) );
  INV_X1 U811 ( .A(n738), .ZN(n741) );
  NOR2_X1 U812 ( .A1(G1971), .A2(G303), .ZN(n739) );
  NOR2_X1 U813 ( .A1(G1976), .A2(G288), .ZN(n1034) );
  NOR2_X1 U814 ( .A1(n739), .A2(n1034), .ZN(n740) );
  NAND2_X1 U815 ( .A1(n741), .A2(n740), .ZN(n745) );
  AND2_X1 U816 ( .A1(n742), .A2(KEYINPUT100), .ZN(n743) );
  NAND2_X1 U817 ( .A1(G1976), .A2(G288), .ZN(n1026) );
  AND2_X1 U818 ( .A1(n743), .A2(n1026), .ZN(n744) );
  NOR2_X1 U819 ( .A1(KEYINPUT33), .A2(n746), .ZN(n753) );
  INV_X1 U820 ( .A(KEYINPUT100), .ZN(n747) );
  NAND2_X1 U821 ( .A1(n747), .A2(n1034), .ZN(n750) );
  NAND2_X1 U822 ( .A1(n1034), .A2(KEYINPUT33), .ZN(n748) );
  NAND2_X1 U823 ( .A1(n748), .A2(KEYINPUT100), .ZN(n749) );
  NAND2_X1 U824 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U825 ( .A1(n705), .A2(n751), .ZN(n752) );
  NOR2_X1 U826 ( .A1(n753), .A2(n752), .ZN(n756) );
  XOR2_X1 U827 ( .A(G1981), .B(G305), .Z(n1019) );
  AND2_X1 U828 ( .A1(n1019), .A2(n754), .ZN(n755) );
  NAND2_X1 U829 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U830 ( .A1(n758), .A2(n757), .ZN(n769) );
  XOR2_X1 U831 ( .A(G2067), .B(KEYINPUT37), .Z(n770) );
  NAND2_X1 U832 ( .A1(G140), .A2(n902), .ZN(n760) );
  NAND2_X1 U833 ( .A1(G104), .A2(n903), .ZN(n759) );
  NAND2_X1 U834 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U835 ( .A(KEYINPUT34), .B(n761), .ZN(n766) );
  NAND2_X1 U836 ( .A1(n897), .A2(G116), .ZN(n763) );
  NAND2_X1 U837 ( .A1(G128), .A2(n898), .ZN(n762) );
  NAND2_X1 U838 ( .A1(n763), .A2(n762), .ZN(n764) );
  XOR2_X1 U839 ( .A(KEYINPUT35), .B(n764), .Z(n765) );
  NOR2_X1 U840 ( .A1(n766), .A2(n765), .ZN(n767) );
  XOR2_X1 U841 ( .A(KEYINPUT36), .B(n767), .Z(n911) );
  AND2_X1 U842 ( .A1(n770), .A2(n911), .ZN(n990) );
  NAND2_X1 U843 ( .A1(n990), .A2(n771), .ZN(n768) );
  NAND2_X1 U844 ( .A1(n769), .A2(n768), .ZN(n773) );
  NOR2_X1 U845 ( .A1(n770), .A2(n911), .ZN(n1000) );
  NAND2_X1 U846 ( .A1(n1000), .A2(n771), .ZN(n772) );
  XNOR2_X1 U847 ( .A(n774), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U848 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U849 ( .A(G57), .ZN(G237) );
  INV_X1 U850 ( .A(G132), .ZN(G219) );
  INV_X1 U851 ( .A(G82), .ZN(G220) );
  NAND2_X1 U852 ( .A1(G7), .A2(G661), .ZN(n775) );
  XNOR2_X1 U853 ( .A(n775), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U854 ( .A(G223), .ZN(n839) );
  NAND2_X1 U855 ( .A1(n839), .A2(G567), .ZN(n776) );
  XOR2_X1 U856 ( .A(KEYINPUT11), .B(n776), .Z(G234) );
  INV_X1 U857 ( .A(G860), .ZN(n782) );
  OR2_X1 U858 ( .A1(n782), .A2(n1012), .ZN(G153) );
  NOR2_X1 U859 ( .A1(n1009), .A2(G868), .ZN(n777) );
  XNOR2_X1 U860 ( .A(n777), .B(KEYINPUT77), .ZN(n779) );
  NAND2_X1 U861 ( .A1(G868), .A2(G301), .ZN(n778) );
  NAND2_X1 U862 ( .A1(n779), .A2(n778), .ZN(G284) );
  NAND2_X1 U863 ( .A1(G868), .A2(G286), .ZN(n781) );
  INV_X1 U864 ( .A(G868), .ZN(n815) );
  NAND2_X1 U865 ( .A1(G299), .A2(n815), .ZN(n780) );
  NAND2_X1 U866 ( .A1(n781), .A2(n780), .ZN(G297) );
  NAND2_X1 U867 ( .A1(n782), .A2(G559), .ZN(n783) );
  NAND2_X1 U868 ( .A1(n783), .A2(n1009), .ZN(n784) );
  XNOR2_X1 U869 ( .A(n784), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U870 ( .A1(n1012), .A2(G868), .ZN(n787) );
  NAND2_X1 U871 ( .A1(G868), .A2(n1009), .ZN(n785) );
  NOR2_X1 U872 ( .A1(G559), .A2(n785), .ZN(n786) );
  NOR2_X1 U873 ( .A1(n787), .A2(n786), .ZN(G282) );
  NAND2_X1 U874 ( .A1(G123), .A2(n898), .ZN(n788) );
  XNOR2_X1 U875 ( .A(n788), .B(KEYINPUT18), .ZN(n790) );
  NAND2_X1 U876 ( .A1(G111), .A2(n897), .ZN(n789) );
  NAND2_X1 U877 ( .A1(n790), .A2(n789), .ZN(n794) );
  NAND2_X1 U878 ( .A1(G135), .A2(n902), .ZN(n792) );
  NAND2_X1 U879 ( .A1(G99), .A2(n903), .ZN(n791) );
  NAND2_X1 U880 ( .A1(n792), .A2(n791), .ZN(n793) );
  NOR2_X1 U881 ( .A1(n794), .A2(n793), .ZN(n976) );
  XNOR2_X1 U882 ( .A(n976), .B(G2096), .ZN(n796) );
  INV_X1 U883 ( .A(G2100), .ZN(n795) );
  NAND2_X1 U884 ( .A1(n796), .A2(n795), .ZN(G156) );
  NAND2_X1 U885 ( .A1(G93), .A2(n797), .ZN(n800) );
  NAND2_X1 U886 ( .A1(G80), .A2(n798), .ZN(n799) );
  NAND2_X1 U887 ( .A1(n800), .A2(n799), .ZN(n806) );
  NAND2_X1 U888 ( .A1(n801), .A2(G55), .ZN(n804) );
  NAND2_X1 U889 ( .A1(G67), .A2(n802), .ZN(n803) );
  NAND2_X1 U890 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U891 ( .A1(n806), .A2(n805), .ZN(n807) );
  XOR2_X1 U892 ( .A(KEYINPUT82), .B(n807), .Z(n847) );
  XOR2_X1 U893 ( .A(n847), .B(KEYINPUT19), .Z(n809) );
  XNOR2_X1 U894 ( .A(G166), .B(n1025), .ZN(n808) );
  XNOR2_X1 U895 ( .A(n809), .B(n808), .ZN(n810) );
  XOR2_X1 U896 ( .A(n810), .B(G305), .Z(n811) );
  XNOR2_X1 U897 ( .A(G288), .B(n811), .ZN(n812) );
  XNOR2_X1 U898 ( .A(G290), .B(n812), .ZN(n918) );
  NAND2_X1 U899 ( .A1(G559), .A2(n1009), .ZN(n813) );
  XNOR2_X1 U900 ( .A(n813), .B(n1012), .ZN(n845) );
  XOR2_X1 U901 ( .A(n918), .B(n845), .Z(n814) );
  NOR2_X1 U902 ( .A1(n815), .A2(n814), .ZN(n817) );
  NOR2_X1 U903 ( .A1(n847), .A2(G868), .ZN(n816) );
  NOR2_X1 U904 ( .A1(n817), .A2(n816), .ZN(G295) );
  NAND2_X1 U905 ( .A1(G2084), .A2(G2078), .ZN(n818) );
  XOR2_X1 U906 ( .A(KEYINPUT20), .B(n818), .Z(n819) );
  NAND2_X1 U907 ( .A1(G2090), .A2(n819), .ZN(n820) );
  XNOR2_X1 U908 ( .A(KEYINPUT21), .B(n820), .ZN(n821) );
  NAND2_X1 U909 ( .A1(n821), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U910 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U911 ( .A1(G220), .A2(G219), .ZN(n822) );
  XOR2_X1 U912 ( .A(KEYINPUT22), .B(n822), .Z(n823) );
  NOR2_X1 U913 ( .A1(G218), .A2(n823), .ZN(n824) );
  NAND2_X1 U914 ( .A1(G96), .A2(n824), .ZN(n849) );
  NAND2_X1 U915 ( .A1(n849), .A2(G2106), .ZN(n828) );
  NAND2_X1 U916 ( .A1(G69), .A2(G120), .ZN(n825) );
  NOR2_X1 U917 ( .A1(G237), .A2(n825), .ZN(n826) );
  NAND2_X1 U918 ( .A1(G108), .A2(n826), .ZN(n848) );
  NAND2_X1 U919 ( .A1(n848), .A2(G567), .ZN(n827) );
  NAND2_X1 U920 ( .A1(n828), .A2(n827), .ZN(n873) );
  NAND2_X1 U921 ( .A1(G483), .A2(G661), .ZN(n829) );
  NOR2_X1 U922 ( .A1(n873), .A2(n829), .ZN(n844) );
  NAND2_X1 U923 ( .A1(n844), .A2(G36), .ZN(G176) );
  XNOR2_X1 U924 ( .A(G1348), .B(G2435), .ZN(n830) );
  XNOR2_X1 U925 ( .A(n830), .B(G2438), .ZN(n831) );
  XNOR2_X1 U926 ( .A(n831), .B(G1341), .ZN(n837) );
  XOR2_X1 U927 ( .A(G2451), .B(G2446), .Z(n833) );
  XNOR2_X1 U928 ( .A(G2427), .B(G2443), .ZN(n832) );
  XNOR2_X1 U929 ( .A(n833), .B(n832), .ZN(n835) );
  XOR2_X1 U930 ( .A(G2430), .B(G2454), .Z(n834) );
  XNOR2_X1 U931 ( .A(n835), .B(n834), .ZN(n836) );
  XNOR2_X1 U932 ( .A(n837), .B(n836), .ZN(n838) );
  NAND2_X1 U933 ( .A1(n838), .A2(G14), .ZN(n924) );
  XNOR2_X1 U934 ( .A(KEYINPUT103), .B(n924), .ZN(G401) );
  NAND2_X1 U935 ( .A1(G2106), .A2(n839), .ZN(G217) );
  INV_X1 U936 ( .A(G661), .ZN(n841) );
  NAND2_X1 U937 ( .A1(G2), .A2(G15), .ZN(n840) );
  NOR2_X1 U938 ( .A1(n841), .A2(n840), .ZN(n842) );
  XOR2_X1 U939 ( .A(KEYINPUT104), .B(n842), .Z(G259) );
  NAND2_X1 U940 ( .A1(G3), .A2(G1), .ZN(n843) );
  NAND2_X1 U941 ( .A1(n844), .A2(n843), .ZN(G188) );
  NOR2_X1 U943 ( .A1(n845), .A2(G860), .ZN(n846) );
  XOR2_X1 U944 ( .A(n847), .B(n846), .Z(G145) );
  INV_X1 U945 ( .A(G120), .ZN(G236) );
  INV_X1 U946 ( .A(G96), .ZN(G221) );
  INV_X1 U947 ( .A(G69), .ZN(G235) );
  NOR2_X1 U948 ( .A1(n849), .A2(n848), .ZN(n850) );
  XNOR2_X1 U949 ( .A(n850), .B(KEYINPUT105), .ZN(G261) );
  INV_X1 U950 ( .A(G261), .ZN(G325) );
  XOR2_X1 U951 ( .A(KEYINPUT107), .B(KEYINPUT106), .Z(n852) );
  XNOR2_X1 U952 ( .A(G2678), .B(KEYINPUT43), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U954 ( .A(KEYINPUT42), .B(G2072), .Z(n854) );
  XNOR2_X1 U955 ( .A(G2067), .B(G2090), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U957 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U958 ( .A(G2096), .B(G2100), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(n860) );
  XOR2_X1 U960 ( .A(G2084), .B(G2078), .Z(n859) );
  XNOR2_X1 U961 ( .A(n860), .B(n859), .ZN(G227) );
  XOR2_X1 U962 ( .A(G1986), .B(G1956), .Z(n862) );
  XNOR2_X1 U963 ( .A(G1976), .B(G1961), .ZN(n861) );
  XNOR2_X1 U964 ( .A(n862), .B(n861), .ZN(n872) );
  XOR2_X1 U965 ( .A(KEYINPUT110), .B(G2474), .Z(n864) );
  XNOR2_X1 U966 ( .A(G1991), .B(KEYINPUT108), .ZN(n863) );
  XNOR2_X1 U967 ( .A(n864), .B(n863), .ZN(n868) );
  XOR2_X1 U968 ( .A(G1996), .B(G1966), .Z(n866) );
  XNOR2_X1 U969 ( .A(G1981), .B(G1971), .ZN(n865) );
  XNOR2_X1 U970 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U971 ( .A(n868), .B(n867), .Z(n870) );
  XNOR2_X1 U972 ( .A(KEYINPUT109), .B(KEYINPUT41), .ZN(n869) );
  XNOR2_X1 U973 ( .A(n870), .B(n869), .ZN(n871) );
  XNOR2_X1 U974 ( .A(n872), .B(n871), .ZN(G229) );
  INV_X1 U975 ( .A(n873), .ZN(G319) );
  NAND2_X1 U976 ( .A1(G124), .A2(n898), .ZN(n874) );
  XNOR2_X1 U977 ( .A(n874), .B(KEYINPUT44), .ZN(n876) );
  NAND2_X1 U978 ( .A1(G112), .A2(n897), .ZN(n875) );
  NAND2_X1 U979 ( .A1(n876), .A2(n875), .ZN(n880) );
  NAND2_X1 U980 ( .A1(G136), .A2(n902), .ZN(n878) );
  NAND2_X1 U981 ( .A1(G100), .A2(n903), .ZN(n877) );
  NAND2_X1 U982 ( .A1(n878), .A2(n877), .ZN(n879) );
  NOR2_X1 U983 ( .A1(n880), .A2(n879), .ZN(G162) );
  XOR2_X1 U984 ( .A(G162), .B(n976), .Z(n881) );
  XNOR2_X1 U985 ( .A(n882), .B(n881), .ZN(n887) );
  XOR2_X1 U986 ( .A(KEYINPUT112), .B(KEYINPUT46), .Z(n885) );
  XOR2_X1 U987 ( .A(n883), .B(KEYINPUT48), .Z(n884) );
  XNOR2_X1 U988 ( .A(n885), .B(n884), .ZN(n886) );
  XOR2_X1 U989 ( .A(n887), .B(n886), .Z(n889) );
  XNOR2_X1 U990 ( .A(G164), .B(G160), .ZN(n888) );
  XNOR2_X1 U991 ( .A(n889), .B(n888), .ZN(n913) );
  NAND2_X1 U992 ( .A1(n897), .A2(G118), .ZN(n891) );
  NAND2_X1 U993 ( .A1(G130), .A2(n898), .ZN(n890) );
  NAND2_X1 U994 ( .A1(n891), .A2(n890), .ZN(n896) );
  NAND2_X1 U995 ( .A1(G142), .A2(n902), .ZN(n893) );
  NAND2_X1 U996 ( .A1(G106), .A2(n903), .ZN(n892) );
  NAND2_X1 U997 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U998 ( .A(n894), .B(KEYINPUT45), .Z(n895) );
  NOR2_X1 U999 ( .A1(n896), .A2(n895), .ZN(n909) );
  NAND2_X1 U1000 ( .A1(n897), .A2(G115), .ZN(n900) );
  NAND2_X1 U1001 ( .A1(G127), .A2(n898), .ZN(n899) );
  NAND2_X1 U1002 ( .A1(n900), .A2(n899), .ZN(n901) );
  XNOR2_X1 U1003 ( .A(KEYINPUT47), .B(n901), .ZN(n908) );
  NAND2_X1 U1004 ( .A1(G139), .A2(n902), .ZN(n905) );
  NAND2_X1 U1005 ( .A1(G103), .A2(n903), .ZN(n904) );
  NAND2_X1 U1006 ( .A1(n905), .A2(n904), .ZN(n906) );
  XNOR2_X1 U1007 ( .A(KEYINPUT111), .B(n906), .ZN(n907) );
  NAND2_X1 U1008 ( .A1(n908), .A2(n907), .ZN(n992) );
  XNOR2_X1 U1009 ( .A(n909), .B(n992), .ZN(n910) );
  XNOR2_X1 U1010 ( .A(n911), .B(n910), .ZN(n912) );
  XNOR2_X1 U1011 ( .A(n913), .B(n912), .ZN(n914) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n914), .ZN(G395) );
  INV_X1 U1013 ( .A(G301), .ZN(G171) );
  XOR2_X1 U1014 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n916) );
  XNOR2_X1 U1015 ( .A(G171), .B(n1009), .ZN(n915) );
  XNOR2_X1 U1016 ( .A(n916), .B(n915), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(n918), .B(n917), .ZN(n920) );
  XNOR2_X1 U1018 ( .A(G286), .B(n1012), .ZN(n919) );
  XNOR2_X1 U1019 ( .A(n920), .B(n919), .ZN(n921) );
  NOR2_X1 U1020 ( .A1(G37), .A2(n921), .ZN(G397) );
  NOR2_X1 U1021 ( .A1(G227), .A2(G229), .ZN(n923) );
  XNOR2_X1 U1022 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n922) );
  XNOR2_X1 U1023 ( .A(n923), .B(n922), .ZN(n927) );
  NAND2_X1 U1024 ( .A1(G319), .A2(n924), .ZN(n925) );
  XOR2_X1 U1025 ( .A(KEYINPUT115), .B(n925), .Z(n926) );
  NOR2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n929) );
  NOR2_X1 U1027 ( .A1(G395), .A2(G397), .ZN(n928) );
  NAND2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(G225) );
  INV_X1 U1029 ( .A(G225), .ZN(G308) );
  INV_X1 U1030 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1031 ( .A(G25), .B(G1991), .Z(n930) );
  NAND2_X1 U1032 ( .A1(n930), .A2(G28), .ZN(n933) );
  XNOR2_X1 U1033 ( .A(KEYINPUT122), .B(G2072), .ZN(n931) );
  XNOR2_X1 U1034 ( .A(G33), .B(n931), .ZN(n932) );
  NOR2_X1 U1035 ( .A1(n933), .A2(n932), .ZN(n941) );
  XOR2_X1 U1036 ( .A(G2067), .B(G26), .Z(n936) );
  XNOR2_X1 U1037 ( .A(n934), .B(G32), .ZN(n935) );
  NAND2_X1 U1038 ( .A1(n936), .A2(n935), .ZN(n939) );
  XNOR2_X1 U1039 ( .A(G27), .B(n937), .ZN(n938) );
  NOR2_X1 U1040 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1041 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1042 ( .A(n942), .B(KEYINPUT53), .ZN(n945) );
  XOR2_X1 U1043 ( .A(G2084), .B(G34), .Z(n943) );
  XNOR2_X1 U1044 ( .A(KEYINPUT54), .B(n943), .ZN(n944) );
  NAND2_X1 U1045 ( .A1(n945), .A2(n944), .ZN(n947) );
  XNOR2_X1 U1046 ( .A(G35), .B(G2090), .ZN(n946) );
  NOR2_X1 U1047 ( .A1(n947), .A2(n946), .ZN(n972) );
  NOR2_X1 U1048 ( .A1(G29), .A2(n972), .ZN(n948) );
  XNOR2_X1 U1049 ( .A(KEYINPUT55), .B(KEYINPUT121), .ZN(n1002) );
  NAND2_X1 U1050 ( .A1(n948), .A2(n1002), .ZN(n949) );
  NAND2_X1 U1051 ( .A1(G11), .A2(n949), .ZN(n1008) );
  XNOR2_X1 U1052 ( .A(G20), .B(n950), .ZN(n954) );
  XNOR2_X1 U1053 ( .A(G1981), .B(G6), .ZN(n952) );
  XNOR2_X1 U1054 ( .A(G1341), .B(G19), .ZN(n951) );
  NOR2_X1 U1055 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1056 ( .A1(n954), .A2(n953), .ZN(n957) );
  XOR2_X1 U1057 ( .A(KEYINPUT59), .B(G1348), .Z(n955) );
  XNOR2_X1 U1058 ( .A(G4), .B(n955), .ZN(n956) );
  NOR2_X1 U1059 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1060 ( .A(KEYINPUT60), .B(n958), .ZN(n962) );
  XNOR2_X1 U1061 ( .A(G1966), .B(G21), .ZN(n960) );
  XNOR2_X1 U1062 ( .A(G1961), .B(G5), .ZN(n959) );
  NOR2_X1 U1063 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1064 ( .A1(n962), .A2(n961), .ZN(n969) );
  XNOR2_X1 U1065 ( .A(G1976), .B(G23), .ZN(n964) );
  XNOR2_X1 U1066 ( .A(G1971), .B(G22), .ZN(n963) );
  NOR2_X1 U1067 ( .A1(n964), .A2(n963), .ZN(n966) );
  XOR2_X1 U1068 ( .A(G1986), .B(G24), .Z(n965) );
  NAND2_X1 U1069 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1070 ( .A(KEYINPUT58), .B(n967), .ZN(n968) );
  NOR2_X1 U1071 ( .A1(n969), .A2(n968), .ZN(n970) );
  XOR2_X1 U1072 ( .A(KEYINPUT61), .B(n970), .Z(n971) );
  NOR2_X1 U1073 ( .A1(G16), .A2(n971), .ZN(n975) );
  INV_X1 U1074 ( .A(n972), .ZN(n973) );
  NOR2_X1 U1075 ( .A1(n973), .A2(n1002), .ZN(n974) );
  NOR2_X1 U1076 ( .A1(n975), .A2(n974), .ZN(n1006) );
  XNOR2_X1 U1077 ( .A(G160), .B(G2084), .ZN(n980) );
  NOR2_X1 U1078 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1079 ( .A(KEYINPUT117), .B(n978), .Z(n979) );
  NAND2_X1 U1080 ( .A1(n980), .A2(n979), .ZN(n986) );
  XOR2_X1 U1081 ( .A(G2090), .B(G162), .Z(n981) );
  NOR2_X1 U1082 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1083 ( .A(KEYINPUT118), .B(n983), .Z(n984) );
  XOR2_X1 U1084 ( .A(KEYINPUT51), .B(n984), .Z(n985) );
  NOR2_X1 U1085 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1086 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1087 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1088 ( .A(KEYINPUT119), .B(n991), .Z(n998) );
  XNOR2_X1 U1089 ( .A(G2072), .B(KEYINPUT120), .ZN(n993) );
  XNOR2_X1 U1090 ( .A(n993), .B(n992), .ZN(n995) );
  XOR2_X1 U1091 ( .A(G164), .B(G2078), .Z(n994) );
  NOR2_X1 U1092 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1093 ( .A(KEYINPUT50), .B(n996), .ZN(n997) );
  NAND2_X1 U1094 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1095 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1096 ( .A(KEYINPUT52), .B(n1001), .ZN(n1003) );
  NAND2_X1 U1097 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1098 ( .A1(n1004), .A2(G29), .ZN(n1005) );
  NAND2_X1 U1099 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1100 ( .A1(n1008), .A2(n1007), .ZN(n1039) );
  XOR2_X1 U1101 ( .A(KEYINPUT56), .B(G16), .Z(n1036) );
  XNOR2_X1 U1102 ( .A(n1009), .B(KEYINPUT124), .ZN(n1011) );
  XNOR2_X1 U1103 ( .A(n1011), .B(n1010), .ZN(n1016) );
  XOR2_X1 U1104 ( .A(n1012), .B(G1341), .Z(n1014) );
  XNOR2_X1 U1105 ( .A(G171), .B(G1961), .ZN(n1013) );
  NAND2_X1 U1106 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1107 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1108 ( .A1(n1018), .A2(n1017), .ZN(n1024) );
  XNOR2_X1 U1109 ( .A(G168), .B(G1966), .ZN(n1020) );
  NAND2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1111 ( .A(n1021), .B(KEYINPUT57), .ZN(n1022) );
  XNOR2_X1 U1112 ( .A(n1022), .B(KEYINPUT123), .ZN(n1023) );
  NOR2_X1 U1113 ( .A1(n1024), .A2(n1023), .ZN(n1032) );
  XNOR2_X1 U1114 ( .A(G1956), .B(n1025), .ZN(n1027) );
  NAND2_X1 U1115 ( .A1(n1027), .A2(n1026), .ZN(n1030) );
  XNOR2_X1 U1116 ( .A(G166), .B(G1971), .ZN(n1028) );
  XNOR2_X1 U1117 ( .A(KEYINPUT125), .B(n1028), .ZN(n1029) );
  NOR2_X1 U1118 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1119 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NOR2_X1 U1120 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NOR2_X1 U1121 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XOR2_X1 U1122 ( .A(KEYINPUT126), .B(n1037), .Z(n1038) );
  NAND2_X1 U1123 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  XNOR2_X1 U1124 ( .A(n1040), .B(KEYINPUT62), .ZN(n1041) );
  XNOR2_X1 U1125 ( .A(KEYINPUT127), .B(n1041), .ZN(G311) );
  INV_X1 U1126 ( .A(G311), .ZN(G150) );
endmodule

