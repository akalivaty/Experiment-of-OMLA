//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1 0 0 1 0 0 1 0 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n856,
    new_n857, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206));
  INV_X1    g005(.A(G211gat), .ZN(new_n207));
  INV_X1    g006(.A(G218gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n206), .B1(KEYINPUT22), .B2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G211gat), .B(G218gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n211), .B(new_n206), .C1(KEYINPUT22), .C2(new_n209), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(G226gat), .A2(G233gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT27), .B(G183gat), .ZN(new_n218));
  INV_X1    g017(.A(G190gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT69), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(new_n221), .A3(KEYINPUT28), .ZN(new_n222));
  OR2_X1    g021(.A1(new_n221), .A2(KEYINPUT28), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(KEYINPUT28), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n218), .A2(new_n219), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n227), .B(KEYINPUT26), .ZN(new_n228));
  NAND2_X1  g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT65), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n229), .B(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(G183gat), .A2(G190gat), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n231), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n229), .B(KEYINPUT65), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT66), .ZN(new_n238));
  NAND3_X1  g037(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n240));
  OR2_X1    g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(new_n233), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n239), .A2(new_n240), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n241), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT25), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT23), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n227), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n246), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n236), .A2(new_n238), .A3(new_n245), .A4(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n248), .A2(new_n249), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n231), .A2(new_n253), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n243), .A2(new_n239), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n252), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n226), .A2(new_n234), .B1(new_n251), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n217), .B1(new_n257), .B2(KEYINPUT29), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n251), .A2(new_n256), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT68), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n251), .A2(new_n256), .A3(new_n261), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n260), .A2(new_n262), .B1(new_n234), .B2(new_n226), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n258), .B(KEYINPUT72), .C1(new_n263), .C2(new_n217), .ZN(new_n264));
  INV_X1    g063(.A(new_n217), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n222), .A2(new_n232), .A3(new_n233), .A4(new_n225), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT29), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n265), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT72), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n216), .B1(new_n264), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n265), .A2(KEYINPUT29), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  OAI221_X1 g073(.A(new_n216), .B1(new_n217), .B2(new_n267), .C1(new_n263), .C2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n205), .B1(new_n272), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n258), .A2(KEYINPUT72), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n260), .A2(new_n262), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(new_n266), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(new_n265), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n269), .A2(new_n270), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n278), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n204), .B(new_n275), .C1(new_n283), .C2(new_n216), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n277), .A2(new_n284), .A3(KEYINPUT30), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n272), .A2(new_n276), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT30), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n286), .A2(new_n287), .A3(new_n204), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n290));
  XOR2_X1   g089(.A(G155gat), .B(G162gat), .Z(new_n291));
  OR2_X1    g090(.A1(KEYINPUT73), .A2(G141gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(KEYINPUT73), .A2(G141gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n292), .A2(G148gat), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G141gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n295), .A2(G148gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n291), .B1(new_n294), .B2(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(KEYINPUT74), .B(G162gat), .Z(new_n299));
  INV_X1    g098(.A(G155gat), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT2), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT2), .ZN(new_n303));
  INV_X1    g102(.A(G148gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n304), .A2(G141gat), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n303), .B1(new_n296), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(new_n291), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G113gat), .B(G120gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n309), .A2(KEYINPUT1), .ZN(new_n310));
  XNOR2_X1  g109(.A(G127gat), .B(G134gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n310), .B(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT75), .B1(new_n308), .B2(new_n312), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n298), .A2(new_n301), .B1(new_n291), .B2(new_n306), .ZN(new_n314));
  INV_X1    g113(.A(new_n311), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n310), .B(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n314), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n308), .A2(new_n312), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n313), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G225gat), .A2(G233gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n290), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n316), .B1(new_n308), .B2(KEYINPUT3), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT3), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n314), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n322), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT4), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n313), .A2(new_n328), .A3(new_n318), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n308), .A2(new_n312), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT4), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n327), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n323), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n313), .A2(KEYINPUT4), .A3(new_n318), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT76), .B1(new_n330), .B2(new_n328), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n313), .A2(KEYINPUT76), .A3(KEYINPUT4), .A4(new_n318), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n336), .A2(new_n290), .A3(new_n327), .A4(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G1gat), .B(G29gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(KEYINPUT0), .ZN(new_n340));
  XNOR2_X1  g139(.A(G57gat), .B(G85gat), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n340), .B(new_n341), .Z(new_n342));
  NAND3_X1  g141(.A1(new_n333), .A2(new_n338), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT77), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT6), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n344), .B1(new_n343), .B2(new_n345), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n342), .B1(new_n333), .B2(new_n338), .ZN(new_n348));
  NOR3_X1   g147(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(KEYINPUT6), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n289), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G15gat), .B(G43gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(KEYINPUT70), .ZN(new_n354));
  INV_X1    g153(.A(G71gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n354), .B(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(G99gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(G227gat), .ZN(new_n359));
  INV_X1    g158(.A(G233gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n280), .A2(new_n312), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n263), .A2(new_n316), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n358), .B1(new_n365), .B2(KEYINPUT33), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT32), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  OR2_X1    g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n363), .A2(new_n364), .A3(new_n362), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n370), .B(KEYINPUT34), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n363), .A2(new_n364), .ZN(new_n373));
  AOI221_X4 g172(.A(new_n367), .B1(KEYINPUT33), .B2(new_n358), .C1(new_n373), .C2(new_n361), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n369), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n213), .A2(KEYINPUT79), .A3(new_n214), .ZN(new_n377));
  OR2_X1    g176(.A1(new_n214), .A2(KEYINPUT79), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(new_n378), .A3(new_n268), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT80), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT3), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n377), .A2(new_n378), .A3(KEYINPUT80), .A4(new_n268), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n314), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n215), .B1(new_n326), .B2(new_n268), .ZN(new_n384));
  INV_X1    g183(.A(G228gat), .ZN(new_n385));
  OAI22_X1  g184(.A1(new_n383), .A2(new_n384), .B1(new_n385), .B2(new_n360), .ZN(new_n386));
  INV_X1    g185(.A(G22gat), .ZN(new_n387));
  INV_X1    g186(.A(new_n384), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT29), .B1(new_n213), .B2(new_n214), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n308), .B1(KEYINPUT3), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT81), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n385), .A2(new_n360), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT81), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n308), .B(new_n393), .C1(KEYINPUT3), .C2(new_n389), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n388), .A2(new_n391), .A3(new_n392), .A4(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n386), .A2(new_n387), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT82), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n386), .A2(new_n395), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(G22gat), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n386), .A2(KEYINPUT82), .A3(new_n387), .A4(new_n395), .ZN(new_n401));
  XNOR2_X1  g200(.A(G78gat), .B(G106gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT31), .B(G50gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n398), .A2(new_n400), .A3(new_n401), .A4(new_n404), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n404), .B(KEYINPUT78), .Z(new_n406));
  INV_X1    g205(.A(new_n396), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n387), .B1(new_n386), .B2(new_n395), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n366), .A2(new_n368), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n371), .B1(new_n411), .B2(new_n374), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n376), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT35), .B1(new_n352), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT89), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n343), .A2(new_n345), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n350), .B1(new_n416), .B2(new_n348), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT35), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n410), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  AND3_X1   g218(.A1(new_n285), .A2(new_n288), .A3(KEYINPUT83), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT83), .B1(new_n285), .B2(new_n288), .ZN(new_n421));
  NOR3_X1   g220(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n376), .A2(new_n412), .A3(KEYINPUT71), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT71), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n424), .B(new_n371), .C1(new_n411), .C2(new_n374), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  AOI22_X1  g225(.A1(new_n414), .A2(new_n415), .B1(new_n422), .B2(new_n426), .ZN(new_n427));
  OAI211_X1 g226(.A(KEYINPUT89), .B(KEYINPUT35), .C1(new_n352), .C2(new_n413), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n350), .B(new_n284), .C1(new_n416), .C2(new_n348), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT87), .B(KEYINPUT37), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n204), .B1(new_n286), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT37), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n431), .B1(new_n432), .B2(new_n286), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n429), .B1(new_n433), .B2(KEYINPUT38), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n283), .A2(new_n216), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT86), .ZN(new_n436));
  OAI22_X1  g235(.A1(new_n263), .A2(new_n274), .B1(new_n217), .B2(new_n267), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n436), .B1(new_n437), .B2(new_n215), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT37), .B1(new_n435), .B2(KEYINPUT86), .ZN(new_n440));
  OR2_X1    g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT88), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT38), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n441), .A2(new_n442), .A3(new_n443), .A4(new_n431), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n431), .A2(new_n443), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n439), .A2(new_n440), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT88), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n434), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n313), .A2(new_n318), .A3(new_n321), .A4(new_n319), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT85), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT39), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n451), .B1(new_n450), .B2(new_n449), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n324), .A2(new_n326), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n336), .A2(new_n453), .A3(new_n337), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n322), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(KEYINPUT84), .B(KEYINPUT39), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n456), .B(new_n342), .C1(new_n455), .C2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT40), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n348), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  OAI221_X1 g260(.A(new_n461), .B1(new_n460), .B2(new_n459), .C1(new_n420), .C2(new_n421), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n448), .A2(new_n462), .A3(new_n410), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT36), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n423), .A2(new_n464), .A3(new_n425), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n376), .A2(new_n412), .A3(KEYINPUT36), .ZN(new_n466));
  INV_X1    g265(.A(new_n410), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n465), .A2(new_n466), .B1(new_n467), .B2(new_n352), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n427), .A2(new_n428), .B1(new_n463), .B2(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(G15gat), .B(G22gat), .ZN(new_n470));
  OR2_X1    g269(.A1(new_n470), .A2(G1gat), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT92), .ZN(new_n472));
  AOI21_X1  g271(.A(G8gat), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT16), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n470), .B1(new_n474), .B2(G1gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n471), .B(new_n475), .C1(new_n472), .C2(G8gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(G43gat), .A2(G50gat), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(G43gat), .A2(G50gat), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT90), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OR2_X1    g282(.A1(G43gat), .A2(G50gat), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT90), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(new_n485), .A3(new_n480), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n483), .A2(new_n486), .A3(KEYINPUT15), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT14), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n488), .B1(G29gat), .B2(G36gat), .ZN(new_n489));
  INV_X1    g288(.A(G29gat), .ZN(new_n490));
  INV_X1    g289(.A(G36gat), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(new_n491), .A3(KEYINPUT14), .ZN(new_n492));
  XNOR2_X1  g291(.A(KEYINPUT91), .B(G36gat), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n489), .B(new_n492), .C1(new_n493), .C2(new_n490), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n484), .A2(new_n480), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n495), .A2(KEYINPUT15), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n487), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT15), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n498), .B1(new_n495), .B2(KEYINPUT90), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n492), .A2(new_n489), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n491), .A2(KEYINPUT91), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n491), .A2(KEYINPUT91), .ZN(new_n502));
  OAI21_X1  g301(.A(G29gat), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n499), .A2(new_n500), .A3(new_n486), .A4(new_n503), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n497), .A2(new_n504), .A3(KEYINPUT17), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT17), .B1(new_n497), .B2(new_n504), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n479), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(G229gat), .A2(G233gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n497), .A2(new_n504), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n510), .A2(new_n478), .A3(new_n477), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n507), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT18), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n507), .A2(KEYINPUT18), .A3(new_n511), .A4(new_n508), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n479), .A2(new_n509), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  XOR2_X1   g316(.A(new_n508), .B(KEYINPUT13), .Z(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n514), .A2(new_n515), .A3(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G113gat), .B(G141gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(G197gat), .ZN(new_n522));
  XOR2_X1   g321(.A(KEYINPUT11), .B(G169gat), .Z(new_n523));
  XNOR2_X1  g322(.A(new_n522), .B(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n524), .B(KEYINPUT12), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n520), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n514), .A2(new_n525), .A3(new_n515), .A4(new_n519), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT104), .ZN(new_n531));
  XOR2_X1   g330(.A(G99gat), .B(G106gat), .Z(new_n532));
  INV_X1    g331(.A(G106gat), .ZN(new_n533));
  OAI21_X1  g332(.A(KEYINPUT8), .B1(new_n357), .B2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(KEYINPUT97), .B(G92gat), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n534), .B1(new_n535), .B2(G85gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(G85gat), .A2(G92gat), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n537), .A2(KEYINPUT96), .A3(KEYINPUT7), .ZN(new_n538));
  NAND2_X1  g337(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n539), .A2(G85gat), .A3(G92gat), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n532), .B1(new_n536), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(G71gat), .A2(G78gat), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT9), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OR2_X1    g344(.A1(G57gat), .A2(G64gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(G57gat), .A2(G64gat), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n546), .A2(KEYINPUT93), .A3(new_n547), .ZN(new_n549));
  XNOR2_X1  g348(.A(G71gat), .B(G78gat), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AND2_X1   g350(.A1(G57gat), .A2(G64gat), .ZN(new_n552));
  NOR2_X1   g351(.A1(G57gat), .A2(G64gat), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AND2_X1   g353(.A1(G71gat), .A2(G78gat), .ZN(new_n555));
  NOR2_X1   g354(.A1(G71gat), .A2(G78gat), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n545), .B(new_n554), .C1(new_n557), .C2(KEYINPUT93), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT8), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n560), .B1(G99gat), .B2(G106gat), .ZN(new_n561));
  AND2_X1   g360(.A1(KEYINPUT97), .A2(G92gat), .ZN(new_n562));
  NOR2_X1   g361(.A1(KEYINPUT97), .A2(G92gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(G85gat), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n561), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n532), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n538), .A2(new_n540), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n542), .A2(new_n559), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT10), .ZN(new_n572));
  AND2_X1   g371(.A1(new_n551), .A2(new_n558), .ZN(new_n573));
  NOR3_X1   g372(.A1(new_n536), .A2(new_n541), .A3(new_n532), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n567), .B1(new_n566), .B2(new_n568), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT102), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n576), .A2(new_n577), .A3(new_n570), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n542), .A2(new_n569), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n579), .A2(KEYINPUT102), .A3(new_n573), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(KEYINPUT103), .B(KEYINPUT10), .Z(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n531), .B(new_n572), .C1(new_n581), .C2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G230gat), .A2(G233gat), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n583), .B1(new_n578), .B2(new_n580), .ZN(new_n586));
  INV_X1    g385(.A(new_n572), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT104), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n584), .A2(new_n585), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n585), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n581), .A2(new_n590), .ZN(new_n591));
  XOR2_X1   g390(.A(G120gat), .B(G148gat), .Z(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT105), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT106), .ZN(new_n594));
  XNOR2_X1  g393(.A(G176gat), .B(G204gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  AND2_X1   g395(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n589), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT107), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(new_n591), .ZN(new_n601));
  INV_X1    g400(.A(new_n596), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n599), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AOI211_X1 g402(.A(KEYINPUT107), .B(new_n596), .C1(new_n600), .C2(new_n591), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n598), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT21), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n573), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G127gat), .B(G155gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n611), .B(KEYINPUT94), .Z(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n610), .A2(new_n613), .ZN(new_n615));
  XNOR2_X1  g414(.A(G183gat), .B(G211gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT95), .ZN(new_n617));
  OR3_X1    g416(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n617), .B1(new_n614), .B2(new_n615), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n479), .B1(new_n607), .B2(new_n573), .ZN(new_n621));
  XOR2_X1   g420(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n618), .A2(new_n623), .A3(new_n619), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT98), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n542), .A2(new_n628), .A3(new_n569), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n628), .B1(new_n542), .B2(new_n569), .ZN(new_n630));
  OAI22_X1  g429(.A1(new_n505), .A2(new_n506), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(G232gat), .A2(G233gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(KEYINPUT41), .ZN(new_n633));
  XOR2_X1   g432(.A(G190gat), .B(G218gat), .Z(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT99), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT100), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n579), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n637), .B1(new_n510), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n631), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n635), .A2(new_n636), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT101), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n632), .A2(KEYINPUT41), .ZN(new_n645));
  XNOR2_X1  g444(.A(G134gat), .B(G162gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n631), .A2(new_n641), .A3(new_n639), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n643), .A2(new_n644), .A3(new_n647), .A4(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n647), .B(KEYINPUT101), .ZN(new_n650));
  AND3_X1   g449(.A1(new_n631), .A2(new_n641), .A3(new_n639), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n641), .B1(new_n631), .B2(new_n639), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n606), .A2(new_n627), .A3(new_n654), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n469), .A2(new_n530), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n349), .A2(new_n351), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g458(.A1(new_n420), .A2(new_n421), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT16), .B(G8gat), .Z(new_n662));
  NAND3_X1  g461(.A1(new_n656), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n656), .ZN(new_n664));
  OAI21_X1  g463(.A(G8gat), .B1(new_n664), .B2(new_n660), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n663), .ZN(new_n666));
  MUX2_X1   g465(.A(new_n663), .B(new_n666), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g466(.A1(new_n465), .A2(new_n466), .ZN(new_n668));
  OAI21_X1  g467(.A(G15gat), .B1(new_n664), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n426), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n670), .A2(G15gat), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n669), .B1(new_n664), .B2(new_n671), .ZN(G1326gat));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n467), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT43), .B(G22gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1327gat));
  NOR2_X1   g474(.A1(new_n469), .A2(new_n530), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n627), .A2(new_n605), .A3(new_n654), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n676), .A2(new_n490), .A3(new_n657), .A4(new_n677), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n678), .A2(KEYINPUT108), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(KEYINPUT108), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT45), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n679), .A2(KEYINPUT45), .A3(new_n680), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n685), .B1(new_n469), .B2(new_n654), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n463), .A2(new_n468), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n414), .A2(new_n415), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n422), .A2(new_n426), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n688), .A2(new_n428), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n654), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(KEYINPUT44), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n686), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n627), .A2(new_n530), .A3(new_n605), .ZN(new_n696));
  AND3_X1   g495(.A1(new_n695), .A2(new_n657), .A3(new_n696), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n683), .B(new_n684), .C1(new_n490), .C2(new_n697), .ZN(G1328gat));
  AND2_X1   g497(.A1(new_n676), .A2(new_n677), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n699), .A2(new_n493), .A3(new_n661), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT46), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n695), .A2(new_n661), .A3(new_n696), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT109), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OAI22_X1  g504(.A1(new_n703), .A2(new_n704), .B1(new_n501), .B2(new_n502), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n702), .B1(new_n705), .B2(new_n706), .ZN(G1329gat));
  NOR2_X1   g506(.A1(new_n670), .A2(G43gat), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n699), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT110), .ZN(new_n710));
  AOI21_X1  g509(.A(KEYINPUT47), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n668), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n686), .A2(new_n693), .A3(new_n712), .A4(new_n696), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(G43gat), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n709), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n711), .B(new_n715), .ZN(G1330gat));
  NOR2_X1   g515(.A1(new_n410), .A2(G50gat), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n699), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n686), .A2(new_n693), .A3(new_n467), .A4(new_n696), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT112), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(G50gat), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n719), .A2(new_n720), .ZN(new_n723));
  OAI211_X1 g522(.A(KEYINPUT48), .B(new_n718), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT111), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n719), .A2(G50gat), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n718), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT48), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n725), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI211_X1 g528(.A(KEYINPUT111), .B(KEYINPUT48), .C1(new_n726), .C2(new_n718), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n724), .B1(new_n729), .B2(new_n730), .ZN(G1331gat));
  AOI211_X1 g530(.A(new_n529), .B(new_n692), .C1(new_n625), .C2(new_n626), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n732), .A2(new_n605), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n733), .B(KEYINPUT113), .Z(new_n734));
  OAI21_X1  g533(.A(KEYINPUT114), .B1(new_n469), .B2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT114), .ZN(new_n736));
  INV_X1    g535(.A(new_n734), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n691), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n657), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g540(.A(new_n660), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT115), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n744), .B(new_n745), .Z(G1333gat));
  NAND3_X1  g545(.A1(new_n735), .A2(new_n738), .A3(new_n426), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT116), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT116), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n735), .A2(new_n738), .A3(new_n749), .A4(new_n426), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n748), .A2(new_n355), .A3(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n739), .A2(G71gat), .A3(new_n712), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT50), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n751), .A2(new_n752), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(G1334gat));
  NAND2_X1  g556(.A1(new_n739), .A2(new_n467), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(G78gat), .ZN(G1335gat));
  INV_X1    g558(.A(new_n657), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n760), .A2(G85gat), .A3(new_n606), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n627), .A2(new_n529), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n469), .A2(new_n654), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n763), .B1(new_n764), .B2(KEYINPUT117), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT117), .B1(new_n691), .B2(new_n692), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT51), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n691), .A2(KEYINPUT117), .A3(new_n692), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n762), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT51), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n770), .A2(new_n771), .A3(new_n766), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n761), .B1(new_n768), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n763), .A2(new_n606), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n694), .A2(new_n760), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n773), .B1(new_n565), .B2(new_n776), .ZN(G1336gat));
  NOR3_X1   g576(.A1(new_n660), .A2(G92gat), .A3(new_n606), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(new_n768), .B2(new_n772), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n686), .A2(new_n693), .A3(new_n661), .A4(new_n774), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n535), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n779), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n778), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n765), .A2(KEYINPUT51), .A3(new_n767), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n771), .B1(new_n770), .B2(new_n766), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n782), .ZN(new_n788));
  OAI21_X1  g587(.A(KEYINPUT52), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n783), .A2(new_n789), .ZN(G1337gat));
  NOR3_X1   g589(.A1(new_n670), .A2(G99gat), .A3(new_n606), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n791), .B1(new_n768), .B2(new_n772), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n694), .A2(new_n668), .A3(new_n775), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n792), .B1(new_n357), .B2(new_n793), .ZN(G1338gat));
  NOR3_X1   g593(.A1(new_n410), .A2(new_n606), .A3(G106gat), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n795), .B1(new_n768), .B2(new_n772), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n686), .A2(new_n693), .A3(new_n467), .A4(new_n774), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(G106gat), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n796), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n795), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(new_n785), .B2(new_n786), .ZN(new_n802));
  INV_X1    g601(.A(new_n799), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT53), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n800), .A2(new_n804), .ZN(G1339gat));
  NAND2_X1  g604(.A1(new_n732), .A2(new_n606), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT118), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n732), .A2(KEYINPUT118), .A3(new_n606), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n627), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n586), .A2(new_n587), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n812), .B1(new_n813), .B2(new_n590), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n589), .A2(new_n814), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n812), .B(new_n585), .C1(new_n586), .C2(new_n587), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n602), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n815), .A2(KEYINPUT55), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n598), .ZN(new_n820));
  INV_X1    g619(.A(new_n518), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n511), .A2(new_n516), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n508), .B1(new_n507), .B2(new_n511), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n524), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AND4_X1   g623(.A1(new_n528), .A2(new_n649), .A3(new_n653), .A4(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n817), .B1(new_n589), .B2(new_n814), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n825), .B1(new_n826), .B2(KEYINPUT55), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n820), .A2(new_n827), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n528), .A2(new_n824), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n605), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n529), .B1(new_n826), .B2(KEYINPUT55), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n830), .B1(new_n820), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n828), .B1(new_n832), .B2(new_n654), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n811), .B1(new_n833), .B2(KEYINPUT119), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT119), .ZN(new_n835));
  AOI211_X1 g634(.A(new_n835), .B(new_n828), .C1(new_n654), .C2(new_n832), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n810), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT120), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n839), .B(new_n810), .C1(new_n834), .C2(new_n836), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n841), .A2(new_n657), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n661), .A2(new_n413), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(new_n529), .A3(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(G113gat), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n670), .A2(new_n467), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n841), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n660), .A2(new_n657), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n530), .A2(new_n845), .ZN(new_n850));
  AOI22_X1  g649(.A1(new_n844), .A2(new_n845), .B1(new_n849), .B2(new_n850), .ZN(G1340gat));
  NAND3_X1  g650(.A1(new_n842), .A2(new_n605), .A3(new_n843), .ZN(new_n852));
  INV_X1    g651(.A(G120gat), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n606), .A2(new_n853), .ZN(new_n854));
  AOI22_X1  g653(.A1(new_n852), .A2(new_n853), .B1(new_n849), .B2(new_n854), .ZN(G1341gat));
  INV_X1    g654(.A(new_n849), .ZN(new_n856));
  OAI21_X1  g655(.A(G127gat), .B1(new_n856), .B2(new_n811), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n843), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n811), .A2(G127gat), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(G1342gat));
  OR2_X1    g659(.A1(new_n654), .A2(G134gat), .ZN(new_n861));
  XOR2_X1   g660(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  OR3_X1    g662(.A1(new_n858), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n863), .B1(new_n858), .B2(new_n861), .ZN(new_n865));
  OAI21_X1  g664(.A(G134gat), .B1(new_n856), .B2(new_n654), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(G1343gat));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n841), .A2(new_n868), .A3(new_n467), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n668), .A2(new_n657), .A3(new_n660), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n833), .A2(new_n627), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n810), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n467), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n870), .B1(new_n873), .B2(KEYINPUT57), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n869), .A2(new_n529), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n292), .A2(new_n293), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n712), .A2(new_n410), .A3(new_n661), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n842), .A2(new_n295), .A3(new_n529), .A4(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT58), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT58), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n877), .A2(new_n882), .A3(new_n879), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(new_n883), .ZN(G1344gat));
  NAND4_X1  g683(.A1(new_n842), .A2(new_n304), .A3(new_n605), .A4(new_n878), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n467), .A2(new_n868), .ZN(new_n887));
  XOR2_X1   g686(.A(new_n806), .B(KEYINPUT123), .Z(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n888), .B2(new_n871), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n870), .A2(KEYINPUT122), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT122), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n668), .A2(new_n891), .A3(new_n657), .A4(new_n660), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n890), .A2(new_n605), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n838), .A2(new_n467), .A3(new_n840), .ZN(new_n894));
  AOI211_X1 g693(.A(new_n889), .B(new_n893), .C1(new_n894), .C2(KEYINPUT57), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n304), .B1(new_n895), .B2(KEYINPUT124), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT124), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n894), .A2(KEYINPUT57), .ZN(new_n898));
  INV_X1    g697(.A(new_n889), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n897), .B1(new_n900), .B2(new_n893), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n886), .B1(new_n896), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n886), .A2(G148gat), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n869), .A2(new_n874), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n903), .B1(new_n904), .B2(new_n605), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n885), .B1(new_n902), .B2(new_n905), .ZN(G1345gat));
  NAND4_X1  g705(.A1(new_n842), .A2(new_n300), .A3(new_n627), .A4(new_n878), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n904), .A2(new_n627), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n908), .B2(new_n300), .ZN(G1346gat));
  NAND3_X1  g708(.A1(new_n842), .A2(new_n692), .A3(new_n878), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n654), .A2(new_n299), .ZN(new_n911));
  AOI22_X1  g710(.A1(new_n299), .A2(new_n910), .B1(new_n904), .B2(new_n911), .ZN(G1347gat));
  NOR2_X1   g711(.A1(new_n660), .A2(new_n657), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n838), .A2(new_n840), .A3(new_n846), .A4(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(G169gat), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n914), .A2(new_n915), .A3(new_n530), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n838), .A2(new_n840), .ZN(new_n917));
  INV_X1    g716(.A(new_n913), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n917), .A2(new_n413), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(new_n529), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n916), .B1(new_n920), .B2(new_n915), .ZN(G1348gat));
  AOI21_X1  g720(.A(G176gat), .B1(new_n919), .B2(new_n605), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n922), .A2(KEYINPUT125), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(KEYINPUT125), .ZN(new_n924));
  INV_X1    g723(.A(new_n914), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n605), .A2(G176gat), .ZN(new_n926));
  AOI22_X1  g725(.A1(new_n923), .A2(new_n924), .B1(new_n925), .B2(new_n926), .ZN(G1349gat));
  NAND3_X1  g726(.A1(new_n919), .A2(new_n218), .A3(new_n627), .ZN(new_n928));
  OAI21_X1  g727(.A(KEYINPUT126), .B1(new_n914), .B2(new_n811), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(G183gat), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n914), .A2(KEYINPUT126), .A3(new_n811), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g732(.A1(new_n919), .A2(new_n219), .A3(new_n692), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n925), .A2(new_n692), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n935), .A2(new_n936), .A3(G190gat), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n936), .B1(new_n935), .B2(G190gat), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n934), .B1(new_n938), .B2(new_n939), .ZN(G1351gat));
  AOI21_X1  g739(.A(new_n889), .B1(new_n894), .B2(KEYINPUT57), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n712), .A2(new_n918), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(G197gat), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n943), .A2(new_n944), .A3(new_n530), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n841), .A2(new_n467), .A3(new_n942), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(G197gat), .B1(new_n947), .B2(new_n529), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n945), .A2(new_n948), .ZN(G1352gat));
  NOR3_X1   g748(.A1(new_n946), .A2(G204gat), .A3(new_n606), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT62), .ZN(new_n951));
  OAI21_X1  g750(.A(G204gat), .B1(new_n943), .B2(new_n606), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1353gat));
  NAND3_X1  g752(.A1(new_n947), .A2(new_n207), .A3(new_n627), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT127), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n941), .A2(new_n627), .A3(new_n942), .ZN(new_n956));
  AND4_X1   g755(.A1(new_n955), .A2(new_n956), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT63), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n207), .B1(KEYINPUT127), .B2(new_n958), .ZN(new_n959));
  AOI22_X1  g758(.A1(new_n956), .A2(new_n959), .B1(new_n955), .B2(KEYINPUT63), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n954), .B1(new_n957), .B2(new_n960), .ZN(G1354gat));
  OAI21_X1  g760(.A(G218gat), .B1(new_n943), .B2(new_n654), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n947), .A2(new_n208), .A3(new_n692), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(G1355gat));
endmodule


