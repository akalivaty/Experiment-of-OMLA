//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993;
  INV_X1    g000(.A(KEYINPUT76), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT26), .B(G101), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT72), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT70), .ZN(new_n192));
  INV_X1    g006(.A(G237), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT70), .A2(G237), .ZN(new_n195));
  AOI21_X1  g009(.A(G953), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n191), .B1(new_n196), .B2(G210), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(new_n191), .A3(G210), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n190), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n199), .ZN(new_n201));
  INV_X1    g015(.A(new_n190), .ZN(new_n202));
  NOR3_X1   g016(.A1(new_n201), .A2(new_n197), .A3(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n189), .B1(new_n200), .B2(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n202), .B1(new_n201), .B2(new_n197), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n198), .A2(new_n199), .A3(new_n190), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(new_n188), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(new_n208), .B(KEYINPUT74), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT28), .ZN(new_n210));
  INV_X1    g024(.A(G137), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G134), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT11), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n211), .A2(KEYINPUT11), .A3(G134), .ZN(new_n215));
  INV_X1    g029(.A(G134), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G137), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n214), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  XOR2_X1   g032(.A(KEYINPUT66), .B(G131), .Z(new_n219));
  NOR2_X1   g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n218), .A2(G131), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n224));
  AND2_X1   g038(.A1(KEYINPUT0), .A2(G128), .ZN(new_n225));
  INV_X1    g039(.A(G146), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G143), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT64), .ZN(new_n228));
  INV_X1    g042(.A(G143), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n228), .B1(new_n229), .B2(G146), .ZN(new_n230));
  NOR3_X1   g044(.A1(new_n226), .A2(KEYINPUT64), .A3(G143), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n225), .B(new_n227), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT65), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n229), .A2(G146), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT64), .B1(new_n226), .B2(G143), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n228), .A2(new_n229), .A3(G146), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(KEYINPUT65), .A3(new_n225), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(G143), .B(G146), .ZN(new_n241));
  NOR2_X1   g055(.A1(KEYINPUT0), .A2(G128), .ZN(new_n242));
  NOR3_X1   g056(.A1(new_n241), .A2(new_n225), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n224), .B1(new_n240), .B2(new_n244), .ZN(new_n245));
  AOI211_X1 g059(.A(KEYINPUT69), .B(new_n243), .C1(new_n234), .C2(new_n239), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n223), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT75), .ZN(new_n248));
  INV_X1    g062(.A(G131), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n249), .B1(new_n212), .B2(new_n217), .ZN(new_n250));
  XOR2_X1   g064(.A(new_n250), .B(KEYINPUT67), .Z(new_n251));
  INV_X1    g065(.A(G128), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n252), .B1(new_n227), .B2(KEYINPUT1), .ZN(new_n253));
  OR2_X1    g067(.A1(new_n253), .A2(new_n241), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n238), .A2(new_n253), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n251), .A2(new_n256), .A3(new_n221), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n247), .A2(new_n248), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G119), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT68), .B1(new_n259), .B2(G116), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT68), .ZN(new_n261));
  INV_X1    g075(.A(G116), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(new_n262), .A3(G119), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n260), .A2(new_n263), .B1(G116), .B2(new_n259), .ZN(new_n264));
  XOR2_X1   g078(.A(KEYINPUT2), .B(G113), .Z(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n258), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n248), .B1(new_n247), .B2(new_n257), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n210), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n247), .A2(new_n267), .A3(new_n257), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n223), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n236), .A2(new_n237), .ZN(new_n274));
  AND4_X1   g088(.A1(KEYINPUT65), .A2(new_n274), .A3(new_n225), .A4(new_n227), .ZN(new_n275));
  AOI21_X1  g089(.A(KEYINPUT65), .B1(new_n238), .B2(new_n225), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n244), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n257), .B1(new_n273), .B2(new_n277), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n278), .A2(new_n266), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT28), .B1(new_n272), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n209), .B1(new_n270), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n271), .A2(new_n208), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT73), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n247), .A2(KEYINPUT30), .A3(new_n257), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT30), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n278), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n284), .A2(new_n266), .A3(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT73), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n271), .A2(new_n288), .A3(new_n208), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n283), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT31), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n283), .A2(KEYINPUT31), .A3(new_n287), .A4(new_n289), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n281), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(G472), .A2(G902), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n187), .B(KEYINPUT32), .C1(new_n294), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n270), .A2(new_n280), .ZN(new_n298));
  INV_X1    g112(.A(new_n209), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n271), .A2(new_n288), .A3(new_n208), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n288), .B1(new_n271), .B2(new_n208), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(KEYINPUT31), .B1(new_n303), .B2(new_n287), .ZN(new_n304));
  INV_X1    g118(.A(new_n293), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n300), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT76), .B1(new_n306), .B2(new_n295), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n297), .B1(new_n307), .B2(KEYINPUT32), .ZN(new_n308));
  INV_X1    g122(.A(new_n257), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n277), .A2(KEYINPUT69), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n243), .B1(new_n234), .B2(new_n239), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n224), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n309), .B1(new_n313), .B2(new_n223), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n266), .B1(new_n314), .B2(new_n248), .ZN(new_n315));
  INV_X1    g129(.A(new_n269), .ZN(new_n316));
  AOI21_X1  g130(.A(KEYINPUT28), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n267), .B1(new_n247), .B2(new_n257), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n210), .B1(new_n319), .B2(new_n271), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT77), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n321), .A2(new_n322), .A3(KEYINPUT29), .A4(new_n208), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT29), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n287), .A2(new_n271), .ZN(new_n325));
  INV_X1    g139(.A(new_n208), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n324), .B(new_n327), .C1(new_n298), .C2(new_n299), .ZN(new_n328));
  INV_X1    g142(.A(G902), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT28), .B1(new_n272), .B2(new_n318), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n270), .A2(new_n330), .A3(KEYINPUT29), .A4(new_n208), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT77), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n323), .A2(new_n328), .A3(new_n329), .A4(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G472), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n308), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G469), .ZN(new_n336));
  INV_X1    g150(.A(G953), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G227), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(KEYINPUT84), .ZN(new_n339));
  XNOR2_X1  g153(.A(G110), .B(G140), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n339), .B(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G104), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT3), .B1(new_n343), .B2(G107), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT3), .ZN(new_n345));
  INV_X1    g159(.A(G107), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n346), .A3(G104), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n343), .A2(G107), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n344), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT85), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n344), .A2(new_n347), .A3(KEYINPUT85), .A4(new_n348), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(G101), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G101), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n344), .A2(new_n347), .A3(new_n354), .A4(new_n348), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n353), .A2(KEYINPUT4), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT86), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT86), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n353), .A2(new_n358), .A3(KEYINPUT4), .A4(new_n355), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT4), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n351), .A2(new_n361), .A3(G101), .A4(new_n352), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n360), .A2(new_n313), .A3(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n343), .A2(G107), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n346), .A2(G104), .ZN(new_n365));
  OAI21_X1  g179(.A(G101), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n355), .A2(new_n366), .ZN(new_n367));
  OR2_X1    g181(.A1(new_n238), .A2(new_n253), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n367), .B1(new_n368), .B2(new_n255), .ZN(new_n369));
  OR2_X1    g183(.A1(new_n369), .A2(KEYINPUT10), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT87), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n367), .B(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n373));
  INV_X1    g187(.A(new_n256), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n363), .A2(new_n370), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n223), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n363), .A2(new_n273), .A3(new_n370), .A4(new_n376), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n342), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n367), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n256), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n223), .B1(new_n382), .B2(new_n369), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT12), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g199(.A(KEYINPUT12), .B(new_n223), .C1(new_n382), .C2(new_n369), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT88), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT88), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n385), .A2(new_n389), .A3(new_n386), .ZN(new_n390));
  AND4_X1   g204(.A1(new_n379), .A2(new_n388), .A3(new_n342), .A4(new_n390), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n336), .B(new_n329), .C1(new_n380), .C2(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n336), .A2(new_n329), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n378), .A2(new_n379), .A3(new_n342), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n379), .A2(new_n387), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n341), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(new_n397), .A3(G469), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n392), .A2(new_n394), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G221), .ZN(new_n400));
  XOR2_X1   g214(.A(KEYINPUT9), .B(G234), .Z(new_n401));
  AOI21_X1  g215(.A(new_n400), .B1(new_n401), .B2(new_n329), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(G214), .B1(G237), .B2(G902), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n266), .A2(new_n362), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n407), .B1(new_n357), .B2(new_n359), .ZN(new_n408));
  XOR2_X1   g222(.A(G110), .B(G122), .Z(new_n409));
  NAND2_X1  g223(.A1(new_n264), .A2(new_n265), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n264), .A2(KEYINPUT5), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n259), .A2(G116), .ZN(new_n413));
  OAI21_X1  g227(.A(G113), .B1(new_n413), .B2(KEYINPUT5), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n410), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n372), .A2(new_n415), .ZN(new_n416));
  OR3_X1    g230(.A1(new_n408), .A2(new_n409), .A3(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n409), .B1(new_n408), .B2(new_n416), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(KEYINPUT6), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G125), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n374), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n421), .B1(new_n311), .B2(new_n420), .ZN(new_n422));
  INV_X1    g236(.A(G224), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(G953), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n422), .B(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT6), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n426), .B(new_n409), .C1(new_n408), .C2(new_n416), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n419), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT7), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n424), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n422), .B1(KEYINPUT91), .B2(new_n424), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n414), .B(KEYINPUT89), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n411), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(new_n410), .A3(new_n381), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT90), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n415), .A2(new_n367), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n433), .A2(KEYINPUT90), .A3(new_n410), .A4(new_n381), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  XOR2_X1   g253(.A(new_n409), .B(KEYINPUT8), .Z(new_n440));
  AOI22_X1  g254(.A1(new_n430), .A2(new_n431), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n441), .B(new_n417), .C1(new_n430), .C2(new_n431), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n428), .A2(new_n442), .A3(new_n329), .ZN(new_n443));
  OAI21_X1  g257(.A(G210), .B1(G237), .B2(G902), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n428), .A2(new_n442), .A3(new_n329), .A4(new_n444), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n406), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G140), .ZN(new_n449));
  AOI21_X1  g263(.A(KEYINPUT16), .B1(new_n449), .B2(G125), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(KEYINPUT79), .A2(G125), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(new_n449), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT16), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n451), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n455), .A2(G146), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n452), .B(G140), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT16), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n226), .B1(new_n458), .B2(new_n451), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n195), .ZN(new_n461));
  NOR2_X1   g275(.A1(KEYINPUT70), .A2(G237), .ZN(new_n462));
  OAI211_X1 g276(.A(G214), .B(new_n337), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(KEYINPUT92), .A2(G143), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(KEYINPUT92), .A2(G143), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n464), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  OAI211_X1 g281(.A(KEYINPUT17), .B(new_n219), .C1(new_n465), .C2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n463), .A2(new_n464), .ZN(new_n469));
  INV_X1    g283(.A(new_n219), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n463), .A2(new_n466), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n469), .B(new_n470), .C1(new_n471), .C2(new_n464), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n219), .B1(new_n465), .B2(new_n467), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n460), .B(new_n468), .C1(new_n474), .C2(KEYINPUT17), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n457), .A2(G146), .ZN(new_n476));
  XNOR2_X1  g290(.A(G125), .B(G140), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n226), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT18), .ZN(new_n480));
  NOR4_X1   g294(.A1(new_n465), .A2(new_n467), .A3(new_n480), .A4(new_n249), .ZN(new_n481));
  OAI22_X1  g295(.A1(new_n465), .A2(new_n467), .B1(new_n480), .B2(new_n249), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n479), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(G113), .B(G122), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n485), .B(new_n343), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n475), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n486), .B1(new_n475), .B2(new_n484), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n329), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT93), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT93), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n492), .B(new_n329), .C1(new_n488), .C2(new_n489), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n491), .A2(G475), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n486), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n465), .A2(new_n467), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(KEYINPUT18), .A3(G131), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n497), .A2(new_n482), .B1(new_n478), .B2(new_n476), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n455), .A2(G146), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT19), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n477), .A2(new_n500), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n501), .B(new_n226), .C1(new_n453), .C2(new_n500), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n503), .B1(new_n473), .B2(new_n472), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n495), .B1(new_n498), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n487), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G475), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(new_n507), .A3(new_n329), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT20), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT20), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n506), .A2(new_n510), .A3(new_n507), .A4(new_n329), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n494), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n401), .A2(G217), .A3(new_n337), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n262), .A2(G122), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n346), .B1(new_n516), .B2(KEYINPUT14), .ZN(new_n517));
  XNOR2_X1  g331(.A(G116), .B(G122), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n517), .B1(new_n519), .B2(KEYINPUT14), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n229), .A2(G128), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n252), .A2(G143), .ZN(new_n522));
  OAI21_X1  g336(.A(G134), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n252), .A2(G143), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n229), .A2(G128), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n525), .A3(new_n216), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n520), .B(new_n527), .C1(G107), .C2(new_n519), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT94), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT13), .B1(new_n229), .B2(G128), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n529), .B1(new_n530), .B2(new_n521), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n524), .B1(new_n522), .B2(KEYINPUT13), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT13), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT94), .B1(new_n525), .B2(new_n533), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n531), .B(G134), .C1(new_n532), .C2(new_n534), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n518), .B(new_n346), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(new_n536), .A3(new_n526), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT95), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n528), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n538), .B1(new_n528), .B2(new_n537), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n515), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n528), .A2(new_n537), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n514), .B1(new_n542), .B2(KEYINPUT95), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n329), .ZN(new_n545));
  INV_X1    g359(.A(G478), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n546), .A2(KEYINPUT15), .ZN(new_n547));
  XOR2_X1   g361(.A(new_n545), .B(new_n547), .Z(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n337), .A2(G952), .ZN(new_n550));
  INV_X1    g364(.A(G234), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n550), .B1(new_n551), .B2(new_n193), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  XOR2_X1   g367(.A(KEYINPUT21), .B(G898), .Z(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(KEYINPUT96), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  AOI211_X1 g370(.A(new_n329), .B(new_n337), .C1(G234), .C2(G237), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n553), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n513), .A2(new_n549), .A3(new_n558), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n404), .A2(new_n448), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n252), .A2(G119), .ZN(new_n561));
  OR2_X1    g375(.A1(new_n561), .A2(KEYINPUT23), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n259), .A2(G128), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n561), .A2(new_n563), .A3(KEYINPUT23), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(G110), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n563), .A2(KEYINPUT78), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT78), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(new_n259), .A3(G128), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n568), .A2(new_n570), .B1(G119), .B2(new_n252), .ZN(new_n571));
  XOR2_X1   g385(.A(KEYINPUT24), .B(G110), .Z(new_n572));
  OAI211_X1 g386(.A(new_n567), .B(KEYINPUT80), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT80), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n571), .A2(new_n572), .ZN(new_n575));
  AOI21_X1  g389(.A(G110), .B1(new_n562), .B2(new_n564), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n573), .A2(new_n577), .A3(new_n499), .A4(new_n478), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n571), .A2(new_n572), .ZN(new_n579));
  OAI221_X1 g393(.A(new_n579), .B1(new_n566), .B2(new_n565), .C1(new_n456), .C2(new_n459), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT22), .B(G137), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n400), .A2(new_n551), .A3(G953), .ZN(new_n583));
  XOR2_X1   g397(.A(new_n582), .B(new_n583), .Z(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n578), .A2(new_n580), .A3(new_n584), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(new_n329), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(KEYINPUT81), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT25), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n588), .A2(KEYINPUT81), .A3(KEYINPUT25), .ZN(new_n592));
  INV_X1    g406(.A(G217), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n593), .B1(G234), .B2(new_n329), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT82), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n591), .A2(new_n592), .A3(KEYINPUT82), .A4(new_n594), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n594), .A2(G902), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(KEYINPUT83), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n586), .A2(new_n587), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n597), .A2(new_n598), .A3(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n335), .A2(new_n560), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G101), .ZN(G3));
  OAI21_X1  g419(.A(G472), .B1(new_n294), .B2(G902), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT97), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n448), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n399), .A2(new_n403), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n609), .A2(new_n610), .A3(new_n602), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n292), .A2(new_n293), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n296), .B1(new_n612), .B2(new_n300), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n608), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(KEYINPUT33), .B1(new_n541), .B2(new_n543), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n542), .B1(KEYINPUT98), .B2(new_n514), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n514), .A2(KEYINPUT98), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n528), .B2(new_n537), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT33), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n617), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(KEYINPUT99), .B1(new_n616), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT99), .ZN(new_n623));
  OR2_X1    g437(.A1(new_n617), .A2(new_n619), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n623), .B1(new_n624), .B2(new_n620), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n622), .A2(G478), .A3(new_n625), .A4(new_n329), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n545), .A2(new_n546), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n513), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n629), .A2(new_n558), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n615), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(G104), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  NAND2_X1  g448(.A1(new_n512), .A2(KEYINPUT101), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT101), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n509), .A2(new_n636), .A3(new_n511), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n494), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n639), .A2(new_n558), .A3(new_n548), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n615), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT35), .B(G107), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G9));
  NOR2_X1   g457(.A1(new_n585), .A2(KEYINPUT36), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n581), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n600), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT102), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n597), .A2(new_n598), .A3(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT103), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n560), .A2(new_n608), .A3(new_n614), .A4(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT104), .B(KEYINPUT105), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT37), .B(G110), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G12));
  NOR2_X1   g470(.A1(new_n609), .A2(new_n610), .ZN(new_n657));
  INV_X1    g471(.A(G900), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n557), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n552), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n639), .A2(new_n548), .A3(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n335), .A2(new_n657), .A3(new_n651), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  INV_X1    g478(.A(new_n649), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n660), .B(KEYINPUT39), .Z(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n404), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n665), .B1(new_n668), .B2(KEYINPUT40), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n209), .B1(new_n271), .B2(new_n319), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n287), .B2(new_n303), .ZN(new_n671));
  OAI21_X1  g485(.A(G472), .B1(new_n671), .B2(G902), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n308), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  AOI211_X1 g488(.A(new_n669), .B(new_n674), .C1(KEYINPUT40), .C2(new_n668), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n446), .A2(new_n447), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n676), .B(KEYINPUT38), .Z(new_n677));
  NOR2_X1   g491(.A1(new_n677), .A2(new_n406), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n513), .A2(new_n549), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n675), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(KEYINPUT106), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT106), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n675), .A2(new_n683), .A3(new_n678), .A4(new_n680), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G143), .ZN(G45));
  AOI221_X4 g500(.A(new_n661), .B1(new_n626), .B2(new_n627), .C1(new_n494), .C2(new_n512), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n335), .A2(new_n657), .A3(new_n651), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  NAND2_X1  g503(.A1(new_n392), .A2(KEYINPUT107), .ZN(new_n690));
  INV_X1    g504(.A(new_n379), .ZN(new_n691));
  INV_X1    g505(.A(new_n362), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n310), .B2(new_n312), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n375), .B1(new_n693), .B2(new_n360), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n273), .B1(new_n694), .B2(new_n370), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n341), .B1(new_n691), .B2(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n379), .A2(new_n388), .A3(new_n342), .A4(new_n390), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n336), .B1(new_n698), .B2(new_n329), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n690), .A2(new_n699), .ZN(new_n700));
  AOI211_X1 g514(.A(KEYINPUT107), .B(new_n336), .C1(new_n698), .C2(new_n329), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n448), .B(new_n403), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n335), .A2(new_n703), .A3(new_n603), .A4(new_n630), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT41), .B(G113), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G15));
  NAND4_X1  g520(.A1(new_n335), .A2(new_n703), .A3(new_n603), .A4(new_n640), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G116), .ZN(G18));
  NAND4_X1  g522(.A1(new_n335), .A2(new_n703), .A3(new_n559), .A4(new_n651), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G119), .ZN(G21));
  OAI21_X1  g524(.A(new_n612), .B1(new_n209), .B2(new_n321), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n295), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n606), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n602), .ZN(new_n714));
  INV_X1    g528(.A(new_n700), .ZN(new_n715));
  INV_X1    g529(.A(new_n701), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n402), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n558), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n609), .A2(new_n679), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n714), .A2(new_n717), .A3(new_n718), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G122), .ZN(G24));
  NAND3_X1  g535(.A1(new_n513), .A2(new_n628), .A3(new_n660), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n713), .A2(new_n665), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n703), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G125), .ZN(G27));
  INV_X1    g539(.A(KEYINPUT32), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n726), .B1(new_n613), .B2(KEYINPUT76), .ZN(new_n727));
  AOI22_X1  g541(.A1(new_n727), .A2(new_n297), .B1(new_n333), .B2(G472), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n446), .A2(new_n405), .A3(new_n447), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n729), .A2(new_n687), .A3(new_n403), .A4(new_n399), .ZN(new_n730));
  NOR4_X1   g544(.A1(new_n728), .A2(new_n730), .A3(KEYINPUT42), .A4(new_n602), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT42), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n613), .A2(new_n726), .ZN(new_n733));
  OAI21_X1  g547(.A(KEYINPUT32), .B1(new_n294), .B2(new_n296), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n602), .B1(new_n735), .B2(new_n334), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n446), .A2(new_n405), .A3(new_n447), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n610), .A2(new_n737), .A3(new_n722), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n732), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g553(.A(KEYINPUT108), .B1(new_n731), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n726), .B1(new_n306), .B2(new_n295), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n294), .A2(KEYINPUT32), .A3(new_n296), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n334), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n738), .A3(new_n603), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(KEYINPUT42), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n335), .A2(new_n732), .A3(new_n603), .A4(new_n738), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT108), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n740), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G131), .ZN(G33));
  NOR2_X1   g564(.A1(new_n610), .A2(new_n737), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n335), .A2(new_n603), .A3(new_n662), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G134), .ZN(G36));
  AOI21_X1  g567(.A(new_n665), .B1(new_n608), .B2(new_n614), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(KEYINPUT113), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n513), .B1(new_n627), .B2(new_n626), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(KEYINPUT43), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(KEYINPUT112), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT43), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n512), .B(new_n494), .C1(new_n628), .C2(KEYINPUT111), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n628), .A2(KEYINPUT111), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n755), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n392), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT45), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n398), .B1(new_n768), .B2(new_n336), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(KEYINPUT109), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n395), .A2(new_n397), .A3(KEYINPUT45), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT110), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n393), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n767), .B1(new_n774), .B2(KEYINPUT46), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT46), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n776), .B1(new_n773), .B2(new_n393), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n403), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n666), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n755), .A2(KEYINPUT44), .A3(new_n763), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n766), .A2(new_n780), .A3(new_n729), .A4(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G137), .ZN(G39));
  INV_X1    g597(.A(KEYINPUT47), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n779), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n402), .B1(new_n775), .B2(new_n777), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT47), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n603), .A2(new_n737), .A3(new_n722), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(new_n728), .A3(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G140), .ZN(G42));
  INV_X1    g605(.A(new_n677), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n792), .A2(new_n673), .A3(new_n406), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n602), .A2(new_n402), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n715), .A2(new_n716), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT49), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n793), .A2(new_n756), .A3(new_n794), .A4(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n552), .B1(new_n758), .B2(new_n762), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n798), .A2(new_n714), .A3(new_n729), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT118), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n785), .A2(new_n787), .A3(KEYINPUT119), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n795), .A2(new_n402), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT119), .B1(new_n785), .B2(new_n787), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n800), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n717), .A2(new_n729), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n603), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n674), .A2(new_n553), .ZN(new_n808));
  NOR4_X1   g622(.A1(new_n807), .A2(new_n808), .A3(new_n513), .A4(new_n628), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n798), .A2(new_n806), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n810), .A2(new_n665), .A3(new_n713), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n792), .A2(new_n405), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n798), .A2(new_n717), .A3(new_n714), .A4(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT50), .ZN(new_n814));
  OR2_X1    g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n813), .A2(new_n814), .ZN(new_n816));
  AOI211_X1 g630(.A(new_n809), .B(new_n811), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT51), .B1(new_n805), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n785), .A2(new_n787), .A3(new_n802), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n800), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n817), .A2(new_n820), .A3(KEYINPUT51), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n550), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n638), .A2(new_n494), .A3(new_n548), .A4(new_n660), .ZN(new_n824));
  OR2_X1    g638(.A1(new_n824), .A2(KEYINPUT114), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(KEYINPUT114), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n335), .A2(new_n825), .A3(new_n651), .A4(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n723), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n751), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n629), .B1(new_n513), .B2(new_n548), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n831), .A2(new_n718), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n608), .A2(new_n611), .A3(new_n832), .A4(new_n614), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n652), .A2(new_n833), .A3(new_n604), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n704), .A2(new_n709), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n707), .A2(new_n720), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n830), .A2(new_n834), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n747), .B1(new_n745), .B2(new_n746), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n752), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT115), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n661), .A2(KEYINPUT116), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n661), .A2(KEYINPUT116), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n610), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n673), .A2(new_n844), .A3(new_n665), .A4(new_n719), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n663), .A2(new_n688), .A3(new_n845), .A4(new_n724), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n704), .A2(new_n707), .A3(new_n709), .A4(new_n720), .ZN(new_n849));
  INV_X1    g663(.A(new_n751), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n850), .B1(new_n827), .B2(new_n828), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n652), .A2(new_n833), .A3(new_n604), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n849), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n752), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(new_n740), .B2(new_n748), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n853), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n841), .A2(new_n848), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n858), .B(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT54), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n798), .A2(new_n703), .A3(new_n714), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n752), .A2(KEYINPUT53), .ZN(new_n863));
  NOR4_X1   g677(.A1(new_n849), .A2(new_n851), .A3(new_n852), .A4(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT117), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n731), .A2(new_n739), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n848), .A2(new_n864), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n663), .A2(new_n724), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n868), .A2(new_n847), .A3(new_n688), .A4(new_n845), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n846), .A2(KEYINPUT52), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n869), .A2(new_n866), .A3(new_n870), .ZN(new_n871));
  AND4_X1   g685(.A1(new_n704), .A2(new_n707), .A3(new_n709), .A4(new_n720), .ZN(new_n872));
  INV_X1    g686(.A(new_n863), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n872), .A2(new_n830), .A3(new_n834), .A4(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT117), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  AOI22_X1  g689(.A1(new_n858), .A2(new_n859), .B1(new_n867), .B2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n823), .A2(new_n861), .A3(new_n862), .A4(new_n878), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n807), .A2(new_n808), .A3(new_n629), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n798), .A2(new_n736), .A3(new_n806), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT48), .Z(new_n882));
  NOR3_X1   g696(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(G952), .A2(G953), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n797), .B1(new_n883), .B2(new_n884), .ZN(G75));
  NAND2_X1  g699(.A1(new_n419), .A2(new_n427), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(new_n425), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT55), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT56), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n858), .A2(new_n859), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n867), .A2(new_n875), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(G902), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT120), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n876), .A2(new_n329), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT120), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n890), .B1(new_n899), .B2(new_n445), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n337), .A2(G952), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT56), .B1(new_n896), .B2(G210), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n902), .B1(new_n903), .B2(new_n888), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n900), .A2(new_n904), .ZN(G51));
  XNOR2_X1  g719(.A(new_n393), .B(KEYINPUT57), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n893), .A2(KEYINPUT54), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n907), .B1(new_n908), .B2(new_n878), .ZN(new_n909));
  INV_X1    g723(.A(new_n698), .ZN(new_n910));
  OAI21_X1  g724(.A(KEYINPUT121), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n894), .A2(KEYINPUT120), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n896), .A2(new_n897), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n773), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n891), .A2(new_n877), .A3(new_n892), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n877), .B1(new_n891), .B2(new_n892), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n906), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT121), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n917), .A2(new_n918), .A3(new_n698), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n911), .A2(new_n914), .A3(new_n919), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n920), .A2(new_n902), .ZN(G54));
  NAND2_X1  g735(.A1(KEYINPUT58), .A2(G475), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT122), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n506), .B1(new_n899), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n506), .ZN(new_n926));
  AOI211_X1 g740(.A(new_n926), .B(new_n923), .C1(new_n895), .C2(new_n898), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n925), .A2(new_n927), .A3(new_n901), .ZN(G60));
  AND2_X1   g742(.A1(new_n622), .A2(new_n625), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n929), .B1(new_n915), .B2(new_n916), .ZN(new_n930));
  NAND2_X1  g744(.A1(G478), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT59), .Z(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n861), .B2(new_n878), .ZN(new_n933));
  OAI221_X1 g747(.A(new_n902), .B1(new_n930), .B2(new_n932), .C1(new_n933), .C2(new_n929), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(G63));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n936));
  NAND2_X1  g750(.A1(G217), .A2(G902), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT60), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n893), .A2(new_n936), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(KEYINPUT123), .B1(new_n876), .B2(new_n938), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n645), .ZN(new_n943));
  INV_X1    g757(.A(new_n587), .ZN(new_n944));
  INV_X1    g758(.A(new_n586), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n940), .B(new_n941), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n943), .A2(new_n902), .A3(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n943), .A2(KEYINPUT61), .A3(new_n946), .A4(new_n902), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(G66));
  NAND2_X1  g765(.A1(new_n872), .A2(new_n834), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n337), .ZN(new_n953));
  OAI21_X1  g767(.A(G953), .B1(new_n556), .B2(new_n423), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n886), .B1(G898), .B2(new_n337), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(G69));
  AND2_X1   g771(.A1(new_n868), .A2(new_n688), .ZN(new_n958));
  XNOR2_X1  g772(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n682), .A2(new_n684), .A3(new_n958), .A4(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n335), .A2(new_n603), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n962), .A2(new_n667), .A3(new_n751), .A4(new_n831), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n790), .A2(new_n960), .A3(new_n782), .A4(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n965), .B1(new_n685), .B2(new_n958), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n337), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n284), .A2(new_n286), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n501), .B1(new_n453), .B2(new_n500), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT124), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n968), .B(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n967), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n337), .A2(G900), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n766), .A2(new_n729), .A3(new_n781), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n736), .A2(new_n719), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n780), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n977), .A2(new_n790), .A3(new_n958), .A4(new_n855), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n973), .B1(new_n978), .B2(new_n337), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n972), .B1(new_n979), .B2(new_n971), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n337), .B1(G227), .B2(G900), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT126), .Z(new_n982));
  XNOR2_X1  g796(.A(new_n980), .B(new_n982), .ZN(G72));
  NAND2_X1  g797(.A1(G472), .A2(G902), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT63), .Z(new_n985));
  NAND2_X1  g799(.A1(new_n290), .A2(new_n327), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n860), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n985), .B1(new_n978), .B2(new_n952), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n326), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n964), .A2(new_n966), .A3(new_n952), .ZN(new_n990));
  INV_X1    g804(.A(new_n985), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n325), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  AOI211_X1 g807(.A(new_n901), .B(new_n987), .C1(new_n993), .C2(new_n327), .ZN(G57));
endmodule


