//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 0 1 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 1 1 1 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n782, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978, new_n979;
  NOR3_X1   g000(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT90), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n202), .A2(KEYINPUT90), .ZN(new_n207));
  AOI22_X1  g006(.A1(new_n206), .A2(new_n207), .B1(G29gat), .B2(G36gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(G43gat), .B(G50gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT15), .ZN(new_n210));
  AOI22_X1  g009(.A1(new_n209), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(KEYINPUT15), .B2(new_n209), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n202), .A2(KEYINPUT91), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n202), .A2(KEYINPUT91), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n205), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI22_X1  g014(.A1(new_n208), .A2(new_n210), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT92), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT17), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n217), .B(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G15gat), .B(G22gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n220), .B(KEYINPUT93), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G1gat), .ZN(new_n222));
  INV_X1    g021(.A(G8gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT94), .ZN(new_n224));
  INV_X1    g023(.A(G1gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT16), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n222), .B(new_n224), .C1(new_n221), .C2(new_n226), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n223), .A2(KEYINPUT94), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n227), .B(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n219), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G229gat), .A2(G233gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n229), .A2(new_n216), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT18), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n231), .A2(KEYINPUT18), .A3(new_n232), .A4(new_n233), .ZN(new_n237));
  XOR2_X1   g036(.A(new_n232), .B(KEYINPUT13), .Z(new_n238));
  INV_X1    g037(.A(new_n233), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n229), .A2(new_n216), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n236), .A2(new_n237), .A3(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G113gat), .B(G141gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n243), .B(G197gat), .ZN(new_n244));
  XOR2_X1   g043(.A(KEYINPUT11), .B(G169gat), .Z(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n246), .B(KEYINPUT12), .Z(new_n247));
  NAND2_X1  g046(.A1(new_n242), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n247), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n236), .A2(new_n249), .A3(new_n237), .A4(new_n241), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(G1gat), .B(G29gat), .Z(new_n253));
  XNOR2_X1  g052(.A(G57gat), .B(G85gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT84), .B(KEYINPUT0), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n255), .B(new_n256), .Z(new_n257));
  INV_X1    g056(.A(KEYINPUT5), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT83), .ZN(new_n259));
  INV_X1    g058(.A(G113gat), .ZN(new_n260));
  INV_X1    g059(.A(G120gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(G113gat), .A2(G120gat), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XOR2_X1   g063(.A(KEYINPUT72), .B(KEYINPUT1), .Z(new_n265));
  XNOR2_X1  g064(.A(G127gat), .B(G134gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G134gat), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n268), .A2(KEYINPUT70), .A3(G127gat), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT70), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n269), .B1(new_n266), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT1), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n262), .A2(new_n272), .A3(new_n263), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT71), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n268), .A2(G127gat), .ZN(new_n275));
  INV_X1    g074(.A(G127gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G134gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n275), .A2(new_n277), .A3(new_n270), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n268), .A2(KEYINPUT70), .A3(G127gat), .ZN(new_n279));
  AND4_X1   g078(.A1(KEYINPUT71), .A2(new_n278), .A3(new_n273), .A4(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n267), .B1(new_n274), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT82), .ZN(new_n282));
  INV_X1    g081(.A(G141gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(G148gat), .ZN(new_n284));
  INV_X1    g083(.A(G148gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(G141gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(G155gat), .A2(G162gat), .ZN(new_n287));
  AOI22_X1  g086(.A1(new_n284), .A2(new_n286), .B1(KEYINPUT2), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G155gat), .ZN(new_n289));
  INV_X1    g088(.A(G162gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(KEYINPUT81), .A3(new_n287), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT81), .B1(new_n291), .B2(new_n287), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n282), .B(new_n288), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n287), .A2(KEYINPUT2), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n285), .A2(G141gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n283), .A2(G148gat), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n291), .A2(new_n287), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT81), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n299), .B1(new_n302), .B2(new_n292), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT82), .B1(new_n288), .B2(new_n300), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n295), .B(KEYINPUT3), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n281), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n288), .B1(new_n293), .B2(new_n294), .ZN(new_n307));
  INV_X1    g106(.A(new_n300), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n282), .B1(new_n299), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT3), .B1(new_n310), .B2(new_n295), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n259), .B1(new_n306), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n295), .B1(new_n303), .B2(new_n304), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT3), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n315), .A2(KEYINPUT83), .A3(new_n281), .A4(new_n305), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G225gat), .A2(G233gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n313), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT4), .B1(new_n319), .B2(new_n281), .ZN(new_n320));
  INV_X1    g119(.A(new_n267), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n271), .A2(KEYINPUT71), .A3(new_n273), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n278), .A2(new_n273), .A3(new_n279), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT71), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n321), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT4), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n326), .A2(new_n313), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n320), .A2(new_n328), .ZN(new_n329));
  AND4_X1   g128(.A1(new_n258), .A2(new_n317), .A3(new_n318), .A4(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n318), .ZN(new_n331));
  AND2_X1   g130(.A1(new_n326), .A2(new_n313), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n326), .A2(new_n313), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT5), .ZN(new_n335));
  AOI22_X1  g134(.A1(new_n312), .A2(new_n316), .B1(new_n320), .B2(new_n328), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n335), .B1(new_n336), .B2(new_n318), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n257), .B1(new_n330), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n317), .A2(new_n329), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT39), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n339), .A2(new_n340), .A3(new_n331), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n332), .A2(new_n333), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n340), .B1(new_n342), .B2(new_n318), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n343), .B1(new_n336), .B2(new_n318), .ZN(new_n344));
  INV_X1    g143(.A(new_n257), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n341), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT40), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n338), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n347), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT87), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n346), .A2(KEYINPUT87), .A3(new_n347), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n348), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AND2_X1   g152(.A1(G211gat), .A2(G218gat), .ZN(new_n354));
  OR2_X1    g153(.A1(new_n354), .A2(KEYINPUT22), .ZN(new_n355));
  XNOR2_X1  g154(.A(G197gat), .B(G204gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(G211gat), .A2(G218gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n355), .B(new_n356), .C1(new_n354), .C2(new_n358), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(G226gat), .A2(G233gat), .ZN(new_n363));
  INV_X1    g162(.A(G183gat), .ZN(new_n364));
  INV_X1    g163(.A(G190gat), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(new_n365), .A3(KEYINPUT64), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT64), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n367), .B1(G183gat), .B2(G190gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G183gat), .A2(G190gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT24), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT24), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n372), .A2(G183gat), .A3(G190gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(G169gat), .ZN(new_n376));
  INV_X1    g175(.A(G176gat), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT23), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT65), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT65), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n380), .A2(new_n376), .A3(new_n377), .A4(KEYINPUT23), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(G169gat), .A2(G176gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT23), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n376), .A2(new_n377), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n375), .A2(new_n382), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT25), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n388), .B1(new_n384), .B2(new_n385), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT66), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n391), .A2(new_n376), .A3(new_n377), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(KEYINPUT23), .A3(new_n393), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT68), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n364), .A2(KEYINPUT24), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n397), .A2(G190gat), .B1(KEYINPUT24), .B2(new_n370), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT67), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n399), .A2(new_n364), .A3(new_n365), .ZN(new_n400));
  OAI21_X1  g199(.A(KEYINPUT67), .B1(G183gat), .B2(G190gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n396), .B1(new_n398), .B2(new_n402), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n374), .A2(KEYINPUT68), .A3(new_n401), .A4(new_n400), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n395), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT28), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n364), .A2(KEYINPUT27), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT69), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n365), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT27), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(G183gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n364), .A2(KEYINPUT27), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT69), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n406), .B1(new_n409), .B2(new_n413), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n411), .A2(new_n412), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n415), .A2(KEYINPUT28), .A3(new_n365), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n383), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n418), .B1(KEYINPUT26), .B2(new_n385), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT26), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n392), .A2(new_n420), .A3(new_n393), .ZN(new_n421));
  AOI22_X1  g220(.A1(new_n419), .A2(new_n421), .B1(G183gat), .B2(G190gat), .ZN(new_n422));
  AOI22_X1  g221(.A1(new_n389), .A2(new_n405), .B1(new_n417), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n363), .B1(new_n423), .B2(KEYINPUT29), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n389), .A2(new_n405), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n417), .A2(new_n422), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n363), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT79), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT79), .ZN(new_n430));
  NOR3_X1   g229(.A1(new_n423), .A2(new_n430), .A3(new_n363), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n362), .B(new_n424), .C1(new_n429), .C2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT77), .B1(new_n423), .B2(new_n363), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT77), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n390), .A2(new_n394), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n374), .A2(new_n401), .A3(new_n400), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n435), .B1(new_n396), .B2(new_n436), .ZN(new_n437));
  AOI22_X1  g236(.A1(new_n437), .A2(new_n404), .B1(new_n388), .B2(new_n387), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n417), .A2(new_n422), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n434), .B(new_n428), .C1(new_n438), .C2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT29), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n441), .B1(new_n438), .B2(new_n439), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n433), .A2(new_n440), .B1(new_n442), .B2(new_n363), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n432), .B(KEYINPUT78), .C1(new_n362), .C2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n434), .B1(new_n427), .B2(new_n428), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n423), .A2(KEYINPUT77), .A3(new_n363), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n424), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT78), .ZN(new_n448));
  INV_X1    g247(.A(new_n362), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n444), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(G8gat), .B(G36gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(G64gat), .B(G92gat), .ZN(new_n453));
  XOR2_X1   g252(.A(new_n452), .B(new_n453), .Z(new_n454));
  AOI21_X1  g253(.A(KEYINPUT80), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT80), .ZN(new_n456));
  INV_X1    g255(.A(new_n454), .ZN(new_n457));
  AOI211_X1 g256(.A(new_n456), .B(new_n457), .C1(new_n444), .C2(new_n450), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n455), .A2(new_n458), .A3(KEYINPUT30), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n451), .A2(KEYINPUT30), .A3(new_n454), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT78), .B1(new_n443), .B2(new_n362), .ZN(new_n461));
  INV_X1    g260(.A(new_n432), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n450), .B(new_n457), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n353), .B1(new_n459), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(KEYINPUT31), .B(G50gat), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n362), .B1(new_n315), .B2(new_n441), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n362), .A2(new_n441), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n313), .B1(new_n468), .B2(new_n314), .ZN(new_n469));
  OAI211_X1 g268(.A(G228gat), .B(G233gat), .C1(new_n467), .C2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(G228gat), .A2(G233gat), .ZN(new_n472));
  INV_X1    g271(.A(new_n361), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT85), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT29), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n360), .A2(new_n361), .A3(KEYINPUT85), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT3), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n472), .B1(new_n477), .B2(new_n313), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n478), .A2(new_n467), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n466), .B1(new_n471), .B2(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(G78gat), .B(G106gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n481), .B(G22gat), .ZN(new_n482));
  INV_X1    g281(.A(new_n466), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n470), .B(new_n483), .C1(new_n467), .C2(new_n478), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n482), .B1(new_n480), .B2(new_n484), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n457), .A2(KEYINPUT37), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n463), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n444), .A2(KEYINPUT37), .A3(new_n450), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT38), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT6), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n336), .A2(new_n258), .A3(new_n318), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n317), .A2(new_n318), .A3(new_n329), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n494), .B(new_n345), .C1(new_n495), .C2(new_n335), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n338), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  OAI211_X1 g296(.A(KEYINPUT6), .B(new_n257), .C1(new_n330), .C2(new_n337), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n455), .A2(new_n458), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n449), .B(new_n424), .C1(new_n429), .C2(new_n431), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n501), .B(KEYINPUT37), .C1(new_n449), .C2(new_n443), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT38), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n489), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n492), .A2(new_n499), .A3(new_n500), .A4(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n465), .A2(new_n487), .A3(new_n505), .ZN(new_n506));
  NOR3_X1   g305(.A1(new_n443), .A2(KEYINPUT78), .A3(new_n362), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n448), .B1(new_n447), .B2(new_n449), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n507), .B1(new_n432), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n456), .B1(new_n509), .B2(new_n457), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT30), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n451), .A2(KEYINPUT80), .A3(new_n454), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n460), .A2(new_n463), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n487), .A2(KEYINPUT86), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT86), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n518), .B1(new_n485), .B2(new_n486), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n326), .B1(new_n438), .B2(new_n439), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n423), .A2(new_n281), .ZN(new_n522));
  INV_X1    g321(.A(G227gat), .ZN(new_n523));
  INV_X1    g322(.A(G233gat), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n521), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT32), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT33), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(G15gat), .B(G43gat), .Z(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT73), .ZN(new_n531));
  XNOR2_X1  g330(.A(G71gat), .B(G99gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n527), .A2(new_n529), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(KEYINPUT74), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(KEYINPUT33), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n526), .A2(KEYINPUT32), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT75), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT75), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n526), .A2(new_n539), .A3(KEYINPUT32), .A4(new_n536), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n533), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n542), .B1(new_n526), .B2(KEYINPUT32), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT74), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n543), .A2(new_n544), .A3(new_n529), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n535), .A2(new_n541), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n521), .A2(new_n522), .ZN(new_n547));
  INV_X1    g346(.A(new_n525), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n549), .A2(KEYINPUT34), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(KEYINPUT34), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n546), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n552), .A2(new_n535), .A3(new_n541), .A4(new_n545), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT36), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n556), .A2(KEYINPUT76), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n556), .A2(KEYINPUT76), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n554), .B(new_n555), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n558), .ZN(new_n560));
  AND3_X1   g359(.A1(new_n543), .A2(new_n544), .A3(new_n529), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n544), .B1(new_n543), .B2(new_n529), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n552), .B1(new_n563), .B2(new_n541), .ZN(new_n564));
  INV_X1    g363(.A(new_n555), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n560), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n516), .A2(new_n520), .B1(new_n559), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n506), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n487), .A2(new_n554), .A3(new_n555), .ZN(new_n569));
  OAI21_X1  g368(.A(KEYINPUT88), .B1(new_n516), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n464), .B1(new_n498), .B2(new_n497), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT88), .ZN(new_n572));
  AND3_X1   g371(.A1(new_n487), .A2(new_n554), .A3(new_n555), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n571), .A2(new_n572), .A3(new_n573), .A4(new_n513), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n570), .A2(KEYINPUT35), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT35), .ZN(new_n576));
  OAI211_X1 g375(.A(KEYINPUT88), .B(new_n576), .C1(new_n516), .C2(new_n569), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n568), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT89), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n574), .A2(KEYINPUT35), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n572), .B1(new_n581), .B2(new_n573), .ZN(new_n582));
  AOI22_X1  g381(.A1(new_n580), .A2(new_n582), .B1(new_n506), .B2(new_n567), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT89), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n583), .A2(new_n584), .A3(new_n575), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n252), .B1(new_n579), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G99gat), .A2(G106gat), .ZN(new_n587));
  INV_X1    g386(.A(G85gat), .ZN(new_n588));
  INV_X1    g387(.A(G92gat), .ZN(new_n589));
  AOI22_X1  g388(.A1(KEYINPUT8), .A2(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT102), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT101), .B(KEYINPUT7), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n588), .A2(new_n589), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G99gat), .B(G106gat), .Z(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT103), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n595), .B(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n219), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n595), .B(new_n597), .Z(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(new_n216), .ZN(new_n601));
  AND2_X1   g400(.A1(G232gat), .A2(G233gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT41), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n599), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(G190gat), .B(G218gat), .Z(new_n605));
  OR2_X1    g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n602), .A2(KEYINPUT41), .ZN(new_n609));
  XNOR2_X1  g408(.A(G134gat), .B(G162gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n606), .A2(new_n611), .A3(new_n607), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G71gat), .A2(G78gat), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT9), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(G64gat), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n621), .A2(G57gat), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(G57gat), .ZN(new_n623));
  OR2_X1    g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G71gat), .B(G78gat), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n625), .A2(KEYINPUT96), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n625), .A2(KEYINPUT96), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n620), .B(new_n624), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n629));
  NOR2_X1   g428(.A1(G71gat), .A2(G78gat), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT95), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n630), .B1(new_n631), .B2(new_n618), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n629), .B(new_n632), .C1(new_n631), .C2(new_n618), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT21), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(G183gat), .B(G211gat), .Z(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g439(.A(G127gat), .B(G155gat), .Z(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT98), .ZN(new_n642));
  NAND2_X1  g441(.A1(G231gat), .A2(G233gat), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n643), .B(KEYINPUT97), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n642), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n640), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n640), .A2(new_n645), .ZN(new_n648));
  INV_X1    g447(.A(new_n634), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n229), .B1(KEYINPUT21), .B2(new_n649), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n647), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n650), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n638), .B(new_n639), .Z(new_n653));
  INV_X1    g452(.A(new_n645), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n652), .B1(new_n655), .B2(new_n646), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n617), .B1(new_n651), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n650), .B1(new_n647), .B2(new_n648), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n655), .A2(new_n652), .A3(new_n646), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(new_n616), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g459(.A(G120gat), .B(G148gat), .Z(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT106), .ZN(new_n662));
  XNOR2_X1  g461(.A(G176gat), .B(G204gat), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n662), .B(new_n663), .Z(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n600), .A2(new_n649), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT10), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n598), .A2(new_n634), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n600), .A2(KEYINPUT10), .A3(new_n649), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(G230gat), .A2(G233gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT104), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n666), .A2(new_n668), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n673), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n665), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n675), .A2(KEYINPUT105), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n671), .A2(new_n680), .A3(new_n674), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n664), .B1(new_n676), .B2(new_n673), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n678), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n615), .A2(new_n657), .A3(new_n660), .A4(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n586), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(new_n514), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT107), .B(G1gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1324gat));
  NOR2_X1   g489(.A1(new_n459), .A2(new_n464), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT16), .B(G8gat), .Z(new_n693));
  AND3_X1   g492(.A1(new_n586), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n223), .B1(new_n586), .B2(new_n692), .ZN(new_n695));
  OAI21_X1  g494(.A(KEYINPUT42), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n696), .B1(KEYINPUT42), .B2(new_n694), .ZN(G1325gat));
  NAND2_X1  g496(.A1(new_n566), .A2(new_n559), .ZN(new_n698));
  OAI21_X1  g497(.A(G15gat), .B1(new_n687), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n554), .A2(new_n555), .ZN(new_n700));
  OR2_X1    g499(.A1(new_n700), .A2(G15gat), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n699), .B1(new_n687), .B2(new_n701), .ZN(G1326gat));
  INV_X1    g501(.A(new_n520), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n687), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(KEYINPUT43), .B(G22gat), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n704), .B(new_n705), .Z(G1327gat));
  INV_X1    g505(.A(G29gat), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n615), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n584), .B1(new_n583), .B2(new_n575), .ZN(new_n710));
  AND4_X1   g509(.A1(new_n584), .A2(new_n568), .A3(new_n575), .A4(new_n577), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n615), .ZN(new_n713));
  AOI21_X1  g512(.A(KEYINPUT44), .B1(new_n578), .B2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n651), .A2(new_n656), .A3(new_n617), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n616), .B1(new_n658), .B2(new_n659), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n684), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n251), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n712), .A2(new_n499), .A3(new_n715), .A4(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n707), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n725), .B1(new_n724), .B2(new_n723), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT45), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n718), .A2(new_n615), .A3(new_n719), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n586), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n514), .A2(G29gat), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n727), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n729), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n733), .A2(KEYINPUT45), .A3(new_n730), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n726), .A2(new_n732), .A3(new_n734), .ZN(G1328gat));
  INV_X1    g534(.A(new_n691), .ZN(new_n736));
  INV_X1    g535(.A(G36gat), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OR3_X1    g537(.A1(new_n729), .A2(KEYINPUT46), .A3(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(KEYINPUT46), .B1(new_n729), .B2(new_n738), .ZN(new_n740));
  INV_X1    g539(.A(new_n709), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n741), .B1(new_n579), .B2(new_n585), .ZN(new_n742));
  NOR4_X1   g541(.A1(new_n742), .A2(new_n691), .A3(new_n714), .A4(new_n721), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n739), .B(new_n740), .C1(new_n737), .C2(new_n743), .ZN(G1329gat));
  NOR4_X1   g543(.A1(new_n742), .A2(new_n698), .A3(new_n714), .A4(new_n721), .ZN(new_n745));
  INV_X1    g544(.A(G43gat), .ZN(new_n746));
  INV_X1    g545(.A(new_n700), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n746), .ZN(new_n748));
  OAI22_X1  g547(.A1(new_n745), .A2(new_n746), .B1(new_n729), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT47), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OAI221_X1 g550(.A(KEYINPUT47), .B1(new_n729), .B2(new_n748), .C1(new_n745), .C2(new_n746), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(G1330gat));
  NOR2_X1   g552(.A1(new_n703), .A2(G50gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n733), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(G50gat), .ZN(new_n756));
  NOR4_X1   g555(.A1(new_n742), .A2(new_n487), .A3(new_n714), .A4(new_n721), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n755), .B(KEYINPUT48), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n742), .A2(new_n714), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n759), .A2(new_n520), .A3(new_n722), .ZN(new_n760));
  AOI22_X1  g559(.A1(new_n760), .A2(G50gat), .B1(new_n733), .B2(new_n754), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n758), .B1(new_n761), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g561(.A(new_n718), .ZN(new_n763));
  NOR4_X1   g562(.A1(new_n763), .A2(new_n713), .A3(new_n251), .A4(new_n684), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n578), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n765), .A2(new_n514), .ZN(new_n766));
  XOR2_X1   g565(.A(new_n766), .B(G57gat), .Z(G1332gat));
  OR2_X1    g566(.A1(new_n765), .A2(KEYINPUT109), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n765), .A2(KEYINPUT109), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n770), .A2(new_n691), .ZN(new_n771));
  XNOR2_X1  g570(.A(KEYINPUT49), .B(G64gat), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n771), .B2(new_n774), .ZN(G1333gat));
  XOR2_X1   g574(.A(new_n700), .B(KEYINPUT110), .Z(new_n776));
  NOR3_X1   g575(.A1(new_n765), .A2(G71gat), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n698), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n768), .A2(new_n778), .A3(new_n769), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n777), .B1(new_n779), .B2(G71gat), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g580(.A1(new_n770), .A2(new_n703), .ZN(new_n782));
  XOR2_X1   g581(.A(new_n782), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g582(.A1(new_n718), .A2(new_n251), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n719), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n742), .A2(new_n714), .A3(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(G85gat), .B1(new_n787), .B2(new_n514), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n615), .B1(new_n583), .B2(new_n575), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n789), .A2(KEYINPUT51), .A3(new_n784), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n578), .A2(new_n713), .A3(new_n784), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n684), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n794), .A2(new_n588), .A3(new_n499), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n788), .A2(new_n795), .ZN(G1336gat));
  NOR3_X1   g595(.A1(new_n691), .A2(G92gat), .A3(new_n684), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT51), .B1(new_n789), .B2(new_n784), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n791), .A2(new_n792), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT111), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n785), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n712), .A2(new_n736), .A3(new_n715), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(G92gat), .ZN(new_n805));
  OAI211_X1 g604(.A(KEYINPUT111), .B(new_n797), .C1(new_n798), .C2(new_n799), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n802), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT52), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n805), .A2(new_n809), .A3(new_n800), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(G1337gat));
  OAI21_X1  g610(.A(G99gat), .B1(new_n787), .B2(new_n698), .ZN(new_n812));
  INV_X1    g611(.A(G99gat), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n794), .A2(new_n813), .A3(new_n747), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(G1338gat));
  NOR2_X1   g614(.A1(new_n487), .A2(G106gat), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n794), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(G106gat), .ZN(new_n820));
  INV_X1    g619(.A(new_n487), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n820), .B1(new_n786), .B2(new_n821), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n712), .A2(new_n520), .A3(new_n715), .A4(new_n803), .ZN(new_n823));
  AOI22_X1  g622(.A1(G106gat), .A2(new_n823), .B1(new_n794), .B2(new_n816), .ZN(new_n824));
  OAI22_X1  g623(.A1(new_n819), .A2(new_n822), .B1(new_n824), .B2(new_n818), .ZN(G1339gat));
  NOR3_X1   g624(.A1(new_n239), .A2(new_n240), .A3(new_n238), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n232), .B1(new_n231), .B2(new_n233), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n246), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n250), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n682), .A2(new_n683), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n669), .A2(new_n670), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n831), .B1(new_n832), .B2(new_n673), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n833), .A2(new_n679), .A3(new_n681), .ZN(new_n834));
  INV_X1    g633(.A(new_n675), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n665), .B1(new_n835), .B2(new_n831), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n834), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n837), .B1(new_n834), .B2(new_n836), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n829), .B(new_n830), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n718), .B1(new_n840), .B2(new_n713), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n251), .B(new_n830), .C1(new_n838), .C2(new_n839), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n719), .A2(new_n829), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(new_n843), .A3(new_n615), .ZN(new_n844));
  AOI22_X1  g643(.A1(new_n841), .A2(new_n844), .B1(new_n252), .B2(new_n686), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n845), .A2(new_n514), .A3(new_n736), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n573), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(new_n260), .A3(new_n251), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n736), .A2(new_n514), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n747), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n841), .A2(new_n844), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n686), .A2(new_n252), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(KEYINPUT112), .A3(new_n703), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n857), .B1(new_n845), .B2(new_n520), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n852), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n251), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n850), .B1(new_n860), .B2(G113gat), .ZN(new_n861));
  AOI211_X1 g660(.A(KEYINPUT113), .B(new_n260), .C1(new_n859), .C2(new_n251), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n849), .B1(new_n861), .B2(new_n862), .ZN(G1340gat));
  AOI21_X1  g662(.A(G120gat), .B1(new_n848), .B2(new_n719), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n684), .A2(new_n261), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n864), .B1(new_n859), .B2(new_n865), .ZN(G1341gat));
  NAND3_X1  g665(.A1(new_n859), .A2(G127gat), .A3(new_n718), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT114), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OR3_X1    g668(.A1(new_n847), .A2(KEYINPUT115), .A3(new_n763), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT115), .B1(new_n847), .B2(new_n763), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(new_n276), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n867), .A2(new_n868), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n869), .A2(new_n872), .A3(new_n873), .ZN(G1342gat));
  NAND4_X1  g673(.A1(new_n846), .A2(new_n268), .A3(new_n573), .A4(new_n713), .ZN(new_n875));
  XOR2_X1   g674(.A(new_n875), .B(KEYINPUT56), .Z(new_n876));
  AOI21_X1  g675(.A(new_n268), .B1(new_n859), .B2(new_n713), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n876), .A2(KEYINPUT116), .A3(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT116), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n875), .B(KEYINPUT56), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n880), .B1(new_n881), .B2(new_n877), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n879), .A2(new_n882), .ZN(G1343gat));
  NAND2_X1  g682(.A1(new_n851), .A2(new_n698), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n845), .A2(new_n885), .A3(new_n703), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n884), .B1(new_n886), .B2(KEYINPUT117), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n855), .A2(KEYINPUT57), .A3(new_n520), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n885), .B1(new_n845), .B2(new_n487), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT117), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n887), .A2(new_n891), .A3(new_n251), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n778), .A2(new_n487), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n846), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n252), .A2(G141gat), .ZN(new_n896));
  AOI22_X1  g695(.A1(new_n892), .A2(G141gat), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  XOR2_X1   g696(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n898));
  XNOR2_X1  g697(.A(new_n897), .B(new_n898), .ZN(G1344gat));
  NAND3_X1  g698(.A1(new_n895), .A2(new_n285), .A3(new_n719), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n887), .A2(new_n891), .ZN(new_n901));
  AOI211_X1 g700(.A(KEYINPUT59), .B(new_n285), .C1(new_n901), .C2(new_n719), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n855), .A2(new_n885), .A3(new_n520), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT57), .B1(new_n845), .B2(new_n487), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n851), .A2(new_n698), .A3(new_n719), .ZN(new_n906));
  OAI21_X1  g705(.A(G148gat), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  XOR2_X1   g706(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n908));
  AND2_X1   g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n900), .B1(new_n902), .B2(new_n909), .ZN(G1345gat));
  NAND3_X1  g709(.A1(new_n895), .A2(new_n289), .A3(new_n718), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n901), .A2(new_n718), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n911), .B1(new_n912), .B2(new_n289), .ZN(G1346gat));
  AOI21_X1  g712(.A(G162gat), .B1(new_n895), .B2(new_n713), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n615), .A2(new_n290), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n914), .B1(new_n901), .B2(new_n915), .ZN(G1347gat));
  NOR2_X1   g715(.A1(new_n691), .A2(new_n499), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n845), .A2(new_n569), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(G169gat), .B1(new_n919), .B2(new_n251), .ZN(new_n920));
  AOI211_X1 g719(.A(new_n776), .B(new_n918), .C1(new_n856), .C2(new_n858), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n252), .A2(new_n376), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(G1348gat));
  NAND3_X1  g722(.A1(new_n921), .A2(G176gat), .A3(new_n719), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT120), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  AOI21_X1  g726(.A(G176gat), .B1(new_n919), .B2(new_n719), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(G1349gat));
  NAND3_X1  g728(.A1(new_n919), .A2(new_n415), .A3(new_n718), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(KEYINPUT121), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n918), .A2(new_n776), .ZN(new_n932));
  INV_X1    g731(.A(new_n856), .ZN(new_n933));
  INV_X1    g732(.A(new_n858), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n718), .B(new_n932), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n931), .B1(new_n935), .B2(G183gat), .ZN(new_n936));
  XNOR2_X1  g735(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n936), .B(new_n938), .ZN(G1350gat));
  NAND3_X1  g738(.A1(new_n919), .A2(new_n365), .A3(new_n713), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT61), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n921), .A2(new_n713), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n941), .B1(new_n942), .B2(G190gat), .ZN(new_n943));
  AOI211_X1 g742(.A(KEYINPUT61), .B(new_n365), .C1(new_n921), .C2(new_n713), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n940), .B1(new_n943), .B2(new_n944), .ZN(G1351gat));
  XNOR2_X1  g744(.A(KEYINPUT124), .B(G197gat), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n918), .A2(new_n778), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n903), .A2(new_n904), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n946), .B1(new_n948), .B2(new_n252), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n845), .A2(new_n918), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(new_n893), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(KEYINPUT123), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT123), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n252), .A2(new_n946), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT125), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AND4_X1   g757(.A1(KEYINPUT125), .A2(new_n953), .A3(new_n955), .A4(new_n957), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n949), .B1(new_n958), .B2(new_n959), .ZN(G1352gat));
  AOI21_X1  g759(.A(G204gat), .B1(KEYINPUT126), .B2(KEYINPUT62), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n952), .A2(new_n719), .A3(new_n961), .ZN(new_n962));
  NOR2_X1   g761(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n962), .B(new_n963), .ZN(new_n964));
  OAI21_X1  g763(.A(G204gat), .B1(new_n948), .B2(new_n684), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1353gat));
  NOR2_X1   g765(.A1(new_n763), .A2(G211gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n953), .A2(new_n955), .A3(new_n967), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n903), .A2(new_n904), .A3(new_n718), .A4(new_n947), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n969), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n970));
  AOI21_X1  g769(.A(KEYINPUT63), .B1(new_n969), .B2(G211gat), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n968), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT127), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI211_X1 g773(.A(new_n968), .B(KEYINPUT127), .C1(new_n970), .C2(new_n971), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(G1354gat));
  INV_X1    g775(.A(G218gat), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n956), .A2(new_n977), .A3(new_n713), .ZN(new_n978));
  OAI21_X1  g777(.A(G218gat), .B1(new_n948), .B2(new_n615), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(G1355gat));
endmodule


