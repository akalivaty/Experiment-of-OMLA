//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 1 1 0 1 0 1 0 0 0 1 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n602, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1130,
    new_n1131;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT66), .B(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT67), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT68), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n463), .B(KEYINPUT69), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G137), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  OR2_X1    g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n474), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(new_n462), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n471), .A2(new_n476), .ZN(G160));
  NOR2_X1   g052(.A1(new_n468), .A2(new_n462), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n482), .B1(G136), .B2(new_n469), .ZN(G162));
  INV_X1    g058(.A(G138), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(KEYINPUT72), .C1(new_n467), .C2(new_n466), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT71), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n462), .A2(G138), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n490), .B1(new_n472), .B2(new_n473), .ZN(new_n491));
  AOI21_X1  g066(.A(KEYINPUT71), .B1(new_n491), .B2(KEYINPUT72), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n485), .B(KEYINPUT71), .C1(new_n467), .C2(new_n466), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n489), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n500));
  AND2_X1   g075(.A1(G126), .A2(G2105), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(new_n474), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n500), .B(new_n501), .C1(new_n466), .C2(new_n467), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n499), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n495), .A2(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n512));
  XOR2_X1   g087(.A(KEYINPUT6), .B(G651), .Z(new_n513));
  OR2_X1    g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n511), .A2(G62), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT73), .ZN(new_n517));
  OAI21_X1  g092(.A(G651), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n519), .A2(KEYINPUT74), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(KEYINPUT74), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(G166));
  AND2_X1   g097(.A1(new_n509), .A2(new_n510), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n523), .A2(new_n513), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G89), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n525), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT75), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n513), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT6), .B(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT75), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n531), .A2(G543), .A3(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n529), .B1(G51), .B2(new_n535), .ZN(G168));
  NAND2_X1  g111(.A1(new_n524), .A2(G90), .ZN(new_n537));
  INV_X1    g112(.A(G651), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G52), .ZN(new_n540));
  OAI221_X1 g115(.A(new_n537), .B1(new_n538), .B2(new_n539), .C1(new_n534), .C2(new_n540), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT76), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND2_X1  g118(.A1(new_n535), .A2(G43), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n538), .ZN(new_n546));
  XNOR2_X1  g121(.A(KEYINPUT77), .B(G81), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n524), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n544), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  NAND2_X1  g130(.A1(new_n524), .A2(G91), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n511), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n531), .A2(G53), .A3(G543), .A4(new_n533), .ZN(new_n558));
  AND2_X1   g133(.A1(KEYINPUT78), .A2(KEYINPUT9), .ZN(new_n559));
  AND2_X1   g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n558), .A2(new_n559), .ZN(new_n561));
  OAI221_X1 g136(.A(new_n556), .B1(new_n538), .B2(new_n557), .C1(new_n560), .C2(new_n561), .ZN(G299));
  INV_X1    g137(.A(G168), .ZN(G286));
  INV_X1    g138(.A(G166), .ZN(G303));
  NAND2_X1  g139(.A1(new_n535), .A2(G49), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n524), .A2(G87), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(G288));
  INV_X1    g143(.A(G61), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(new_n509), .B2(new_n510), .ZN(new_n570));
  AND2_X1   g145(.A1(G73), .A2(G543), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n532), .A2(G48), .A3(G543), .ZN(new_n573));
  AND2_X1   g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n511), .A2(new_n532), .A3(G86), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(G305));
  AOI22_X1  g151(.A1(new_n535), .A2(G47), .B1(G85), .B2(new_n524), .ZN(new_n577));
  NAND2_X1  g152(.A1(G72), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G60), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n523), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT79), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n538), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n582), .B1(new_n581), .B2(new_n580), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n577), .A2(new_n583), .ZN(G290));
  INV_X1    g159(.A(G868), .ZN(new_n585));
  NOR2_X1   g160(.A1(G301), .A2(new_n585), .ZN(new_n586));
  AND3_X1   g161(.A1(new_n511), .A2(new_n532), .A3(G92), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT10), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n511), .A2(G66), .ZN(new_n589));
  NAND2_X1  g164(.A1(G79), .A2(G543), .ZN(new_n590));
  XOR2_X1   g165(.A(new_n590), .B(KEYINPUT80), .Z(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  AND2_X1   g167(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n535), .A2(G54), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT81), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n586), .B1(new_n596), .B2(new_n585), .ZN(G284));
  AOI21_X1  g172(.A(new_n586), .B1(new_n596), .B2(new_n585), .ZN(G321));
  NAND2_X1  g173(.A1(G299), .A2(new_n585), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(new_n585), .B2(G168), .ZN(G297));
  OAI21_X1  g175(.A(new_n599), .B1(new_n585), .B2(G168), .ZN(G280));
  INV_X1    g176(.A(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n596), .B1(new_n602), .B2(G860), .ZN(G148));
  NAND2_X1  g178(.A1(new_n596), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G868), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g182(.A1(new_n464), .A2(new_n474), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT12), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT13), .ZN(new_n610));
  INV_X1    g185(.A(G2100), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n469), .A2(G135), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n478), .A2(G123), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n462), .A2(G111), .ZN(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n614), .B(new_n615), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(G2096), .Z(new_n619));
  NAND3_X1  g194(.A1(new_n612), .A2(new_n613), .A3(new_n619), .ZN(G156));
  XNOR2_X1  g195(.A(KEYINPUT15), .B(G2435), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT82), .B(G2438), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(G2427), .B(G2430), .Z(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n625), .A2(KEYINPUT14), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2443), .B(G2446), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(G1341), .B(G1348), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G2451), .B(G2454), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT16), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT83), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n632), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(G14), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT84), .Z(G401));
  XNOR2_X1  g214(.A(G2072), .B(G2078), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT17), .Z(new_n641));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n642), .B2(new_n640), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT86), .Z(new_n649));
  NAND3_X1  g224(.A1(new_n645), .A2(new_n642), .A3(new_n640), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT85), .B(KEYINPUT18), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n646), .A2(new_n642), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n652), .B1(new_n641), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n649), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2096), .B(G2100), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(G227));
  XOR2_X1   g232(.A(G1971), .B(G1976), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT19), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1956), .B(G2474), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1961), .B(G1966), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g237(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  NOR3_X1   g238(.A1(new_n659), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n659), .A2(new_n662), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT20), .Z(new_n666));
  AOI211_X1 g241(.A(new_n664), .B(new_n666), .C1(new_n659), .C2(new_n663), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1991), .B(G1996), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1981), .B(G1986), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G229));
  NOR2_X1   g248(.A1(G16), .A2(G22), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(G166), .B2(G16), .ZN(new_n675));
  INV_X1    g250(.A(G1971), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(G16), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G23), .ZN(new_n679));
  INV_X1    g254(.A(G288), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n679), .B1(new_n680), .B2(new_n678), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT33), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT89), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(new_n683), .ZN(new_n684));
  MUX2_X1   g259(.A(G6), .B(G305), .S(G16), .Z(new_n685));
  XOR2_X1   g260(.A(KEYINPUT32), .B(G1981), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n677), .A2(new_n684), .A3(new_n687), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n688), .A2(KEYINPUT34), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(KEYINPUT34), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n478), .A2(G119), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT87), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  OAI21_X1  g268(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n694));
  INV_X1    g269(.A(G107), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n694), .B1(new_n695), .B2(G2105), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n469), .B2(G131), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  MUX2_X1   g273(.A(G25), .B(new_n698), .S(G29), .Z(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT88), .Z(new_n700));
  XOR2_X1   g275(.A(KEYINPUT35), .B(G1991), .Z(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n700), .A2(new_n702), .ZN(new_n704));
  MUX2_X1   g279(.A(G24), .B(G290), .S(G16), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G1986), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g282(.A1(new_n689), .A2(new_n690), .A3(new_n703), .A4(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n708), .B(new_n709), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n678), .A2(G19), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n550), .B2(new_n678), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT91), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G1341), .ZN(new_n714));
  INV_X1    g289(.A(G29), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G26), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT92), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT28), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n469), .A2(G140), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n478), .A2(G128), .ZN(new_n720));
  OR2_X1    g295(.A1(G104), .A2(G2105), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n721), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n718), .B1(new_n724), .B2(new_n715), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G2067), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n678), .A2(G4), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n596), .B2(new_n678), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n726), .B1(new_n728), .B2(G1348), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n714), .B(new_n729), .C1(G1348), .C2(new_n728), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT93), .ZN(new_n731));
  NOR2_X1   g306(.A1(G29), .A2(G35), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G162), .B2(G29), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT99), .B(KEYINPUT29), .Z(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G2090), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT100), .ZN(new_n738));
  INV_X1    g313(.A(G27), .ZN(new_n739));
  OR3_X1    g314(.A1(new_n739), .A2(KEYINPUT98), .A3(G29), .ZN(new_n740));
  OAI21_X1  g315(.A(KEYINPUT98), .B1(new_n739), .B2(G29), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n740), .B(new_n741), .C1(G164), .C2(new_n715), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G2078), .ZN(new_n743));
  NOR2_X1   g318(.A1(G168), .A2(new_n678), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n678), .B2(G21), .ZN(new_n745));
  INV_X1    g320(.A(G1966), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT31), .B(G11), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT96), .B(G28), .ZN(new_n749));
  AOI21_X1  g324(.A(G29), .B1(new_n749), .B2(KEYINPUT30), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(KEYINPUT30), .B2(new_n749), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n748), .B(new_n751), .C1(new_n618), .C2(new_n715), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT97), .Z(new_n753));
  INV_X1    g328(.A(new_n745), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n753), .B1(new_n754), .B2(G1966), .ZN(new_n755));
  NOR4_X1   g330(.A1(new_n738), .A2(new_n743), .A3(new_n747), .A4(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n735), .A2(new_n736), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT101), .Z(new_n758));
  NAND2_X1  g333(.A1(new_n678), .A2(G20), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT23), .Z(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G299), .B2(G16), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(G1956), .Z(new_n762));
  NOR2_X1   g337(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G5), .A2(G16), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G171), .B2(G16), .ZN(new_n765));
  INV_X1    g340(.A(G1961), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(G29), .A2(G32), .ZN(new_n768));
  AOI22_X1  g343(.A1(G105), .A2(new_n464), .B1(new_n469), .B2(G141), .ZN(new_n769));
  NAND3_X1  g344(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT26), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G129), .B2(new_n478), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT94), .Z(new_n774));
  AOI21_X1  g349(.A(new_n768), .B1(new_n774), .B2(G29), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT27), .B(G1996), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT95), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n775), .A2(new_n777), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n715), .A2(G33), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT25), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n474), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n783), .A2(new_n462), .ZN(new_n784));
  AOI211_X1 g359(.A(new_n782), .B(new_n784), .C1(G139), .C2(new_n469), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n780), .B1(new_n785), .B2(new_n715), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G2072), .ZN(new_n787));
  AND2_X1   g362(.A1(KEYINPUT24), .A2(G34), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n715), .B1(KEYINPUT24), .B2(G34), .ZN(new_n789));
  OAI22_X1  g364(.A1(G160), .A2(new_n715), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G2084), .ZN(new_n791));
  NOR4_X1   g366(.A1(new_n778), .A2(new_n779), .A3(new_n787), .A4(new_n791), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n756), .A2(new_n763), .A3(new_n767), .A4(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n731), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n710), .A2(new_n794), .ZN(G150));
  INV_X1    g370(.A(G150), .ZN(G311));
  NAND2_X1  g371(.A1(new_n524), .A2(G93), .ZN(new_n797));
  INV_X1    g372(.A(G55), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n534), .B2(new_n798), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT102), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(new_n538), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT103), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n550), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n804), .B2(new_n803), .ZN(new_n806));
  INV_X1    g381(.A(new_n803), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n807), .A2(KEYINPUT103), .A3(new_n550), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT38), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n596), .A2(G559), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT39), .ZN(new_n813));
  AOI21_X1  g388(.A(G860), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n813), .B2(new_n812), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n803), .A2(G860), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT37), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n817), .ZN(G145));
  XNOR2_X1  g393(.A(new_n698), .B(KEYINPUT105), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(new_n609), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n478), .A2(G130), .ZN(new_n821));
  OR2_X1    g396(.A1(G106), .A2(G2105), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n822), .B(G2104), .C1(G118), .C2(new_n462), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(G142), .B2(new_n469), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n820), .B(new_n825), .ZN(new_n826));
  MUX2_X1   g401(.A(new_n773), .B(new_n774), .S(new_n785), .Z(new_n827));
  NAND2_X1  g402(.A1(new_n505), .A2(KEYINPUT104), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n501), .B1(new_n466), .B2(new_n467), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(KEYINPUT70), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(new_n503), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT104), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n831), .A2(new_n832), .A3(new_n499), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n495), .B1(new_n828), .B2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n723), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n827), .B(new_n835), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n826), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(G160), .B(new_n618), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(G162), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n826), .A2(new_n836), .ZN(new_n841));
  AOI21_X1  g416(.A(G37), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT106), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n837), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n841), .ZN(new_n845));
  INV_X1    g420(.A(new_n839), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n842), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g423(.A(new_n604), .B(KEYINPUT107), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n809), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n593), .A2(new_n594), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(G299), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n852), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n854), .A2(KEYINPUT41), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(KEYINPUT41), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n850), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(G166), .B(G288), .ZN(new_n858));
  XOR2_X1   g433(.A(G290), .B(G305), .Z(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT108), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n860), .B1(new_n861), .B2(KEYINPUT42), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(KEYINPUT42), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n862), .B(new_n863), .Z(new_n864));
  AND3_X1   g439(.A1(new_n853), .A2(new_n857), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n864), .B1(new_n853), .B2(new_n857), .ZN(new_n866));
  OAI21_X1  g441(.A(G868), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(G868), .B2(new_n807), .ZN(G295));
  OAI21_X1  g443(.A(new_n867), .B1(G868), .B2(new_n807), .ZN(G331));
  INV_X1    g444(.A(KEYINPUT44), .ZN(new_n870));
  XNOR2_X1  g445(.A(G301), .B(G168), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n809), .B(new_n871), .Z(new_n872));
  NAND2_X1  g447(.A1(new_n855), .A2(new_n856), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n809), .B(new_n871), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n852), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n874), .A2(new_n860), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(G37), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n860), .B1(new_n874), .B2(new_n876), .ZN(new_n880));
  XNOR2_X1  g455(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  OR3_X1    g457(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT110), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n855), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n856), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n855), .A2(new_n884), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n872), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n860), .B1(new_n888), .B2(new_n876), .ZN(new_n889));
  OAI21_X1  g464(.A(KEYINPUT43), .B1(new_n879), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n870), .B1(new_n883), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n889), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n892), .A2(new_n878), .A3(new_n877), .A4(new_n881), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n882), .B1(new_n879), .B2(new_n880), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n893), .A2(new_n894), .A3(new_n870), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n891), .A2(new_n895), .ZN(G397));
  INV_X1    g471(.A(KEYINPUT45), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(new_n834), .B2(G1384), .ZN(new_n898));
  OR2_X1    g473(.A1(new_n475), .A2(new_n462), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n899), .A2(new_n465), .A3(G40), .A4(new_n470), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  OR3_X1    g477(.A1(new_n902), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n903));
  OAI21_X1  g478(.A(KEYINPUT46), .B1(new_n902), .B2(G1996), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n723), .B(G2067), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n905), .A2(new_n773), .ZN(new_n906));
  AOI22_X1  g481(.A1(new_n903), .A2(new_n904), .B1(new_n901), .B2(new_n906), .ZN(new_n907));
  XOR2_X1   g482(.A(new_n907), .B(KEYINPUT47), .Z(new_n908));
  INV_X1    g483(.A(G1996), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n909), .B1(new_n769), .B2(new_n772), .ZN(new_n910));
  AOI211_X1 g485(.A(new_n905), .B(new_n910), .C1(new_n774), .C2(new_n909), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n698), .A2(new_n702), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n723), .A2(G2067), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n902), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n698), .A2(new_n702), .ZN(new_n916));
  INV_X1    g491(.A(new_n912), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n911), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n918), .A2(new_n901), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT48), .ZN(new_n920));
  OR3_X1    g495(.A1(new_n902), .A2(G1986), .A3(G290), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n921), .A2(new_n920), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n915), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n908), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g500(.A(new_n925), .B(KEYINPUT127), .Z(new_n926));
  INV_X1    g501(.A(G8), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT50), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(new_n834), .B2(G1384), .ZN(new_n929));
  INV_X1    g504(.A(G1384), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n930), .B1(new_n495), .B2(new_n505), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n931), .A2(new_n928), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n900), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n736), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n832), .B1(new_n831), .B2(new_n499), .ZN(new_n935));
  AOI211_X1 g510(.A(KEYINPUT104), .B(new_n498), .C1(new_n830), .C2(new_n503), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI211_X1 g512(.A(KEYINPUT45), .B(new_n930), .C1(new_n937), .C2(new_n495), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n900), .B1(new_n931), .B2(new_n897), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n676), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n927), .B1(new_n934), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(G166), .A2(new_n927), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n943), .B(KEYINPUT55), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(G1981), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n572), .A2(new_n946), .A3(new_n575), .A4(new_n573), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT112), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n947), .B(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n524), .ZN(new_n950));
  XOR2_X1   g525(.A(KEYINPUT113), .B(G86), .Z(new_n951));
  OAI21_X1  g526(.A(new_n574), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(G1981), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n949), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT49), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n492), .A2(new_n494), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n957), .B(new_n489), .C1(new_n935), .C2(new_n936), .ZN(new_n958));
  INV_X1    g533(.A(G40), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n471), .A2(new_n959), .A3(new_n476), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n958), .A2(new_n930), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n949), .A2(new_n953), .A3(KEYINPUT49), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n956), .A2(G8), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n961), .A2(G8), .ZN(new_n964));
  INV_X1    g539(.A(G1976), .ZN(new_n965));
  NOR2_X1   g540(.A1(G288), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT52), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n680), .A2(G1976), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT52), .B1(G288), .B2(new_n965), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n968), .A2(new_n969), .A3(new_n961), .A4(G8), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n963), .A2(new_n967), .A3(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n949), .ZN(new_n972));
  NOR2_X1   g547(.A1(G288), .A2(G1976), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n972), .B1(new_n963), .B2(new_n973), .ZN(new_n974));
  OAI22_X1  g549(.A1(new_n945), .A2(new_n971), .B1(new_n964), .B2(new_n974), .ZN(new_n975));
  XOR2_X1   g550(.A(new_n943), .B(KEYINPUT55), .Z(new_n976));
  OAI211_X1 g551(.A(new_n928), .B(new_n930), .C1(new_n495), .C2(new_n505), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n960), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n834), .A2(G1384), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n979), .B1(new_n980), .B2(new_n928), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n982));
  AOI21_X1  g557(.A(G2090), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n979), .B(KEYINPUT114), .C1(new_n980), .C2(new_n928), .ZN(new_n984));
  AOI22_X1  g559(.A1(new_n983), .A2(new_n984), .B1(new_n676), .B2(new_n940), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n976), .B(KEYINPUT115), .C1(new_n985), .C2(new_n927), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT115), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n928), .B1(new_n958), .B2(new_n930), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n982), .B1(new_n988), .B2(new_n978), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n984), .A2(new_n989), .A3(new_n736), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n927), .B1(new_n990), .B2(new_n941), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n987), .B1(new_n991), .B2(new_n944), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n971), .B1(new_n942), .B2(new_n944), .ZN(new_n993));
  INV_X1    g568(.A(G2078), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n938), .A2(new_n939), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI211_X1 g572(.A(KEYINPUT45), .B(new_n930), .C1(new_n495), .C2(new_n505), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n960), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n1000), .A2(new_n898), .A3(KEYINPUT53), .A4(new_n994), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n997), .B(new_n1001), .C1(G1961), .C2(new_n933), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(G171), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n986), .A2(new_n992), .A3(new_n993), .A4(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1966), .B1(new_n1000), .B2(new_n898), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n900), .A2(G2084), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1007), .B1(new_n929), .B2(new_n932), .ZN(new_n1008));
  OAI21_X1  g583(.A(G286), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT45), .B1(new_n958), .B2(new_n930), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n746), .B1(new_n1010), .B2(new_n999), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n900), .A2(G2084), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT50), .B1(new_n958), .B2(new_n930), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n931), .A2(new_n928), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1011), .A2(new_n1015), .A3(G168), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1009), .A2(G8), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT51), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT122), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT51), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1016), .A2(new_n1020), .A3(G8), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n1018), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1019), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1005), .B1(new_n1024), .B2(KEYINPUT62), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT62), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1026), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n975), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n986), .A2(new_n992), .A3(new_n993), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n471), .A2(new_n959), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT123), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n462), .B1(new_n475), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1032), .B1(new_n1031), .B2(new_n475), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT124), .B1(new_n1010), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT124), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n898), .A2(new_n1036), .A3(new_n1030), .A4(new_n1033), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n994), .A2(KEYINPUT53), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1038), .B1(new_n980), .B2(KEYINPUT45), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1035), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n960), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n766), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1040), .A2(G301), .A3(new_n1042), .A4(new_n997), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT54), .B1(new_n1003), .B2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1040), .A2(new_n997), .A3(new_n1042), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT125), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1040), .A2(KEYINPUT125), .A3(new_n1042), .A4(new_n997), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1047), .A2(G171), .A3(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1002), .A2(G171), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1044), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1023), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1018), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1055));
  AND4_X1   g630(.A1(new_n1029), .A2(new_n1053), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT121), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT57), .ZN(new_n1058));
  XNOR2_X1  g633(.A(G299), .B(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT56), .B(G2072), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n938), .A2(new_n939), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n958), .A2(new_n930), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n978), .B1(new_n1062), .B2(KEYINPUT50), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1059), .B(new_n1061), .C1(G1956), .C2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n961), .A2(G2067), .ZN(new_n1066));
  INV_X1    g641(.A(G1348), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1066), .B1(new_n1041), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT117), .B1(new_n1068), .B2(new_n595), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n933), .A2(G1348), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1070), .B(new_n851), .C1(new_n1071), .C2(new_n1066), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1061), .B1(new_n1063), .B2(G1956), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1059), .B1(new_n1074), .B2(KEYINPUT118), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT118), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1076), .B(new_n1061), .C1(new_n1063), .C2(G1956), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT119), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1073), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1075), .A2(KEYINPUT119), .A3(new_n1077), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1065), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n595), .A2(KEYINPUT60), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1068), .A2(new_n1082), .ZN(new_n1083));
  XOR2_X1   g658(.A(KEYINPUT58), .B(G1341), .Z(new_n1084));
  NAND2_X1  g659(.A1(new_n961), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1085), .B1(new_n940), .B2(G1996), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n549), .A2(KEYINPUT120), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1086), .A2(KEYINPUT59), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT59), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1089));
  NOR3_X1   g664(.A1(new_n1083), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n1071), .A2(new_n851), .A3(new_n1066), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1068), .A2(new_n595), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT60), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(G299), .B(KEYINPUT57), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT61), .B1(new_n1074), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n1064), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT61), .ZN(new_n1097));
  OR3_X1    g672(.A1(new_n1074), .A2(new_n1094), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1090), .A2(new_n1093), .A3(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1057), .B1(new_n1081), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1104), .A2(new_n1080), .A3(new_n1069), .A4(new_n1072), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n1064), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1090), .A2(new_n1099), .A3(new_n1093), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(KEYINPUT121), .A3(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1056), .A2(new_n1101), .A3(new_n1108), .ZN(new_n1109));
  OAI211_X1 g684(.A(G8), .B(G168), .C1(new_n1006), .C2(new_n1008), .ZN(new_n1110));
  AOI211_X1 g685(.A(new_n1110), .B(new_n971), .C1(new_n944), .C2(new_n942), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1111), .A2(new_n986), .A3(new_n992), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(KEYINPUT116), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT63), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT116), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1111), .A2(new_n1115), .A3(new_n986), .A4(new_n992), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1113), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1111), .B(KEYINPUT63), .C1(new_n944), .C2(new_n942), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1028), .A2(new_n1109), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT126), .ZN(new_n1121));
  INV_X1    g696(.A(new_n919), .ZN(new_n1122));
  XOR2_X1   g697(.A(G290), .B(G1986), .Z(new_n1123));
  OAI21_X1  g698(.A(new_n1122), .B1(new_n902), .B2(new_n1123), .ZN(new_n1124));
  XOR2_X1   g699(.A(new_n1124), .B(KEYINPUT111), .Z(new_n1125));
  AND3_X1   g700(.A1(new_n1120), .A2(new_n1121), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1121), .B1(new_n1120), .B2(new_n1125), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n926), .B1(new_n1126), .B2(new_n1127), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g703(.A1(new_n893), .A2(new_n894), .ZN(new_n1130));
  NOR4_X1   g704(.A1(G229), .A2(G401), .A3(new_n460), .A4(G227), .ZN(new_n1131));
  NAND3_X1  g705(.A1(new_n1130), .A2(new_n847), .A3(new_n1131), .ZN(G225));
  INV_X1    g706(.A(G225), .ZN(G308));
endmodule


