//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 0 0 1 1 0 0 0 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 1 1 0 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n805, new_n806, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1012, new_n1013;
  INV_X1    g000(.A(KEYINPUT86), .ZN(new_n202));
  INV_X1    g001(.A(G120gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G113gat), .ZN(new_n204));
  INV_X1    g003(.A(G113gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G120gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT67), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT1), .ZN(new_n209));
  XNOR2_X1  g008(.A(G127gat), .B(G134gat), .ZN(new_n210));
  AND3_X1   g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G113gat), .B(G120gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n212), .A2(new_n207), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n212), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(new_n209), .ZN(new_n216));
  INV_X1    g015(.A(G127gat), .ZN(new_n217));
  AND3_X1   g016(.A1(new_n217), .A2(KEYINPUT66), .A3(G134gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n218), .B1(new_n210), .B2(new_n219), .ZN(new_n220));
  AOI22_X1  g019(.A1(new_n211), .A2(new_n214), .B1(new_n216), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G141gat), .B(G148gat), .ZN(new_n222));
  OR2_X1    g021(.A1(new_n222), .A2(KEYINPUT2), .ZN(new_n223));
  INV_X1    g022(.A(G162gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G155gat), .ZN(new_n225));
  INV_X1    g024(.A(G155gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G162gat), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n223), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT75), .ZN(new_n231));
  INV_X1    g030(.A(G148gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(G141gat), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT74), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n236), .B1(new_n232), .B2(G141gat), .ZN(new_n237));
  INV_X1    g036(.A(G141gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n238), .A2(KEYINPUT74), .A3(G148gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n235), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT2), .B1(new_n226), .B2(KEYINPUT76), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n241), .A2(new_n225), .A3(new_n227), .ZN(new_n242));
  AND3_X1   g041(.A1(new_n240), .A2(KEYINPUT77), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT77), .B1(new_n240), .B2(new_n242), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n221), .B(new_n230), .C1(new_n243), .C2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT80), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT77), .ZN(new_n247));
  AND2_X1   g046(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n248));
  NOR2_X1   g047(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n249));
  NOR3_X1   g048(.A1(new_n248), .A2(new_n249), .A3(new_n238), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n237), .A2(new_n239), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n228), .A2(new_n241), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n247), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n240), .A2(KEYINPUT77), .A3(new_n242), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n254), .A2(new_n255), .B1(new_n229), .B2(new_n223), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT80), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n256), .A2(new_n257), .A3(new_n221), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n246), .A2(new_n258), .A3(KEYINPUT4), .ZN(new_n259));
  INV_X1    g058(.A(new_n245), .ZN(new_n260));
  XOR2_X1   g059(.A(KEYINPUT79), .B(KEYINPUT4), .Z(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G225gat), .A2(G233gat), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n230), .B1(new_n243), .B2(new_n244), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT78), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT78), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n268), .B(new_n230), .C1(new_n243), .C2(new_n244), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(KEYINPUT3), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT3), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n221), .B1(new_n256), .B2(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n265), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n263), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n217), .A2(G134gat), .ZN(new_n277));
  INV_X1    g076(.A(G134gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(G127gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n279), .A3(new_n219), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n280), .B1(new_n219), .B2(new_n277), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n212), .A2(KEYINPUT1), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n283));
  OAI22_X1  g082(.A1(new_n281), .A2(new_n282), .B1(new_n283), .B2(new_n213), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n267), .A2(new_n269), .A3(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(new_n246), .A3(new_n258), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT81), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n286), .A2(new_n287), .A3(new_n265), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n287), .B1(new_n286), .B2(new_n265), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT4), .B1(new_n246), .B2(new_n258), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n260), .A2(new_n261), .ZN(new_n292));
  OR2_X1    g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n274), .B1(new_n293), .B2(new_n273), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n276), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G1gat), .B(G29gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n296), .B(KEYINPUT0), .ZN(new_n297));
  XNOR2_X1  g096(.A(G57gat), .B(G85gat), .ZN(new_n298));
  XOR2_X1   g097(.A(new_n297), .B(new_n298), .Z(new_n299));
  OAI21_X1  g098(.A(new_n202), .B1(new_n295), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT6), .B1(new_n295), .B2(new_n299), .ZN(new_n301));
  AND3_X1   g100(.A1(new_n267), .A2(new_n269), .A3(new_n284), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n246), .A2(new_n258), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n265), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT81), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n270), .A2(new_n272), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n306), .B(new_n264), .C1(new_n291), .C2(new_n292), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n286), .A2(new_n287), .A3(new_n265), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n305), .A2(KEYINPUT5), .A3(new_n307), .A4(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n299), .B1(new_n309), .B2(new_n275), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT86), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n300), .A2(new_n301), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n309), .A2(new_n275), .ZN(new_n313));
  INV_X1    g112(.A(new_n299), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n313), .A2(KEYINPUT6), .A3(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G8gat), .B(G36gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(G64gat), .B(G92gat), .ZN(new_n317));
  XOR2_X1   g116(.A(new_n316), .B(new_n317), .Z(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(G169gat), .A2(G176gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT23), .ZN(new_n321));
  NAND2_X1  g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT23), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n323), .B1(G169gat), .B2(G176gat), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n321), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(G183gat), .A2(G190gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(KEYINPUT64), .ZN(new_n327));
  NAND2_X1  g126(.A1(G183gat), .A2(G190gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT24), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT24), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n330), .A2(G183gat), .A3(G190gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n325), .B1(new_n327), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n326), .B1(new_n329), .B2(new_n331), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n321), .A2(KEYINPUT25), .A3(new_n324), .A4(new_n322), .ZN(new_n335));
  OAI22_X1  g134(.A1(new_n333), .A2(KEYINPUT25), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT26), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n337), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n338), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n320), .A2(new_n337), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT65), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n341), .B1(new_n342), .B2(new_n320), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n339), .A2(new_n340), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(G183gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT27), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT27), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(G183gat), .ZN(new_n348));
  INV_X1    g147(.A(G190gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n346), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  OR2_X1    g149(.A1(new_n350), .A2(KEYINPUT28), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n350), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n344), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT29), .B1(new_n336), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(G226gat), .A2(G233gat), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT72), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n326), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT64), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT64), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n326), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n359), .A2(new_n332), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n325), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT25), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n335), .B1(new_n332), .B2(new_n358), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n353), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT71), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n336), .A2(KEYINPUT71), .A3(new_n353), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n368), .A2(new_n356), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT29), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT72), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n372), .A2(new_n373), .A3(new_n355), .ZN(new_n374));
  XNOR2_X1  g173(.A(G197gat), .B(G204gat), .ZN(new_n375));
  INV_X1    g174(.A(G211gat), .ZN(new_n376));
  INV_X1    g175(.A(G218gat), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n375), .B1(KEYINPUT22), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G211gat), .B(G218gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n379), .B(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n357), .A2(new_n370), .A3(new_n374), .A4(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n336), .A2(new_n356), .A3(new_n353), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n355), .A2(new_n371), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n381), .B(new_n384), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n319), .B1(new_n388), .B2(KEYINPUT37), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n389), .B1(KEYINPUT37), .B2(new_n388), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT38), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n383), .A2(new_n387), .A3(new_n318), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT37), .B1(new_n394), .B2(new_n381), .ZN(new_n395));
  AND4_X1   g194(.A1(new_n381), .A2(new_n357), .A3(new_n370), .A4(new_n374), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n391), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n393), .B1(new_n389), .B2(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n392), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n312), .A2(new_n315), .A3(new_n399), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n271), .B(new_n230), .C1(new_n243), .C2(new_n244), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n371), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT82), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n401), .A2(KEYINPUT82), .A3(new_n371), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n404), .A2(new_n381), .A3(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n271), .B1(new_n381), .B2(KEYINPUT29), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n267), .A2(new_n269), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(G228gat), .ZN(new_n409));
  INV_X1    g208(.A(G233gat), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(KEYINPUT83), .B1(new_n406), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n412), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT83), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n404), .A2(new_n381), .A3(new_n405), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n381), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n407), .A2(new_n266), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n411), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  XOR2_X1   g221(.A(KEYINPUT84), .B(G22gat), .Z(new_n423));
  XNOR2_X1  g222(.A(G78gat), .B(G106gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT31), .B(G50gat), .ZN(new_n425));
  XOR2_X1   g224(.A(new_n424), .B(new_n425), .Z(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT85), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n418), .A2(new_n422), .A3(new_n423), .A4(new_n427), .ZN(new_n428));
  NOR3_X1   g227(.A1(new_n406), .A2(new_n412), .A3(KEYINPUT83), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n415), .B1(new_n414), .B2(new_n416), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n422), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(G22gat), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n426), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n422), .B(new_n423), .C1(new_n429), .C2(new_n430), .ZN(new_n435));
  INV_X1    g234(.A(new_n427), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n423), .B1(new_n418), .B2(new_n422), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n428), .B(new_n434), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT86), .B1(new_n313), .B2(new_n314), .ZN(new_n440));
  AOI211_X1 g239(.A(new_n202), .B(new_n299), .C1(new_n309), .C2(new_n275), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n285), .A2(new_n264), .A3(new_n246), .A4(new_n258), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n259), .A2(new_n262), .B1(new_n270), .B2(new_n272), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n443), .B(KEYINPUT39), .C1(new_n444), .C2(new_n264), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n263), .A2(new_n306), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT39), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(new_n447), .A3(new_n265), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n445), .A2(new_n448), .A3(new_n299), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT40), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n445), .A2(new_n448), .A3(KEYINPUT40), .A4(new_n299), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT30), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n393), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n388), .A2(new_n319), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n383), .A2(new_n387), .A3(KEYINPUT30), .A4(new_n318), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n451), .A2(new_n452), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n439), .B1(new_n442), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n400), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT68), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n284), .A2(new_n461), .ZN(new_n462));
  OAI221_X1 g261(.A(KEYINPUT68), .B1(new_n283), .B2(new_n213), .C1(new_n282), .C2(new_n281), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n366), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(G227gat), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n465), .A2(new_n410), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n336), .A2(new_n461), .A3(new_n284), .A4(new_n353), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT32), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT69), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n468), .A2(KEYINPUT69), .A3(KEYINPUT32), .ZN(new_n472));
  XNOR2_X1  g271(.A(G15gat), .B(G43gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(G71gat), .B(G99gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n473), .B(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT33), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n475), .B1(new_n468), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n471), .A2(new_n472), .A3(new_n477), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n468), .B(KEYINPUT32), .C1(new_n476), .C2(new_n475), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT34), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n464), .A2(new_n467), .ZN(new_n482));
  INV_X1    g281(.A(new_n466), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI211_X1 g283(.A(KEYINPUT34), .B(new_n466), .C1(new_n464), .C2(new_n467), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n480), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT70), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n478), .A2(new_n486), .A3(new_n479), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n486), .B1(new_n478), .B2(new_n479), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT70), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(KEYINPUT36), .A3(new_n493), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n478), .A2(new_n486), .A3(new_n479), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n495), .A2(new_n492), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT36), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n309), .A2(new_n299), .A3(new_n275), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT6), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n315), .B1(new_n502), .B2(new_n310), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n455), .A2(KEYINPUT73), .A3(new_n456), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n454), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT73), .B1(new_n455), .B2(new_n456), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n499), .B1(new_n508), .B2(new_n439), .ZN(new_n509));
  INV_X1    g308(.A(new_n423), .ZN(new_n510));
  AOI211_X1 g309(.A(new_n421), .B(new_n510), .C1(new_n413), .C2(new_n417), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n511), .A2(new_n427), .B1(new_n431), .B2(new_n433), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n431), .A2(new_n510), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n513), .A2(new_n435), .A3(new_n436), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n495), .A2(new_n492), .A3(KEYINPUT70), .ZN(new_n515));
  INV_X1    g314(.A(new_n493), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n512), .B(new_n514), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT35), .B1(new_n508), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT35), .ZN(new_n519));
  INV_X1    g318(.A(new_n457), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n496), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n439), .A2(new_n521), .ZN(new_n522));
  NOR3_X1   g321(.A1(new_n440), .A2(new_n441), .A3(new_n502), .ZN(new_n523));
  INV_X1    g322(.A(new_n315), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI22_X1  g324(.A1(new_n460), .A2(new_n509), .B1(new_n518), .B2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G113gat), .B(G141gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(KEYINPUT87), .B(G197gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(KEYINPUT11), .B(G169gat), .Z(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT12), .ZN(new_n532));
  XOR2_X1   g331(.A(G43gat), .B(G50gat), .Z(new_n533));
  XNOR2_X1  g332(.A(KEYINPUT89), .B(KEYINPUT15), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT90), .ZN(new_n536));
  NOR2_X1   g335(.A1(G29gat), .A2(G36gat), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT14), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT15), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n533), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n541), .B1(G29gat), .B2(G36gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n536), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT88), .ZN(new_n544));
  AOI22_X1  g343(.A1(new_n539), .A2(new_n544), .B1(G29gat), .B2(G36gat), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(new_n544), .B2(new_n539), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(new_n541), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT91), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n543), .A2(new_n547), .A3(KEYINPUT91), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G15gat), .B(G22gat), .ZN(new_n553));
  INV_X1    g352(.A(G1gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT16), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n556), .B1(G1gat), .B2(new_n553), .ZN(new_n557));
  OR2_X1    g356(.A1(new_n557), .A2(G8gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(G8gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT93), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT93), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n552), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G229gat), .A2(G233gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT92), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT17), .B1(new_n550), .B2(new_n551), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT17), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n561), .B1(new_n548), .B2(new_n571), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n566), .B(new_n569), .C1(new_n570), .C2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n560), .B(KEYINPUT93), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n575), .A2(new_n550), .A3(new_n551), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n566), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n568), .B(KEYINPUT13), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n574), .A2(KEYINPUT18), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT94), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n573), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n552), .A2(new_n571), .ZN(new_n582));
  INV_X1    g381(.A(new_n572), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n584), .A2(KEYINPUT94), .A3(new_n566), .A4(new_n569), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT18), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n581), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n532), .B1(new_n579), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n577), .A2(new_n578), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n589), .B(new_n532), .C1(new_n573), .C2(new_n586), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n581), .A2(new_n585), .A3(KEYINPUT95), .A4(new_n586), .ZN(new_n592));
  AND2_X1   g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT95), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n587), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n588), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(KEYINPUT96), .B1(new_n526), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n460), .A2(new_n509), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n518), .A2(new_n525), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT96), .ZN(new_n601));
  INV_X1    g400(.A(new_n588), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n595), .A2(new_n592), .A3(new_n591), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n600), .A2(new_n601), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(G57gat), .ZN(new_n606));
  INV_X1    g405(.A(G64gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G57gat), .A2(G64gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(G71gat), .A2(G78gat), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n608), .B(new_n609), .C1(new_n611), .C2(KEYINPUT9), .ZN(new_n612));
  NOR2_X1   g411(.A1(G71gat), .A2(G78gat), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n613), .B1(KEYINPUT97), .B2(new_n610), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n612), .B(new_n614), .C1(KEYINPUT97), .C2(new_n610), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT98), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n607), .B1(new_n616), .B2(new_n606), .ZN(new_n617));
  NAND3_X1  g416(.A1(KEYINPUT98), .A2(G57gat), .A3(G64gat), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n613), .A2(KEYINPUT9), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n617), .B(new_n618), .C1(new_n619), .C2(new_n611), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT21), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(G231gat), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n624), .A2(new_n410), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  OAI211_X1 g425(.A(new_n621), .B(new_n622), .C1(new_n624), .C2(new_n410), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(G127gat), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT99), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n615), .A2(KEYINPUT21), .A3(new_n620), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n575), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n562), .A2(new_n564), .A3(new_n631), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(KEYINPUT99), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n629), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n629), .A3(new_n632), .ZN(new_n637));
  XNOR2_X1  g436(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(new_n226), .ZN(new_n639));
  XNOR2_X1  g438(.A(G183gat), .B(G211gat), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n639), .B(new_n640), .Z(new_n641));
  NAND3_X1  g440(.A1(new_n636), .A2(new_n637), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n641), .ZN(new_n643));
  INV_X1    g442(.A(new_n637), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n643), .B1(new_n644), .B2(new_n635), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(G134gat), .B(G162gat), .Z(new_n647));
  AND2_X1   g446(.A1(G232gat), .A2(G233gat), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n648), .A2(KEYINPUT41), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n647), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT100), .ZN(new_n651));
  NAND2_X1  g450(.A1(G85gat), .A2(G92gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT7), .ZN(new_n653));
  NAND2_X1  g452(.A1(G99gat), .A2(G106gat), .ZN(new_n654));
  INV_X1    g453(.A(G85gat), .ZN(new_n655));
  INV_X1    g454(.A(G92gat), .ZN(new_n656));
  AOI22_X1  g455(.A1(KEYINPUT8), .A2(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(G99gat), .B(G106gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n548), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n660), .B1(new_n661), .B2(KEYINPUT17), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n582), .A2(new_n662), .ZN(new_n663));
  AOI22_X1  g462(.A1(new_n552), .A2(new_n660), .B1(KEYINPUT41), .B2(new_n648), .ZN(new_n664));
  XOR2_X1   g463(.A(G190gat), .B(G218gat), .Z(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n663), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n666), .B1(new_n663), .B2(new_n664), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n651), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n669), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n650), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n671), .A2(new_n673), .A3(new_n667), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n646), .B1(new_n670), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(G230gat), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(new_n410), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n660), .B(new_n621), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT10), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n660), .A2(KEYINPUT10), .A3(new_n615), .A4(new_n620), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n677), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  OR3_X1    g482(.A1(new_n678), .A2(new_n676), .A3(new_n410), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(G120gat), .B(G148gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(G176gat), .B(G204gat), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n686), .B(new_n687), .Z(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n683), .A2(new_n684), .A3(new_n688), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n675), .A2(KEYINPUT101), .A3(new_n693), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n642), .A2(new_n645), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n671), .A2(new_n673), .A3(new_n667), .ZN(new_n696));
  INV_X1    g495(.A(new_n651), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n697), .B1(new_n671), .B2(new_n667), .ZN(new_n698));
  OAI211_X1 g497(.A(new_n695), .B(new_n693), .C1(new_n696), .C2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT101), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI22_X1  g500(.A1(new_n597), .A2(new_n605), .B1(new_n694), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n503), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT102), .B(G1gat), .Z(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1324gat));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n707));
  XOR2_X1   g506(.A(KEYINPUT16), .B(G8gat), .Z(new_n708));
  NAND3_X1  g507(.A1(new_n702), .A2(new_n457), .A3(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT42), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n597), .A2(new_n605), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n701), .A2(new_n694), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(G8gat), .B1(new_n714), .B2(new_n520), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n715), .A2(new_n709), .ZN(new_n716));
  OAI211_X1 g515(.A(new_n707), .B(new_n711), .C1(new_n716), .C2(new_n710), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n710), .B1(new_n715), .B2(new_n709), .ZN(new_n718));
  INV_X1    g517(.A(new_n711), .ZN(new_n719));
  OAI21_X1  g518(.A(KEYINPUT103), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n717), .A2(new_n720), .ZN(G1325gat));
  INV_X1    g520(.A(new_n496), .ZN(new_n722));
  OR3_X1    g521(.A1(new_n714), .A2(G15gat), .A3(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n499), .ZN(new_n724));
  OAI21_X1  g523(.A(G15gat), .B1(new_n714), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n725), .ZN(G1326gat));
  NAND2_X1  g525(.A1(new_n702), .A2(new_n439), .ZN(new_n727));
  XNOR2_X1  g526(.A(KEYINPUT43), .B(G22gat), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1327gat));
  NOR2_X1   g528(.A1(new_n695), .A2(new_n692), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n696), .A2(new_n698), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n712), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(G29gat), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n733), .A2(new_n734), .A3(new_n703), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT45), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n604), .A2(new_n730), .ZN(new_n738));
  INV_X1    g537(.A(new_n731), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n739), .B1(new_n598), .B2(new_n599), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT104), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT104), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n743), .B(KEYINPUT44), .C1(new_n526), .C2(new_n739), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n600), .A2(KEYINPUT105), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT105), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n526), .A2(new_n747), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n749));
  NAND4_X1  g548(.A1(new_n746), .A2(new_n748), .A3(new_n731), .A4(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n738), .B1(new_n745), .B2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(G29gat), .B1(new_n752), .B2(new_n503), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n735), .A2(new_n736), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n737), .A2(new_n753), .A3(new_n754), .ZN(G1328gat));
  INV_X1    g554(.A(G36gat), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n733), .A2(new_n756), .A3(new_n457), .ZN(new_n757));
  OR2_X1    g556(.A1(new_n757), .A2(KEYINPUT46), .ZN(new_n758));
  OAI21_X1  g557(.A(G36gat), .B1(new_n752), .B2(new_n520), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(KEYINPUT46), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(G1329gat));
  INV_X1    g560(.A(KEYINPUT47), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n751), .A2(new_n499), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G43gat), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n722), .A2(G43gat), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n712), .A2(new_n732), .A3(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n762), .B1(new_n764), .B2(new_n767), .ZN(new_n768));
  AOI211_X1 g567(.A(KEYINPUT47), .B(new_n766), .C1(new_n763), .C2(G43gat), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n768), .A2(new_n769), .ZN(G1330gat));
  INV_X1    g569(.A(G50gat), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n771), .B1(new_n751), .B2(new_n439), .ZN(new_n772));
  INV_X1    g571(.A(new_n439), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n773), .A2(G50gat), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n733), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT107), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT48), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n772), .B2(new_n776), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(G1331gat));
  AND2_X1   g582(.A1(new_n746), .A2(new_n748), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n604), .A2(new_n646), .A3(new_n731), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n785), .A2(new_n692), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  OR3_X1    g586(.A1(new_n787), .A2(KEYINPUT109), .A3(new_n503), .ZN(new_n788));
  OAI21_X1  g587(.A(KEYINPUT109), .B1(new_n787), .B2(new_n503), .ZN(new_n789));
  XNOR2_X1  g588(.A(KEYINPUT108), .B(G57gat), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n790), .B1(new_n788), .B2(new_n789), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n791), .A2(new_n792), .ZN(G1332gat));
  NOR2_X1   g592(.A1(new_n787), .A2(new_n520), .ZN(new_n794));
  NOR2_X1   g593(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n795));
  AND2_X1   g594(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n797), .B1(new_n794), .B2(new_n795), .ZN(G1333gat));
  OAI21_X1  g597(.A(G71gat), .B1(new_n787), .B2(new_n724), .ZN(new_n799));
  INV_X1    g598(.A(G71gat), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n496), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n799), .B1(new_n787), .B2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n802), .B(new_n803), .ZN(G1334gat));
  NOR2_X1   g603(.A1(new_n787), .A2(new_n773), .ZN(new_n805));
  XOR2_X1   g604(.A(KEYINPUT110), .B(G78gat), .Z(new_n806));
  XNOR2_X1  g605(.A(new_n805), .B(new_n806), .ZN(G1335gat));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n604), .A2(new_n695), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n740), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT51), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n810), .A2(KEYINPUT51), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n808), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n813), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n815), .A2(KEYINPUT111), .A3(new_n811), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n703), .A2(new_n655), .A3(new_n692), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n814), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n809), .A2(new_n692), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n820), .B1(new_n745), .B2(new_n750), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n655), .B1(new_n821), .B2(new_n703), .ZN(new_n822));
  OAI21_X1  g621(.A(KEYINPUT112), .B1(new_n819), .B2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n822), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT112), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n814), .A2(new_n816), .A3(new_n818), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n823), .A2(new_n827), .ZN(G1336gat));
  NAND2_X1  g627(.A1(new_n821), .A2(new_n457), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(G92gat), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n812), .A2(new_n813), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n693), .A2(G92gat), .A3(new_n520), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT52), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n810), .B(new_n835), .ZN(new_n836));
  AOI22_X1  g635(.A1(new_n829), .A2(G92gat), .B1(new_n836), .B2(new_n832), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n834), .B1(new_n837), .B2(new_n838), .ZN(G1337gat));
  INV_X1    g638(.A(new_n821), .ZN(new_n840));
  OAI21_X1  g639(.A(G99gat), .B1(new_n840), .B2(new_n724), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n814), .A2(new_n816), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n722), .A2(new_n693), .A3(G99gat), .ZN(new_n843));
  XOR2_X1   g642(.A(new_n843), .B(KEYINPUT114), .Z(new_n844));
  OAI21_X1  g643(.A(new_n841), .B1(new_n842), .B2(new_n844), .ZN(G1338gat));
  NOR3_X1   g644(.A1(new_n773), .A2(G106gat), .A3(new_n693), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT53), .B1(new_n831), .B2(new_n846), .ZN(new_n847));
  AOI211_X1 g646(.A(new_n773), .B(new_n820), .C1(new_n745), .C2(new_n750), .ZN(new_n848));
  OAI21_X1  g647(.A(G106gat), .B1(new_n848), .B2(KEYINPUT116), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n821), .A2(KEYINPUT116), .A3(new_n439), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n847), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(G106gat), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  XOR2_X1   g652(.A(new_n846), .B(KEYINPUT115), .Z(new_n854));
  AND2_X1   g653(.A1(new_n836), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(KEYINPUT53), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n851), .A2(new_n856), .ZN(G1339gat));
  NOR2_X1   g656(.A1(new_n570), .A2(new_n572), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n575), .B1(new_n550), .B2(new_n551), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n568), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n862), .B1(new_n577), .B2(new_n578), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n860), .A2(new_n861), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n531), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n603), .A2(new_n865), .A3(new_n692), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n680), .A2(new_n681), .A3(new_n677), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n683), .A2(KEYINPUT54), .A3(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n688), .B1(new_n682), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n868), .A2(KEYINPUT55), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n691), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT55), .B1(new_n868), .B2(new_n870), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n866), .B(new_n739), .C1(new_n596), .C2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n603), .A2(new_n865), .A3(new_n874), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n695), .B1(new_n877), .B2(new_n731), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  AND4_X1   g678(.A1(new_n602), .A2(new_n675), .A3(new_n603), .A4(new_n693), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(KEYINPUT118), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT118), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n879), .A2(new_n881), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n439), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n457), .B1(new_n491), .B2(new_n493), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(new_n703), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT119), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n205), .A3(new_n604), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n886), .A2(new_n703), .A3(new_n520), .A4(new_n496), .ZN(new_n891));
  OAI21_X1  g690(.A(G113gat), .B1(new_n891), .B2(new_n596), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(G1340gat));
  NAND3_X1  g692(.A1(new_n889), .A2(new_n203), .A3(new_n692), .ZN(new_n894));
  OAI21_X1  g693(.A(G120gat), .B1(new_n891), .B2(new_n693), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1341gat));
  OAI21_X1  g695(.A(G127gat), .B1(new_n891), .B2(new_n646), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n695), .A2(new_n217), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n897), .B1(new_n888), .B2(new_n898), .ZN(G1342gat));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n885), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n703), .A3(new_n773), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT56), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n739), .A2(G134gat), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n902), .A2(new_n903), .A3(new_n887), .A4(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(G134gat), .B1(new_n891), .B2(new_n739), .ZN(new_n906));
  INV_X1    g705(.A(new_n904), .ZN(new_n907));
  OAI21_X1  g706(.A(KEYINPUT56), .B1(new_n888), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n905), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT120), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n905), .A2(new_n906), .A3(new_n908), .A4(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(G1343gat));
  NOR3_X1   g712(.A1(new_n499), .A2(new_n503), .A3(new_n457), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT121), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n884), .B1(new_n879), .B2(new_n881), .ZN(new_n916));
  AOI211_X1 g715(.A(KEYINPUT118), .B(new_n880), .C1(new_n876), .C2(new_n878), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n439), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  XOR2_X1   g717(.A(KEYINPUT122), .B(KEYINPUT57), .Z(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n882), .A2(KEYINPUT57), .A3(new_n439), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n915), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n238), .B1(new_n922), .B2(new_n604), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n900), .A2(new_n439), .A3(new_n914), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n924), .A2(G141gat), .A3(new_n596), .ZN(new_n925));
  OAI21_X1  g724(.A(KEYINPUT58), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(new_n925), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT58), .ZN(new_n928));
  AOI211_X1 g727(.A(new_n596), .B(new_n915), .C1(new_n920), .C2(new_n921), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n927), .B(new_n928), .C1(new_n929), .C2(new_n238), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n926), .A2(new_n930), .ZN(G1344gat));
  OAI21_X1  g730(.A(KEYINPUT59), .B1(new_n924), .B2(new_n693), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n932), .A2(new_n233), .A3(new_n234), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n920), .A2(new_n921), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT59), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n915), .A2(new_n693), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n919), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n439), .B(new_n938), .C1(new_n916), .C2(new_n917), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT57), .ZN(new_n940));
  AOI22_X1  g739(.A1(new_n876), .A2(new_n878), .B1(new_n713), .B2(new_n596), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n941), .B2(new_n773), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(KEYINPUT123), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT123), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n944), .B(new_n940), .C1(new_n941), .C2(new_n773), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n939), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n946), .A2(new_n936), .ZN(new_n947));
  NAND2_X1  g746(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n933), .B(new_n937), .C1(new_n947), .C2(new_n948), .ZN(G1345gat));
  INV_X1    g748(.A(new_n924), .ZN(new_n950));
  XNOR2_X1  g749(.A(KEYINPUT76), .B(G155gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n950), .A2(new_n695), .A3(new_n951), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n922), .A2(new_n695), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n952), .B1(new_n953), .B2(new_n951), .ZN(G1346gat));
  NAND3_X1  g753(.A1(new_n950), .A2(new_n224), .A3(new_n731), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n922), .A2(new_n731), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n955), .B1(new_n956), .B2(new_n224), .ZN(G1347gat));
  NOR2_X1   g756(.A1(new_n517), .A2(new_n520), .ZN(new_n958));
  XOR2_X1   g757(.A(new_n958), .B(KEYINPUT124), .Z(new_n959));
  OAI211_X1 g758(.A(new_n503), .B(new_n959), .C1(new_n916), .C2(new_n917), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(G169gat), .B1(new_n961), .B2(new_n604), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n703), .A2(new_n520), .A3(new_n722), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n886), .A2(new_n963), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n604), .A2(G169gat), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n962), .B1(new_n965), .B2(new_n966), .ZN(G1348gat));
  OAI21_X1  g766(.A(G176gat), .B1(new_n964), .B2(new_n693), .ZN(new_n968));
  OR2_X1    g767(.A1(new_n693), .A2(G176gat), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n968), .B1(new_n960), .B2(new_n969), .ZN(G1349gat));
  NAND3_X1  g769(.A1(new_n695), .A2(new_n346), .A3(new_n348), .ZN(new_n971));
  OR3_X1    g770(.A1(new_n960), .A2(KEYINPUT125), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g771(.A(KEYINPUT125), .B1(new_n960), .B2(new_n971), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g773(.A(G183gat), .B1(new_n964), .B2(new_n646), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(KEYINPUT60), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT60), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n974), .A2(new_n978), .A3(new_n975), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n977), .A2(new_n979), .ZN(G1350gat));
  NAND3_X1  g779(.A1(new_n961), .A2(new_n349), .A3(new_n731), .ZN(new_n981));
  NOR2_X1   g780(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n965), .A2(new_n731), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n349), .B1(KEYINPUT126), .B2(KEYINPUT61), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n982), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI211_X1 g784(.A(new_n982), .B(new_n984), .C1(new_n964), .C2(new_n739), .ZN(new_n986));
  INV_X1    g785(.A(new_n986), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n981), .B1(new_n985), .B2(new_n987), .ZN(G1351gat));
  NOR3_X1   g787(.A1(new_n703), .A2(new_n499), .A3(new_n520), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n946), .A2(new_n604), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(G197gat), .ZN(new_n991));
  NOR3_X1   g790(.A1(new_n499), .A2(new_n773), .A3(new_n520), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n900), .A2(new_n503), .A3(new_n992), .ZN(new_n993));
  OR3_X1    g792(.A1(new_n993), .A2(G197gat), .A3(new_n596), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n995), .A2(KEYINPUT127), .ZN(new_n996));
  INV_X1    g795(.A(KEYINPUT127), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n991), .A2(new_n997), .A3(new_n994), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n996), .A2(new_n998), .ZN(G1352gat));
  INV_X1    g798(.A(G204gat), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n692), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g800(.A(KEYINPUT62), .B1(new_n993), .B2(new_n1001), .ZN(new_n1002));
  OR3_X1    g801(.A1(new_n993), .A2(KEYINPUT62), .A3(new_n1001), .ZN(new_n1003));
  AND3_X1   g802(.A1(new_n946), .A2(new_n692), .A3(new_n989), .ZN(new_n1004));
  OAI211_X1 g803(.A(new_n1002), .B(new_n1003), .C1(new_n1004), .C2(new_n1000), .ZN(G1353gat));
  INV_X1    g804(.A(new_n993), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n1006), .A2(new_n376), .A3(new_n695), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n946), .A2(new_n695), .A3(new_n989), .ZN(new_n1008));
  AND3_X1   g807(.A1(new_n1008), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1009));
  AOI21_X1  g808(.A(KEYINPUT63), .B1(new_n1008), .B2(G211gat), .ZN(new_n1010));
  OAI21_X1  g809(.A(new_n1007), .B1(new_n1009), .B2(new_n1010), .ZN(G1354gat));
  NAND3_X1  g810(.A1(new_n1006), .A2(new_n377), .A3(new_n731), .ZN(new_n1012));
  AND3_X1   g811(.A1(new_n946), .A2(new_n731), .A3(new_n989), .ZN(new_n1013));
  OAI21_X1  g812(.A(new_n1012), .B1(new_n1013), .B2(new_n377), .ZN(G1355gat));
endmodule


