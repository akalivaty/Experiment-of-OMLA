//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 0 1 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1286, new_n1287, new_n1288, new_n1289, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n206), .A2(new_n207), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(KEYINPUT65), .B(G238), .ZN(new_n220));
  AND2_X1   g0020(.A1(new_n220), .A2(G68), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G107), .A2(G264), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n211), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n214), .B(new_n219), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(G41), .ZN(new_n246));
  AND2_X1   g0046(.A1(KEYINPUT76), .A2(KEYINPUT5), .ZN(new_n247));
  NOR2_X1   g0047(.A1(KEYINPUT76), .A2(KEYINPUT5), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT77), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  OAI211_X1 g0051(.A(KEYINPUT77), .B(new_n246), .C1(new_n247), .C2(new_n248), .ZN(new_n252));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G45), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT5), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n254), .B1(new_n255), .B2(G41), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n251), .A2(new_n252), .A3(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(G1), .A2(G13), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n257), .A2(G257), .A3(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT79), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT4), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  OAI21_X1  g0065(.A(KEYINPUT73), .B1(new_n265), .B2(KEYINPUT3), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT73), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT3), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(new_n268), .A3(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n266), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT66), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT66), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G1698), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n273), .A2(new_n275), .A3(G244), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n264), .B1(new_n271), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n268), .A2(G33), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n278), .A2(new_n270), .A3(G250), .A4(G1698), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G283), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT66), .B(G1698), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT3), .B(G33), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT4), .A4(G244), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n277), .A2(new_n281), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT78), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT76), .B(KEYINPUT5), .ZN(new_n289));
  AOI21_X1  g0089(.A(KEYINPUT77), .B1(new_n289), .B2(new_n246), .ZN(new_n290));
  INV_X1    g0090(.A(new_n252), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n288), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n251), .A2(KEYINPUT78), .A3(new_n252), .ZN(new_n293));
  INV_X1    g0093(.A(G274), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n294), .B1(new_n258), .B2(new_n259), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n256), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n292), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n257), .A2(KEYINPUT79), .A3(G257), .A4(new_n260), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n263), .A2(new_n287), .A3(new_n297), .A4(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT80), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n293), .A2(new_n296), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n302), .A2(new_n292), .B1(new_n286), .B2(new_n285), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n303), .A2(KEYINPUT80), .A3(new_n298), .A4(new_n263), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G169), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n216), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT6), .ZN(new_n310));
  INV_X1    g0110(.A(G97), .ZN(new_n311));
  NOR3_X1   g0111(.A1(new_n310), .A2(new_n311), .A3(G107), .ZN(new_n312));
  XNOR2_X1  g0112(.A(G97), .B(G107), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n312), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G77), .ZN(new_n315));
  NOR2_X1   g0115(.A1(G20), .A2(G33), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n314), .A2(new_n217), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G107), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT7), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(new_n283), .B2(G20), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n278), .A2(new_n270), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n322), .A2(KEYINPUT7), .A3(new_n217), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n319), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n309), .B1(new_n318), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n253), .A2(G13), .A3(G20), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n311), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n308), .A2(new_n216), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n329), .B(new_n326), .C1(G1), .C2(new_n265), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G97), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n325), .A2(new_n328), .A3(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n299), .B2(G179), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n301), .A2(new_n304), .A3(G190), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n333), .B1(new_n299), .B2(G200), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n307), .A2(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n208), .A2(G20), .ZN(new_n339));
  INV_X1    g0139(.A(G150), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT8), .B(G58), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n341), .B(KEYINPUT67), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n217), .A2(G33), .ZN(new_n343));
  OAI221_X1 g0143(.A(new_n339), .B1(new_n340), .B2(new_n317), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n309), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n329), .B1(G1), .B2(new_n217), .ZN(new_n346));
  MUX2_X1   g0146(.A(new_n326), .B(new_n346), .S(G50), .Z(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G45), .ZN(new_n349));
  AOI21_X1  g0149(.A(G1), .B1(new_n246), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n295), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n253), .B1(G41), .B2(G45), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n260), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G226), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n351), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n283), .A2(G223), .A3(G1698), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n282), .A2(new_n283), .ZN(new_n357));
  INV_X1    g0157(.A(G222), .ZN(new_n358));
  OAI221_X1 g0158(.A(new_n356), .B1(new_n315), .B2(new_n283), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n355), .B1(new_n359), .B2(new_n286), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n348), .B1(G169), .B2(new_n360), .ZN(new_n361));
  OR2_X1    g0161(.A1(new_n361), .A2(KEYINPUT68), .ZN(new_n362));
  INV_X1    g0162(.A(G179), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n361), .A2(KEYINPUT68), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n362), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G200), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n360), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g0169(.A(new_n369), .B(KEYINPUT70), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT9), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n348), .A2(new_n371), .B1(G190), .B2(new_n360), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n370), .B(new_n372), .C1(new_n371), .C2(new_n348), .ZN(new_n373));
  OR2_X1    g0173(.A1(new_n373), .A2(KEYINPUT10), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(KEYINPUT10), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n367), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  OAI22_X1  g0177(.A1(new_n317), .A2(new_n207), .B1(new_n217), .B2(G68), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n343), .A2(new_n315), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n309), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT11), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n380), .A2(new_n381), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT12), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n385), .B1(new_n327), .B2(new_n203), .ZN(new_n386));
  NOR3_X1   g0186(.A1(new_n326), .A2(KEYINPUT12), .A3(G68), .ZN(new_n387));
  OAI22_X1  g0187(.A1(new_n346), .A2(new_n203), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NOR3_X1   g0188(.A1(new_n383), .A2(new_n384), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n351), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n286), .A2(new_n350), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n391), .B1(G238), .B2(new_n392), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n278), .A2(new_n270), .A3(G232), .A4(G1698), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT71), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT71), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n283), .A2(new_n396), .A3(G232), .A4(G1698), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n282), .A2(new_n283), .A3(G226), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G33), .A2(G97), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n395), .A2(new_n397), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n400), .A2(KEYINPUT72), .A3(new_n286), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT72), .B1(new_n400), .B2(new_n286), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n393), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT13), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT13), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n405), .B(new_n393), .C1(new_n401), .C2(new_n402), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(G179), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n400), .A2(new_n286), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT72), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n400), .A2(KEYINPUT72), .A3(new_n286), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n405), .B1(new_n412), .B2(new_n393), .ZN(new_n413));
  INV_X1    g0213(.A(new_n406), .ZN(new_n414));
  OAI21_X1  g0214(.A(G169), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n407), .B1(new_n415), .B2(KEYINPUT14), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT14), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n404), .A2(new_n406), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n417), .B1(new_n418), .B2(G169), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n390), .B1(new_n416), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(G190), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n389), .B1(new_n418), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n368), .B1(new_n404), .B2(new_n406), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n392), .A2(G232), .B1(new_n295), .B2(new_n350), .ZN(new_n427));
  INV_X1    g0227(.A(G87), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n265), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n273), .A2(new_n275), .A3(G223), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G226), .A2(G1698), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n266), .A2(new_n269), .A3(new_n270), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n429), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI211_X1 g0234(.A(G179), .B(new_n427), .C1(new_n434), .C2(new_n260), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT75), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n351), .B1(new_n231), .B2(new_n353), .ZN(new_n437));
  INV_X1    g0237(.A(new_n429), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n282), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n438), .B1(new_n439), .B2(new_n271), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n437), .B1(new_n440), .B2(new_n286), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n435), .B(new_n436), .C1(new_n441), .C2(new_n306), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n432), .A2(new_n433), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n260), .B1(new_n444), .B2(new_n438), .ZN(new_n445));
  OAI21_X1  g0245(.A(G169), .B1(new_n445), .B2(new_n437), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n436), .B1(new_n446), .B2(new_n435), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT18), .ZN(new_n449));
  INV_X1    g0249(.A(new_n342), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n346), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(new_n327), .B2(new_n450), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n271), .A2(new_n217), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT7), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n271), .A2(new_n320), .A3(new_n217), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n454), .A2(G68), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G58), .A2(G68), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n204), .A2(new_n205), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G20), .ZN(new_n459));
  INV_X1    g0259(.A(G159), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n460), .A2(G20), .A3(G33), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT74), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n461), .B1(new_n458), .B2(G20), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT74), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n456), .A2(KEYINPUT16), .A3(new_n464), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n309), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n465), .A2(new_n466), .ZN(new_n470));
  AOI211_X1 g0270(.A(KEYINPUT74), .B(new_n461), .C1(new_n458), .C2(G20), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n203), .B1(new_n321), .B2(new_n323), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT16), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n452), .B1(new_n469), .B2(new_n475), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n448), .A2(new_n449), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n449), .B1(new_n448), .B2(new_n476), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR3_X1   g0279(.A1(new_n470), .A2(new_n471), .A3(new_n473), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n468), .B(new_n309), .C1(KEYINPUT16), .C2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n441), .A2(new_n421), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(G200), .B2(new_n441), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n481), .A2(new_n452), .A3(new_n483), .ZN(new_n484));
  XNOR2_X1  g0284(.A(new_n484), .B(KEYINPUT17), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G20), .A2(G77), .ZN(new_n487));
  XNOR2_X1  g0287(.A(KEYINPUT15), .B(G87), .ZN(new_n488));
  OAI221_X1 g0288(.A(new_n487), .B1(new_n488), .B2(new_n343), .C1(new_n317), .C2(new_n341), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n309), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n327), .A2(new_n315), .ZN(new_n491));
  OR2_X1    g0291(.A1(new_n346), .A2(new_n315), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n220), .A2(new_n283), .A3(G1698), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n322), .A2(G107), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n494), .B(new_n495), .C1(new_n357), .C2(new_n231), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n286), .ZN(new_n497));
  INV_X1    g0297(.A(G244), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n351), .B1(new_n353), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n493), .B1(G200), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(new_n421), .B2(new_n501), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n491), .B1(new_n346), .B2(new_n315), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n504), .B1(new_n309), .B2(new_n489), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n505), .B1(new_n501), .B2(new_n306), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n499), .B1(new_n496), .B2(new_n286), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n507), .A2(KEYINPUT69), .A3(new_n363), .ZN(new_n508));
  AOI21_X1  g0308(.A(KEYINPUT69), .B1(new_n507), .B2(new_n363), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n506), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n503), .A2(new_n510), .ZN(new_n511));
  NOR4_X1   g0311(.A1(new_n377), .A2(new_n426), .A3(new_n486), .A4(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n254), .A2(G274), .ZN(new_n513));
  AOI21_X1  g0313(.A(G250), .B1(new_n253), .B2(G45), .ZN(new_n514));
  NOR3_X1   g0314(.A1(new_n513), .A2(new_n286), .A3(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(G116), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT81), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT81), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G116), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G33), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n282), .A2(G238), .B1(G244), .B2(G1698), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n521), .B1(new_n522), .B2(new_n271), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n515), .B1(new_n523), .B2(new_n286), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n524), .A2(G169), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n525), .B1(new_n363), .B2(new_n524), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n266), .A2(new_n269), .A3(new_n217), .A4(new_n270), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT19), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n428), .A2(new_n311), .A3(new_n319), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n399), .A2(new_n217), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR3_X1   g0331(.A1(new_n343), .A2(KEYINPUT19), .A3(new_n311), .ZN(new_n532));
  OAI22_X1  g0332(.A1(new_n203), .A2(new_n527), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n533), .A2(new_n309), .B1(new_n327), .B2(new_n488), .ZN(new_n534));
  INV_X1    g0334(.A(new_n488), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n331), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT82), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT82), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n534), .A2(new_n539), .A3(new_n536), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n331), .A2(G87), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n534), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n524), .A2(new_n368), .ZN(new_n544));
  AOI211_X1 g0344(.A(new_n421), .B(new_n515), .C1(new_n523), .C2(new_n286), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n526), .A2(new_n541), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT83), .ZN(new_n548));
  AOI21_X1  g0348(.A(KEYINPUT25), .B1(new_n327), .B2(new_n319), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n327), .A2(KEYINPUT25), .A3(new_n319), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n331), .A2(G107), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT22), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n217), .A2(G87), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n553), .B1(new_n322), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT23), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n217), .B2(G107), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n319), .A2(KEYINPUT23), .A3(G20), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n555), .B(new_n559), .C1(new_n521), .C2(G20), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n527), .A2(new_n553), .A3(new_n428), .ZN(new_n561));
  OAI21_X1  g0361(.A(KEYINPUT24), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  XNOR2_X1  g0362(.A(KEYINPUT81), .B(G116), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n563), .A2(new_n265), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n564), .A2(new_n217), .B1(new_n557), .B2(new_n558), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n433), .A2(KEYINPUT22), .A3(new_n217), .A4(G87), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT24), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n565), .A2(new_n566), .A3(new_n567), .A4(new_n555), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n562), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n548), .B(new_n552), .C1(new_n569), .C2(new_n329), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n329), .B1(new_n562), .B2(new_n568), .ZN(new_n571));
  INV_X1    g0371(.A(new_n552), .ZN(new_n572));
  OAI21_X1  g0372(.A(KEYINPUT83), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n282), .A2(G250), .B1(G257), .B2(G1698), .ZN(new_n574));
  INV_X1    g0374(.A(G294), .ZN(new_n575));
  OAI22_X1  g0375(.A1(new_n574), .A2(new_n271), .B1(new_n265), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n286), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n257), .A2(G264), .A3(new_n260), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n297), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n579), .A2(KEYINPUT84), .A3(G169), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n297), .A2(new_n577), .A3(G179), .A4(new_n578), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(KEYINPUT84), .B1(new_n579), .B2(G169), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n570), .B(new_n573), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  OAI22_X1  g0384(.A1(new_n330), .A2(new_n516), .B1(new_n326), .B2(new_n520), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n517), .A2(new_n519), .A3(G20), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n280), .B(new_n217), .C1(G33), .C2(new_n311), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n309), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT20), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n587), .A2(KEYINPUT20), .A3(new_n309), .A4(new_n588), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n586), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G179), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n282), .A2(G257), .B1(G264), .B2(G1698), .ZN(new_n596));
  INV_X1    g0396(.A(G303), .ZN(new_n597));
  OAI22_X1  g0397(.A1(new_n596), .A2(new_n271), .B1(new_n597), .B2(new_n283), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n286), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n257), .A2(G270), .A3(new_n260), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n297), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n595), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n306), .B1(new_n586), .B2(new_n593), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n601), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(KEYINPUT21), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT21), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n603), .A2(new_n601), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n602), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n571), .A2(new_n572), .ZN(new_n609));
  OR2_X1    g0409(.A1(new_n579), .A2(new_n421), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n579), .A2(G200), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n594), .B1(new_n601), .B2(G200), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n421), .B2(new_n601), .ZN(new_n614));
  AND4_X1   g0414(.A1(new_n584), .A2(new_n608), .A3(new_n612), .A4(new_n614), .ZN(new_n615));
  AND4_X1   g0415(.A1(new_n338), .A2(new_n512), .A3(new_n547), .A4(new_n615), .ZN(G372));
  NAND2_X1  g0416(.A1(new_n336), .A2(new_n337), .ZN(new_n617));
  AOI21_X1  g0417(.A(G169), .B1(new_n301), .B2(new_n304), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n617), .B(new_n547), .C1(new_n618), .C2(new_n334), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n603), .A2(new_n601), .A3(new_n606), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n606), .B1(new_n603), .B2(new_n601), .ZN(new_n621));
  OAI22_X1  g0421(.A1(new_n620), .A2(new_n621), .B1(new_n601), .B2(new_n595), .ZN(new_n622));
  INV_X1    g0422(.A(new_n609), .ZN(new_n623));
  INV_X1    g0423(.A(new_n583), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n624), .A2(new_n581), .A3(new_n580), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n622), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n612), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n619), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n526), .A2(new_n541), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n334), .B1(new_n305), .B2(new_n306), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n630), .A2(KEYINPUT26), .A3(new_n547), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT26), .B1(new_n630), .B2(new_n547), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n512), .B1(new_n628), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n374), .A2(new_n375), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT17), .ZN(new_n636));
  XNOR2_X1  g0436(.A(new_n484), .B(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n493), .B1(G169), .B2(new_n507), .ZN(new_n638));
  INV_X1    g0438(.A(new_n509), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n507), .A2(KEYINPUT69), .A3(new_n363), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n425), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n637), .B1(new_n642), .B2(new_n420), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n481), .A2(new_n452), .B1(new_n446), .B2(new_n435), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n644), .B(new_n449), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n635), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n646), .A2(new_n366), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n634), .A2(new_n647), .ZN(G369));
  NAND3_X1  g0448(.A1(new_n253), .A2(new_n217), .A3(G13), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n650), .A2(G213), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT85), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n653), .A2(G343), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(G343), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g0457(.A(new_n657), .B(KEYINPUT86), .Z(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n594), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n608), .A2(new_n614), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n622), .A2(new_n594), .A3(new_n659), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT87), .ZN(new_n665));
  INV_X1    g0465(.A(G330), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(KEYINPUT87), .B1(new_n663), .B2(G330), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n570), .A2(new_n573), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n659), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n672), .A2(new_n584), .A3(new_n612), .ZN(new_n673));
  INV_X1    g0473(.A(new_n584), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n659), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n670), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n608), .A2(new_n659), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n678), .A2(new_n584), .A3(new_n612), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n625), .A2(new_n623), .A3(new_n658), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n677), .A2(new_n681), .ZN(G399));
  NOR2_X1   g0482(.A1(new_n529), .A2(G116), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n212), .A2(new_n246), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(new_n684), .A3(G1), .ZN(new_n685));
  INV_X1    g0485(.A(new_n215), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n685), .B1(new_n686), .B2(new_n684), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT28), .ZN(new_n688));
  INV_X1    g0488(.A(new_n629), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n307), .A2(new_n547), .A3(new_n335), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT26), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n630), .A2(KEYINPUT26), .A3(new_n547), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n689), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n625), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n608), .B1(new_n695), .B2(new_n609), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n696), .A2(new_n338), .A3(new_n547), .A4(new_n612), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n659), .B1(new_n694), .B2(new_n697), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n698), .A2(KEYINPUT29), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n622), .B1(new_n671), .B2(new_n625), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n619), .A2(new_n700), .A3(new_n627), .ZN(new_n701));
  OAI211_X1 g0501(.A(KEYINPUT29), .B(new_n658), .C1(new_n633), .C2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n524), .A2(new_n600), .A3(new_n599), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n581), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n301), .A2(new_n304), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT30), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n524), .A2(G179), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n708), .A2(new_n579), .A3(new_n601), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n706), .A2(new_n707), .B1(new_n299), .B2(new_n709), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n301), .A2(new_n304), .A3(new_n705), .A4(KEYINPUT30), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n658), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(KEYINPUT31), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n713), .A2(KEYINPUT88), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(KEYINPUT88), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n710), .A2(new_n711), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n659), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT31), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n615), .A2(new_n338), .A3(new_n547), .A4(new_n658), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n714), .A2(new_n715), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G330), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n703), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n688), .B1(new_n724), .B2(G1), .ZN(G364));
  INV_X1    g0525(.A(new_n684), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n217), .A2(G13), .ZN(new_n727));
  XOR2_X1   g0527(.A(new_n727), .B(KEYINPUT89), .Z(new_n728));
  AOI21_X1  g0528(.A(new_n253), .B1(new_n728), .B2(G45), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OAI221_X1 g0530(.A(new_n669), .B1(G330), .B2(new_n663), .C1(new_n726), .C2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n726), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n283), .A2(new_n212), .ZN(new_n733));
  INV_X1    g0533(.A(G355), .ZN(new_n734));
  OAI22_X1  g0534(.A1(new_n733), .A2(new_n734), .B1(G116), .B2(new_n212), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n241), .A2(new_n349), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n271), .A2(new_n212), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n737), .B1(new_n349), .B2(new_n215), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n735), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n258), .B1(new_n217), .B2(G169), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n740), .A2(KEYINPUT90), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(KEYINPUT90), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G13), .A2(G33), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n732), .B1(new_n739), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n217), .A2(new_n363), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n750), .A2(G190), .A3(new_n368), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(G200), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G190), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI221_X1 g0554(.A(new_n283), .B1(new_n202), .B2(new_n751), .C1(new_n754), .C2(new_n203), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n217), .A2(G179), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n756), .A2(new_n421), .A3(G200), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n319), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n752), .A2(new_n421), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n758), .B1(G50), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n756), .A2(G190), .A3(G200), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n760), .B1(new_n428), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G190), .A2(G200), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n750), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n765), .A2(KEYINPUT91), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(KEYINPUT91), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n755), .B(new_n762), .C1(G77), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n756), .A2(new_n763), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n771), .A2(KEYINPUT92), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(KEYINPUT92), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n460), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT32), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n421), .A2(G179), .A3(G200), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n217), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT93), .Z(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n770), .B(new_n776), .C1(new_n311), .C2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT94), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n759), .B(KEYINPUT95), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  XOR2_X1   g0585(.A(KEYINPUT96), .B(G326), .Z(new_n786));
  XOR2_X1   g0586(.A(new_n761), .B(KEYINPUT97), .Z(new_n787));
  AOI22_X1  g0587(.A1(new_n785), .A2(new_n786), .B1(new_n787), .B2(G303), .ZN(new_n788));
  INV_X1    g0588(.A(new_n751), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n283), .B1(new_n789), .B2(G322), .ZN(new_n790));
  INV_X1    g0590(.A(G311), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n790), .B1(new_n791), .B2(new_n764), .ZN(new_n792));
  INV_X1    g0592(.A(new_n774), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n792), .B1(new_n793), .B2(G329), .ZN(new_n794));
  INV_X1    g0594(.A(new_n757), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G283), .ZN(new_n796));
  INV_X1    g0596(.A(new_n778), .ZN(new_n797));
  XNOR2_X1  g0597(.A(KEYINPUT33), .B(G317), .ZN(new_n798));
  AOI22_X1  g0598(.A1(G294), .A2(new_n797), .B1(new_n753), .B2(new_n798), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n788), .A2(new_n794), .A3(new_n796), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n781), .A2(new_n782), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n783), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n749), .B1(new_n802), .B2(new_n743), .ZN(new_n803));
  INV_X1    g0603(.A(new_n746), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n803), .B1(new_n663), .B2(new_n804), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n731), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(G396));
  OAI211_X1 g0607(.A(new_n503), .B(new_n510), .C1(new_n505), .C2(new_n658), .ZN(new_n808));
  AOI21_X1  g0608(.A(KEYINPUT99), .B1(new_n641), .B2(new_n659), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT99), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n510), .A2(new_n810), .A3(new_n658), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n808), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(KEYINPUT100), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT100), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n814), .B(new_n808), .C1(new_n809), .C2(new_n811), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n698), .B(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n732), .B1(new_n817), .B2(new_n722), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n722), .B2(new_n817), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n743), .A2(new_n744), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n726), .B(new_n730), .C1(new_n315), .C2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n743), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n757), .A2(new_n203), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n271), .B(new_n823), .C1(G58), .C2(new_n797), .ZN(new_n824));
  INV_X1    g0624(.A(G132), .ZN(new_n825));
  INV_X1    g0625(.A(new_n787), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n824), .B1(new_n825), .B2(new_n774), .C1(new_n826), .C2(new_n207), .ZN(new_n827));
  AOI22_X1  g0627(.A1(G137), .A2(new_n759), .B1(new_n789), .B2(G143), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n340), .B2(new_n754), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(G159), .B2(new_n769), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n827), .B1(KEYINPUT34), .B2(new_n830), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n830), .A2(KEYINPUT34), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n768), .A2(new_n563), .B1(new_n791), .B2(new_n774), .ZN(new_n833));
  XNOR2_X1  g0633(.A(KEYINPUT98), .B(G283), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n322), .B1(new_n575), .B2(new_n751), .C1(new_n754), .C2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n795), .A2(G87), .ZN(new_n836));
  INV_X1    g0636(.A(new_n759), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n836), .B1(new_n837), .B2(new_n597), .ZN(new_n838));
  NOR3_X1   g0638(.A1(new_n833), .A2(new_n835), .A3(new_n838), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n779), .A2(G97), .B1(new_n787), .B2(G107), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n831), .A2(new_n832), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n821), .B1(new_n822), .B2(new_n841), .C1(new_n816), .C2(new_n745), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n819), .A2(new_n842), .ZN(G384));
  INV_X1    g0643(.A(new_n314), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n844), .A2(KEYINPUT35), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(KEYINPUT35), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n845), .A2(G116), .A3(new_n218), .A4(new_n846), .ZN(new_n847));
  XOR2_X1   g0647(.A(KEYINPUT101), .B(KEYINPUT36), .Z(new_n848));
  XNOR2_X1  g0648(.A(new_n847), .B(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n215), .A2(G77), .A3(new_n457), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n207), .A2(G68), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n253), .B(G13), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT38), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT16), .B1(new_n472), .B2(new_n456), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n452), .B1(new_n469), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n652), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(new_n479), .B2(new_n485), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n446), .A2(new_n435), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n857), .A2(new_n860), .A3(new_n484), .ZN(new_n861));
  AND3_X1   g0661(.A1(new_n481), .A2(new_n452), .A3(new_n483), .ZN(new_n862));
  INV_X1    g0662(.A(new_n652), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n481), .B2(new_n452), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT37), .B1(new_n448), .B2(new_n476), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n861), .A2(KEYINPUT37), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n854), .B1(new_n858), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT102), .ZN(new_n869));
  INV_X1    g0669(.A(new_n857), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n448), .A2(new_n476), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT18), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n448), .A2(new_n449), .A3(new_n476), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n870), .B1(new_n874), .B2(new_n637), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n861), .A2(KEYINPUT37), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n865), .A2(new_n866), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n875), .A2(KEYINPUT38), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n868), .A2(new_n869), .A3(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(KEYINPUT102), .B(new_n854), .C1(new_n858), .C2(new_n867), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n717), .A2(KEYINPUT106), .A3(new_n718), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT106), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n712), .B2(KEYINPUT31), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n882), .A2(new_n884), .A3(new_n713), .A4(new_n720), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n659), .A2(new_n390), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n420), .A2(new_n425), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n415), .A2(KEYINPUT14), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n418), .A2(new_n417), .A3(G169), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(new_n407), .A3(new_n889), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n390), .B(new_n659), .C1(new_n890), .C2(new_n424), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n887), .A2(new_n891), .B1(new_n815), .B2(new_n813), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n880), .A2(new_n881), .A3(new_n885), .A4(new_n892), .ZN(new_n893));
  XOR2_X1   g0693(.A(KEYINPUT105), .B(KEYINPUT40), .Z(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n476), .A2(new_n652), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n644), .B(KEYINPUT18), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n896), .B1(new_n897), .B2(new_n485), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n476), .A2(new_n859), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n899), .A2(new_n896), .A3(new_n484), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT103), .B1(new_n900), .B2(KEYINPUT37), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n865), .A2(new_n866), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n900), .A2(KEYINPUT103), .A3(KEYINPUT37), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n898), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n879), .B1(new_n905), .B2(KEYINPUT38), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n906), .A2(KEYINPUT40), .A3(new_n885), .A4(new_n892), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n895), .A2(G330), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n512), .A2(G330), .A3(new_n885), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n911), .A2(KEYINPUT107), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT40), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n900), .A2(KEYINPUT103), .A3(KEYINPUT37), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n914), .A2(new_n901), .A3(new_n902), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n854), .B1(new_n915), .B2(new_n898), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n913), .B1(new_n916), .B2(new_n879), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n885), .A2(new_n892), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n893), .A2(new_n894), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(new_n512), .A3(new_n885), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n911), .A2(KEYINPUT107), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n912), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n923), .B(new_n879), .C1(new_n905), .C2(KEYINPUT38), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT104), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n880), .A2(KEYINPUT39), .A3(new_n881), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT104), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n916), .A2(new_n927), .A3(new_n923), .A4(new_n879), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n890), .A2(new_n390), .A3(new_n658), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n658), .B(new_n816), .C1(new_n633), .C2(new_n628), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n641), .A2(new_n658), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n887), .A2(new_n891), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n935), .A2(new_n937), .A3(new_n881), .A4(new_n880), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n645), .A2(new_n863), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n932), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n512), .A2(new_n699), .A3(new_n702), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n647), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n942), .B(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n922), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n253), .B2(new_n728), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n922), .A2(new_n945), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n853), .B1(new_n947), .B2(new_n948), .ZN(G367));
  OAI21_X1  g0749(.A(new_n747), .B1(new_n212), .B2(new_n488), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n237), .A2(new_n737), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n732), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n761), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n753), .A2(G159), .B1(new_n953), .B2(G58), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n768), .B2(new_n207), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n795), .A2(G77), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT116), .B1(new_n956), .B2(new_n283), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n785), .B2(G143), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n956), .A2(KEYINPUT116), .A3(new_n283), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n955), .B(new_n960), .C1(G137), .C2(new_n793), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n779), .A2(G68), .B1(G150), .B2(new_n789), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT115), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n271), .B1(new_n751), .B2(new_n597), .ZN(new_n965));
  INV_X1    g0765(.A(new_n834), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n965), .B1(new_n769), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n761), .A2(new_n563), .ZN(new_n968));
  XOR2_X1   g0768(.A(KEYINPUT114), .B(G317), .Z(new_n969));
  OAI221_X1 g0769(.A(new_n967), .B1(KEYINPUT46), .B2(new_n968), .C1(new_n774), .C2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n785), .A2(G311), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n787), .A2(KEYINPUT46), .A3(G116), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n757), .A2(new_n311), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  AOI22_X1  g0774(.A1(G107), .A2(new_n797), .B1(new_n753), .B2(G294), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n971), .A2(new_n972), .A3(new_n974), .A4(new_n975), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n962), .A2(new_n964), .B1(new_n970), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n978), .A2(KEYINPUT47), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n822), .B1(new_n978), .B2(KEYINPUT47), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n952), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n658), .A2(new_n543), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n547), .A2(new_n982), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n983), .A2(KEYINPUT108), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(KEYINPUT108), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n982), .A2(new_n629), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n987), .A2(new_n804), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n981), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT113), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n987), .B(KEYINPUT43), .Z(new_n991));
  INV_X1    g0791(.A(KEYINPUT42), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n307), .A2(new_n335), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n659), .A2(new_n333), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n993), .A2(new_n617), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n630), .A2(new_n659), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n679), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT110), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n999), .B1(new_n997), .B2(new_n998), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n992), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n997), .A2(new_n998), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(KEYINPUT110), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1005), .A2(KEYINPUT42), .A3(new_n1000), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n995), .A2(KEYINPUT109), .A3(new_n996), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(KEYINPUT109), .B1(new_n995), .B2(new_n996), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n674), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n659), .B1(new_n1011), .B2(new_n993), .ZN(new_n1012));
  OAI211_X1 g0812(.A(KEYINPUT111), .B(new_n991), .C1(new_n1007), .C2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1010), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n584), .B1(new_n1014), .B2(new_n1008), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n658), .B1(new_n1015), .B2(new_n630), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n987), .A2(KEYINPUT43), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1016), .A2(new_n1006), .A3(new_n1003), .A4(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1013), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1016), .A2(new_n1006), .A3(new_n1003), .ZN(new_n1020));
  AOI21_X1  g0820(.A(KEYINPUT111), .B1(new_n1020), .B2(new_n991), .ZN(new_n1021));
  OAI21_X1  g0821(.A(KEYINPUT112), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n991), .B1(new_n1007), .B2(new_n1012), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT111), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT112), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1025), .A2(new_n1026), .A3(new_n1018), .A4(new_n1013), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1022), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1014), .A2(new_n1008), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n677), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1031), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1022), .A2(new_n1033), .A3(new_n1027), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n681), .A2(new_n997), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT44), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n681), .A2(new_n997), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT45), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1038), .B(new_n1039), .ZN(new_n1040));
  AND3_X1   g0840(.A1(new_n1037), .A2(new_n677), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n677), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n679), .B1(new_n676), .B2(new_n678), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n669), .B(new_n1044), .Z(new_n1045));
  AOI21_X1  g0845(.A(new_n723), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n684), .B(KEYINPUT41), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n729), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n990), .B1(new_n1035), .B2(new_n1048), .ZN(new_n1049));
  AND3_X1   g0849(.A1(new_n1022), .A2(new_n1033), .A3(new_n1027), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1033), .B1(new_n1022), .B2(new_n1027), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n990), .B(new_n1048), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n989), .B1(new_n1049), .B2(new_n1053), .ZN(G387));
  NAND3_X1  g0854(.A1(new_n673), .A2(new_n675), .A3(new_n746), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n733), .A2(new_n683), .B1(G107), .B2(new_n212), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n234), .A2(new_n349), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n683), .ZN(new_n1058));
  AOI211_X1 g0858(.A(G45), .B(new_n1058), .C1(G68), .C2(G77), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n341), .A2(G50), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT50), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n737), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1056), .B1(new_n1057), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n732), .B1(new_n1063), .B2(new_n748), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n759), .A2(G159), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT117), .Z(new_n1066));
  AOI22_X1  g0866(.A1(new_n793), .A2(G150), .B1(new_n450), .B2(new_n753), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n779), .A2(new_n535), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n751), .A2(new_n207), .B1(new_n764), .B2(new_n203), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n761), .A2(new_n315), .ZN(new_n1070));
  NOR4_X1   g0870(.A1(new_n1069), .A2(new_n973), .A3(new_n1070), .A4(new_n271), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .A4(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n785), .A2(G322), .B1(G311), .B2(new_n753), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1074), .A2(KEYINPUT118), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n768), .A2(new_n597), .B1(new_n751), .B2(new_n969), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(KEYINPUT118), .B2(new_n1074), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT48), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n778), .A2(new_n834), .B1(new_n761), .B2(new_n575), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1080), .A2(KEYINPUT49), .A3(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n271), .B1(new_n757), .B2(new_n563), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n793), .B2(new_n786), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(KEYINPUT49), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1072), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1064), .B1(new_n1088), .B2(new_n743), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n1055), .A2(new_n1089), .B1(new_n1045), .B2(new_n730), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n724), .A2(new_n1045), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n726), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n724), .A2(new_n1045), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1090), .B1(new_n1092), .B2(new_n1093), .ZN(G393));
  OAI21_X1  g0894(.A(new_n747), .B1(new_n311), .B2(new_n212), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n244), .A2(new_n737), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n732), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n341), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n769), .A2(new_n1098), .B1(G143), .B2(new_n793), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n753), .A2(G50), .B1(new_n953), .B2(G68), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1099), .A2(new_n433), .A3(new_n836), .A4(new_n1100), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n837), .A2(new_n340), .B1(new_n460), .B2(new_n751), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT51), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n779), .A2(G77), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n793), .A2(G322), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n283), .B(new_n758), .C1(G294), .C2(new_n765), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n797), .A2(new_n520), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n753), .A2(G303), .B1(new_n953), .B2(new_n966), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(G317), .A2(new_n759), .B1(new_n789), .B2(G311), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT52), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n1101), .A2(new_n1107), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1097), .B1(new_n1115), .B2(new_n743), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n1029), .B2(new_n804), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1043), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1117), .B1(new_n1118), .B2(new_n729), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1118), .A2(new_n1091), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1120), .A2(new_n684), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1118), .A2(new_n1091), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1119), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(G390));
  OAI211_X1 g0924(.A(new_n658), .B(new_n816), .C1(new_n633), .C2(new_n701), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n934), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n937), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n931), .B1(new_n916), .B2(new_n879), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1127), .A2(new_n1128), .A3(KEYINPUT119), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT119), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n936), .B1(new_n934), .B2(new_n1125), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT103), .ZN(new_n1132));
  NOR3_X1   g0932(.A1(new_n862), .A2(new_n644), .A3(new_n864), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT37), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1135), .A2(new_n877), .A3(new_n904), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n864), .B1(new_n645), .B2(new_n637), .ZN(new_n1137));
  AOI21_X1  g0937(.A(KEYINPUT38), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NOR3_X1   g0938(.A1(new_n858), .A2(new_n854), .A3(new_n867), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n930), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1130), .B1(new_n1131), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1129), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n934), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n698), .B2(new_n816), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n930), .B1(new_n1144), .B2(new_n936), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1145), .A2(new_n925), .A3(new_n926), .A4(new_n928), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n666), .B1(new_n813), .B2(new_n815), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n721), .A2(new_n937), .A3(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1142), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n1142), .A2(new_n1146), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n885), .A2(new_n1147), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1151), .A2(new_n936), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1149), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(KEYINPUT120), .B1(new_n1154), .B2(new_n729), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n1142), .A2(new_n1148), .A3(new_n1146), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1153), .B1(new_n1142), .B2(new_n1146), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT120), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1158), .A2(new_n1159), .A3(new_n730), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1155), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n937), .B1(new_n721), .B2(new_n1147), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n935), .B1(new_n1162), .B2(new_n1152), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1126), .B1(new_n936), .B2(new_n1151), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n1148), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n943), .A2(new_n909), .A3(new_n647), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1154), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1167), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1149), .B(new_n1171), .C1(new_n1150), .C2(new_n1153), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1170), .A2(new_n726), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n820), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n732), .B1(new_n1174), .B2(new_n450), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n769), .A2(G97), .B1(G294), .B2(new_n793), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n283), .B(new_n823), .C1(G116), .C2(new_n789), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(G107), .A2(new_n753), .B1(new_n759), .B2(G283), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1105), .B1(new_n428), .B2(new_n826), .ZN(new_n1180));
  XOR2_X1   g0980(.A(KEYINPUT54), .B(G143), .Z(new_n1181));
  NAND2_X1  g0981(.A1(new_n769), .A2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n283), .B1(new_n751), .B2(new_n825), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(G128), .B2(new_n759), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n753), .A2(G137), .B1(new_n795), .B2(G50), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n793), .A2(G125), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1182), .A2(new_n1184), .A3(new_n1185), .A4(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n761), .A2(new_n340), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT53), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n780), .B2(new_n460), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n1179), .A2(new_n1180), .B1(new_n1187), .B2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1175), .B1(new_n1191), .B2(new_n743), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n929), .B2(new_n745), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1161), .A2(new_n1173), .A3(new_n1193), .ZN(G378));
  XNOR2_X1  g0994(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n348), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1197), .A2(new_n863), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n376), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n376), .A2(new_n1199), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1196), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1202), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1204), .A2(new_n1200), .A3(new_n1195), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n895), .A2(new_n1206), .A3(G330), .A4(new_n907), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1206), .B1(new_n919), .B2(G330), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n942), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1206), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n908), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n940), .B1(new_n929), .B2(new_n931), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1212), .A2(new_n1213), .A3(new_n1207), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1210), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1211), .A2(new_n744), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n732), .B1(new_n1174), .B2(G50), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n433), .A2(G41), .ZN(new_n1218));
  AOI211_X1 g1018(.A(G50), .B(new_n1218), .C1(new_n265), .C2(new_n246), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n757), .A2(new_n202), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n311), .A2(new_n754), .B1(new_n837), .B2(new_n516), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1220), .B(new_n1221), .C1(G68), .C2(new_n779), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n793), .A2(G283), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n751), .A2(new_n319), .B1(new_n764), .B2(new_n488), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1224), .A2(new_n1070), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1222), .A2(new_n1223), .A3(new_n1218), .A4(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT58), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1219), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n753), .A2(G132), .B1(new_n765), .B2(G137), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1229), .B(KEYINPUT121), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n779), .A2(G150), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n953), .A2(new_n1181), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(G125), .A2(new_n759), .B1(new_n789), .B2(G128), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .A4(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1234), .A2(KEYINPUT59), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(KEYINPUT59), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n793), .A2(G124), .ZN(new_n1237));
  AOI211_X1 g1037(.A(G33), .B(G41), .C1(new_n795), .C2(G159), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1228), .B1(new_n1227), .B2(new_n1226), .C1(new_n1235), .C2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1217), .B1(new_n1240), .B2(new_n743), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n1215), .A2(new_n730), .B1(new_n1216), .B2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1167), .B1(new_n1158), .B2(new_n1171), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1212), .A2(new_n1213), .A3(new_n1207), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n1212), .A2(new_n1207), .B1(new_n932), .B2(new_n941), .ZN(new_n1245));
  OAI21_X1  g1045(.A(KEYINPUT57), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(KEYINPUT122), .B1(new_n1243), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1172), .A2(new_n1168), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT122), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1248), .A2(new_n1249), .A3(KEYINPUT57), .A4(new_n1215), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1247), .A2(new_n1250), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1172), .A2(new_n1168), .B1(new_n1210), .B2(new_n1214), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n726), .B1(new_n1252), .B2(KEYINPUT57), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1242), .B1(new_n1251), .B2(new_n1253), .ZN(G375));
  INV_X1    g1054(.A(new_n1166), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1167), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1047), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1256), .A2(new_n1257), .A3(new_n1169), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n936), .A2(new_n744), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n732), .B1(new_n1174), .B2(G68), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n837), .A2(new_n825), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n1220), .B(new_n1261), .C1(new_n753), .C2(new_n1181), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n793), .A2(G128), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n764), .A2(new_n340), .ZN(new_n1264));
  AOI211_X1 g1064(.A(new_n271), .B(new_n1264), .C1(G137), .C2(new_n789), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1262), .A2(new_n1263), .A3(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n779), .A2(G50), .B1(new_n787), .B2(G159), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n769), .A2(G107), .B1(G303), .B2(new_n793), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n283), .B1(new_n789), .B2(G283), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(G294), .A2(new_n759), .B1(new_n753), .B2(new_n520), .ZN(new_n1271));
  AND4_X1   g1071(.A1(new_n956), .A2(new_n1269), .A3(new_n1270), .A4(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1068), .B1(new_n311), .B2(new_n826), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n1267), .A2(new_n1268), .B1(new_n1272), .B2(new_n1274), .ZN(new_n1275));
  OR2_X1    g1075(.A1(new_n1275), .A2(KEYINPUT123), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n822), .B1(new_n1275), .B2(KEYINPUT123), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1260), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(new_n1166), .A2(new_n730), .B1(new_n1259), .B2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1258), .A2(new_n1279), .ZN(G381));
  INV_X1    g1080(.A(G384), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1123), .A2(new_n1281), .ZN(new_n1282));
  OR4_X1    g1082(.A1(G396), .A2(new_n1282), .A3(G393), .A4(G381), .ZN(new_n1283));
  NOR4_X1   g1083(.A1(new_n1283), .A2(G375), .A3(G387), .A4(G378), .ZN(new_n1284));
  XOR2_X1   g1084(.A(new_n1284), .B(KEYINPUT124), .Z(G407));
  AND3_X1   g1085(.A1(new_n1161), .A2(new_n1173), .A3(new_n1193), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n654), .A2(new_n655), .A3(G213), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1289));
  OAI211_X1 g1089(.A(G407), .B(G213), .C1(G375), .C2(new_n1289), .ZN(G409));
  OAI211_X1 g1090(.A(G378), .B(new_n1242), .C1(new_n1251), .C2(new_n1253), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1252), .A2(new_n1257), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1216), .A2(new_n1241), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1215), .A2(KEYINPUT125), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n730), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1215), .A2(KEYINPUT125), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n1292), .B(new_n1293), .C1(new_n1295), .C2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1286), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1291), .A2(new_n1298), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1300), .B1(KEYINPUT60), .B2(new_n1169), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1255), .A2(KEYINPUT60), .A3(new_n1167), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n726), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1279), .B1(new_n1301), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1281), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1304), .A2(new_n1281), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1299), .A2(new_n1287), .A3(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT63), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(G393), .B(new_n806), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1048), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(KEYINPUT113), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(new_n1052), .ZN(new_n1316));
  AOI21_X1  g1116(.A(G390), .B1(new_n1316), .B2(new_n989), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n989), .ZN(new_n1318));
  AOI211_X1 g1118(.A(new_n1318), .B(new_n1123), .C1(new_n1315), .C2(new_n1052), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1313), .B1(new_n1317), .B2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(G387), .A2(new_n1123), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1316), .A2(new_n989), .A3(G390), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1321), .A2(new_n1312), .A3(new_n1322), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1320), .A2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1299), .A2(new_n1287), .ZN(new_n1325));
  OAI211_X1 g1125(.A(G2897), .B(new_n1288), .C1(new_n1306), .C2(new_n1307), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1307), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1288), .A2(G2897), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1327), .A2(new_n1305), .A3(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1326), .A2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1325), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT61), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1311), .A2(new_n1324), .A3(new_n1332), .A4(new_n1333), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1299), .A2(KEYINPUT63), .A3(new_n1287), .A4(new_n1308), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT126), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1288), .B1(new_n1291), .B2(new_n1298), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1338), .A2(KEYINPUT126), .A3(KEYINPUT63), .A4(new_n1308), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1337), .A2(new_n1339), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1334), .A2(new_n1340), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1333), .B1(new_n1338), .B2(new_n1330), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT62), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1343), .B1(new_n1338), .B2(new_n1308), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1342), .A2(new_n1344), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1338), .A2(new_n1343), .A3(new_n1308), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1324), .B1(new_n1345), .B2(new_n1346), .ZN(new_n1347));
  OAI21_X1  g1147(.A(KEYINPUT127), .B1(new_n1341), .B2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1309), .A2(KEYINPUT62), .ZN(new_n1349));
  NAND4_X1  g1149(.A1(new_n1349), .A2(new_n1332), .A3(new_n1333), .A4(new_n1346), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1324), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT127), .ZN(new_n1353));
  OAI211_X1 g1153(.A(new_n1352), .B(new_n1353), .C1(new_n1334), .C2(new_n1340), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1348), .A2(new_n1354), .ZN(G405));
  NAND2_X1  g1155(.A1(G375), .A2(new_n1286), .ZN(new_n1356));
  INV_X1    g1156(.A(new_n1356), .ZN(new_n1357));
  INV_X1    g1157(.A(new_n1291), .ZN(new_n1358));
  NOR2_X1   g1158(.A1(new_n1357), .A2(new_n1358), .ZN(new_n1359));
  XNOR2_X1  g1159(.A(new_n1359), .B(new_n1308), .ZN(new_n1360));
  XNOR2_X1  g1160(.A(new_n1360), .B(new_n1324), .ZN(G402));
endmodule


