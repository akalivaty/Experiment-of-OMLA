//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 1 1 0 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 0 1 0 1 0 1 1 1 1 0 0 0 0 1 1 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1007, new_n1008, new_n1009, new_n1010, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT70), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT70), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G237), .ZN(new_n191));
  AOI21_X1  g005(.A(G953), .B1(new_n189), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT85), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT85), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  AND3_X1   g011(.A1(new_n192), .A2(G214), .A3(new_n197), .ZN(new_n198));
  AOI22_X1  g012(.A1(new_n192), .A2(G214), .B1(new_n195), .B2(G143), .ZN(new_n199));
  OAI21_X1  g013(.A(G131), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT88), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT17), .ZN(new_n202));
  INV_X1    g016(.A(G953), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n190), .A2(G237), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n188), .A2(KEYINPUT70), .ZN(new_n205));
  OAI211_X1 g019(.A(G214), .B(new_n203), .C1(new_n204), .C2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(new_n196), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n192), .A2(G214), .A3(new_n197), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT88), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(G131), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n207), .A2(new_n212), .A3(new_n208), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n201), .A2(new_n202), .A3(new_n211), .A4(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n210), .B1(new_n209), .B2(G131), .ZN(new_n215));
  AOI211_X1 g029(.A(KEYINPUT88), .B(new_n212), .C1(new_n207), .C2(new_n208), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT17), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(G125), .B(G140), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT75), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT16), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n218), .A2(KEYINPUT16), .ZN(new_n221));
  INV_X1    g035(.A(G140), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G125), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT75), .B1(new_n223), .B2(KEYINPUT16), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n220), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G146), .ZN(new_n226));
  INV_X1    g040(.A(G146), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n227), .B(new_n220), .C1(new_n221), .C2(new_n224), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n214), .A2(new_n217), .A3(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(G113), .B(G122), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT90), .B(G104), .ZN(new_n233));
  XOR2_X1   g047(.A(new_n232), .B(new_n233), .Z(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT76), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n236), .B1(new_n218), .B2(new_n227), .ZN(new_n237));
  INV_X1    g051(.A(G125), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G140), .ZN(new_n239));
  AND4_X1   g053(.A1(new_n236), .A2(new_n223), .A3(new_n239), .A4(new_n227), .ZN(new_n240));
  OAI22_X1  g054(.A1(new_n237), .A2(new_n240), .B1(new_n227), .B2(new_n218), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT86), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT86), .ZN(new_n243));
  OAI221_X1 g057(.A(new_n243), .B1(new_n227), .B2(new_n218), .C1(new_n237), .C2(new_n240), .ZN(new_n244));
  NAND2_X1  g058(.A1(KEYINPUT18), .A2(G131), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  AOI22_X1  g060(.A1(new_n242), .A2(new_n244), .B1(new_n246), .B2(new_n209), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT87), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n248), .B1(new_n209), .B2(new_n246), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n207), .A2(KEYINPUT87), .A3(new_n208), .A4(new_n245), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n231), .A2(new_n235), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n235), .B1(new_n231), .B2(new_n252), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n187), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G475), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT91), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n193), .A2(G128), .ZN(new_n258));
  INV_X1    g072(.A(G128), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G143), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT13), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n257), .B(new_n258), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n259), .A2(G143), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n264), .B1(KEYINPUT13), .B2(new_n260), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT91), .B1(new_n258), .B2(new_n262), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n263), .B(G134), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n258), .A2(new_n260), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n268), .A2(G134), .ZN(new_n269));
  INV_X1    g083(.A(G116), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n270), .A2(G122), .ZN(new_n271));
  INV_X1    g085(.A(G122), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n272), .A2(G116), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G107), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(G107), .B1(new_n271), .B2(new_n273), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n269), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n267), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT92), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT92), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n267), .A2(new_n278), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT14), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n273), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n271), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(KEYINPUT93), .A3(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n273), .A2(new_n283), .ZN(new_n287));
  OAI221_X1 g101(.A(G107), .B1(KEYINPUT93), .B2(new_n284), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n269), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n268), .A2(G134), .ZN(new_n290));
  AOI22_X1  g104(.A1(new_n289), .A2(new_n290), .B1(new_n275), .B2(new_n274), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n280), .A2(new_n282), .A3(new_n292), .ZN(new_n293));
  XNOR2_X1  g107(.A(KEYINPUT9), .B(G234), .ZN(new_n294));
  INV_X1    g108(.A(G217), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n294), .A2(new_n295), .A3(G953), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n279), .A2(KEYINPUT92), .B1(new_n288), .B2(new_n291), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n299), .A2(new_n282), .A3(new_n296), .ZN(new_n300));
  AOI21_X1  g114(.A(G902), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G478), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n302), .A2(KEYINPUT15), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n301), .B(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT20), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n201), .A2(new_n211), .A3(new_n213), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n218), .A2(KEYINPUT16), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n307), .B(KEYINPUT75), .C1(KEYINPUT16), .C2(new_n223), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n227), .B1(new_n308), .B2(new_n220), .ZN(new_n309));
  XOR2_X1   g123(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(new_n218), .ZN(new_n311));
  NAND2_X1  g125(.A1(KEYINPUT89), .A2(KEYINPUT19), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n311), .B1(new_n218), .B2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n309), .B1(new_n227), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n306), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n252), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n234), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n231), .A2(new_n235), .A3(new_n252), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(G475), .A2(G902), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n305), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n320), .ZN(new_n322));
  AOI211_X1 g136(.A(KEYINPUT20), .B(new_n322), .C1(new_n317), .C2(new_n318), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n256), .B(new_n304), .C1(new_n321), .C2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G952), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n326), .A2(G953), .ZN(new_n327));
  NAND2_X1  g141(.A1(G234), .A2(G237), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  XOR2_X1   g143(.A(new_n329), .B(KEYINPUT94), .Z(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT21), .B(G898), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n328), .A2(G902), .A3(G953), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n330), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(G214), .B1(G237), .B2(G902), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(G110), .B(G122), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n340), .B(KEYINPUT8), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT83), .ZN(new_n342));
  INV_X1    g156(.A(G119), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT66), .B1(new_n343), .B2(G116), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT66), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(new_n270), .A3(G119), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n270), .A2(G119), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(KEYINPUT2), .B(G113), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT67), .ZN(new_n353));
  AOI211_X1 g167(.A(new_n353), .B(new_n348), .C1(new_n346), .C2(new_n344), .ZN(new_n354));
  AOI21_X1  g168(.A(KEYINPUT67), .B1(new_n347), .B2(new_n349), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT5), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(G113), .B1(new_n349), .B2(KEYINPUT5), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n352), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT3), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(new_n275), .A3(G104), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT79), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT79), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n363), .A2(new_n360), .A3(new_n275), .A4(G104), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n275), .A2(G104), .ZN(new_n366));
  INV_X1    g180(.A(G104), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT3), .B1(new_n367), .B2(G107), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT78), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n366), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G101), .ZN(new_n371));
  OAI211_X1 g185(.A(KEYINPUT78), .B(KEYINPUT3), .C1(new_n367), .C2(G107), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n365), .A2(new_n370), .A3(new_n371), .A4(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n367), .A2(G107), .ZN(new_n374));
  OAI21_X1  g188(.A(G101), .B1(new_n374), .B2(new_n366), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n342), .B1(new_n359), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n373), .A2(new_n375), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n348), .B1(new_n344), .B2(new_n346), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n357), .B1(new_n379), .B2(KEYINPUT5), .ZN(new_n380));
  OR3_X1    g194(.A1(new_n378), .A2(new_n352), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  NOR3_X1   g196(.A1(new_n359), .A2(new_n342), .A3(new_n376), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n341), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n227), .A2(G143), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n193), .A2(G146), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT1), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n385), .A2(new_n386), .A3(new_n387), .A4(G128), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n259), .B1(new_n385), .B2(KEYINPUT1), .ZN(new_n389));
  XNOR2_X1  g203(.A(G143), .B(G146), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n238), .ZN(new_n392));
  NAND2_X1  g206(.A1(KEYINPUT0), .A2(G128), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n385), .A2(new_n386), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n393), .ZN(new_n395));
  NOR2_X1   g209(.A1(KEYINPUT0), .A2(G128), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n394), .B1(new_n397), .B2(new_n390), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G125), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n392), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(G224), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n401), .A2(G953), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n402), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n392), .A2(new_n399), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT7), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n403), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n392), .A2(new_n399), .A3(new_n406), .A4(new_n404), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n362), .A2(new_n364), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n368), .A2(new_n369), .ZN(new_n412));
  INV_X1    g226(.A(new_n366), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(new_n372), .A3(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(G101), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  XOR2_X1   g230(.A(KEYINPUT80), .B(KEYINPUT4), .Z(new_n417));
  NAND2_X1  g231(.A1(new_n350), .A2(new_n353), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n379), .A2(KEYINPUT67), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n419), .A3(new_n351), .ZN(new_n420));
  INV_X1    g234(.A(new_n352), .ZN(new_n421));
  AOI22_X1  g235(.A1(new_n416), .A2(new_n417), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n415), .A2(KEYINPUT4), .A3(new_n373), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n422), .A2(new_n423), .B1(new_n359), .B2(new_n376), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n410), .B1(new_n424), .B2(new_n340), .ZN(new_n425));
  AOI21_X1  g239(.A(G902), .B1(new_n384), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n420), .A2(new_n421), .ZN(new_n427));
  OAI211_X1 g241(.A(G101), .B(new_n417), .C1(new_n411), .C2(new_n414), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n423), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n356), .A2(new_n358), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(new_n421), .A3(new_n376), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n340), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n429), .A2(new_n431), .A3(new_n340), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(KEYINPUT6), .A3(new_n435), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n403), .A2(new_n405), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT6), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n432), .A2(new_n438), .A3(new_n433), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n436), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n426), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G210), .B1(G237), .B2(G902), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT84), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n426), .A2(new_n440), .A3(new_n444), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n339), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G221), .ZN(new_n449));
  INV_X1    g263(.A(new_n294), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n449), .B1(new_n450), .B2(new_n187), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT82), .ZN(new_n452));
  NAND2_X1  g266(.A1(KEYINPUT65), .A2(G131), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G134), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G137), .ZN(new_n456));
  INV_X1    g270(.A(G137), .ZN(new_n457));
  AOI21_X1  g271(.A(KEYINPUT64), .B1(new_n457), .B2(G134), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT11), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n456), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT64), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n461), .B(new_n459), .C1(new_n455), .C2(G137), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n454), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n457), .A2(G134), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n461), .B1(new_n455), .B2(G137), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n465), .B1(new_n466), .B2(KEYINPUT11), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(new_n453), .A3(new_n462), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n391), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n378), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n385), .A2(new_n386), .ZN(new_n473));
  OAI211_X1 g287(.A(KEYINPUT81), .B(KEYINPUT1), .C1(new_n193), .C2(G146), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(G128), .ZN(new_n475));
  AOI21_X1  g289(.A(KEYINPUT81), .B1(new_n385), .B2(KEYINPUT1), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n388), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(new_n373), .A3(new_n375), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n470), .B1(new_n472), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n480), .A2(KEYINPUT12), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT12), .ZN(new_n482));
  AOI211_X1 g296(.A(new_n482), .B(new_n470), .C1(new_n472), .C2(new_n479), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n452), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n398), .A2(KEYINPUT68), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT68), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n394), .B(new_n486), .C1(new_n397), .C2(new_n390), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n423), .A2(new_n488), .A3(new_n428), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n376), .A2(KEYINPUT10), .A3(new_n391), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT10), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n479), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n489), .A2(new_n490), .A3(new_n470), .A4(new_n492), .ZN(new_n493));
  XNOR2_X1  g307(.A(G110), .B(G140), .ZN(new_n494));
  INV_X1    g308(.A(G227), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n495), .A2(G953), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n494), .B(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n479), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n391), .B1(new_n373), .B2(new_n375), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n469), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n482), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n480), .A2(KEYINPUT12), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT82), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n484), .A2(new_n499), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n489), .A2(new_n492), .A3(new_n490), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n469), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n493), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n497), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(G469), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n511), .A2(new_n512), .A3(new_n187), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n493), .B1(new_n481), .B2(new_n483), .ZN(new_n514));
  AOI22_X1  g328(.A1(new_n514), .A2(new_n497), .B1(new_n499), .B2(new_n508), .ZN(new_n515));
  OAI21_X1  g329(.A(G469), .B1(new_n515), .B2(G902), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n451), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n325), .A2(new_n448), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT95), .ZN(new_n519));
  NOR2_X1   g333(.A1(G472), .A2(G902), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT31), .ZN(new_n522));
  INV_X1    g336(.A(new_n487), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT0), .B(G128), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n473), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n486), .B1(new_n525), .B2(new_n394), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n460), .A2(new_n463), .A3(new_n454), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n453), .B1(new_n467), .B2(new_n462), .ZN(new_n528));
  OAI22_X1  g342(.A1(new_n523), .A2(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n387), .B1(G143), .B2(new_n227), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n473), .B1(new_n530), .B2(new_n259), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n457), .A2(G134), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n456), .ZN(new_n533));
  AOI22_X1  g347(.A1(new_n531), .A2(new_n388), .B1(G131), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n466), .A2(KEYINPUT11), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n535), .A2(new_n212), .A3(new_n462), .A4(new_n456), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n529), .A2(KEYINPUT30), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT30), .ZN(new_n539));
  AOI22_X1  g353(.A1(new_n464), .A2(new_n468), .B1(new_n525), .B2(new_n394), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n533), .A2(G131), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n391), .A2(new_n536), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n539), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n538), .A2(new_n427), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT69), .ZN(new_n545));
  AOI22_X1  g359(.A1(new_n488), .A2(new_n469), .B1(new_n536), .B2(new_n534), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n420), .A2(new_n421), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n538), .A2(new_n543), .A3(new_n545), .A4(new_n427), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n192), .A2(G210), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n552), .B1(new_n192), .B2(G210), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT26), .B(G101), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  OR3_X1    g370(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n556), .B1(new_n553), .B2(new_n554), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n522), .B1(new_n551), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n559), .ZN(new_n561));
  AOI211_X1 g375(.A(KEYINPUT31), .B(new_n561), .C1(new_n549), .C2(new_n550), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n540), .A2(new_n542), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n547), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n529), .A2(new_n420), .A3(new_n421), .A4(new_n537), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT28), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT28), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n546), .A2(new_n547), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n565), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  OR2_X1    g384(.A1(new_n570), .A2(new_n559), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n521), .B1(new_n563), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT72), .B1(new_n572), .B2(KEYINPUT32), .ZN(new_n573));
  INV_X1    g387(.A(G472), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT29), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n561), .B1(new_n570), .B2(new_n575), .ZN(new_n576));
  OR2_X1    g390(.A1(new_n546), .A2(new_n547), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n566), .A2(KEYINPUT28), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n568), .B1(new_n546), .B2(new_n547), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT29), .ZN(new_n581));
  AOI21_X1  g395(.A(G902), .B1(new_n576), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n559), .B1(new_n549), .B2(new_n550), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n575), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n574), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n585), .B1(new_n572), .B2(KEYINPUT32), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n551), .A2(new_n559), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT31), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n551), .A2(new_n522), .A3(new_n559), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n588), .A2(new_n571), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n520), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT72), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT32), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n573), .A2(new_n586), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n343), .A2(G128), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n259), .A2(G119), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(KEYINPUT74), .ZN(new_n599));
  XOR2_X1   g413(.A(KEYINPUT24), .B(G110), .Z(new_n600));
  NAND3_X1  g414(.A1(new_n259), .A2(KEYINPUT23), .A3(G119), .ZN(new_n601));
  INV_X1    g415(.A(new_n597), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n596), .B(new_n601), .C1(new_n602), .C2(KEYINPUT23), .ZN(new_n603));
  AOI22_X1  g417(.A1(new_n599), .A2(new_n600), .B1(G110), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n228), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n604), .B1(new_n309), .B2(new_n605), .ZN(new_n606));
  OAI22_X1  g420(.A1(new_n599), .A2(new_n600), .B1(G110), .B2(new_n603), .ZN(new_n607));
  OR2_X1    g421(.A1(new_n237), .A2(new_n240), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n607), .A2(new_n226), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT22), .B(G137), .ZN(new_n611));
  INV_X1    g425(.A(G234), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n449), .A2(new_n612), .A3(G953), .ZN(new_n613));
  XOR2_X1   g427(.A(new_n611), .B(new_n613), .Z(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n606), .A2(new_n609), .A3(new_n614), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n616), .A2(new_n187), .A3(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT25), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n616), .A2(KEYINPUT25), .A3(new_n187), .A4(new_n617), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(G217), .B1(new_n612), .B2(G902), .ZN(new_n623));
  XOR2_X1   g437(.A(new_n623), .B(KEYINPUT73), .Z(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n616), .A2(new_n617), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n623), .A2(new_n187), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(KEYINPUT77), .B1(new_n626), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n624), .B1(new_n620), .B2(new_n621), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT77), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n632), .A2(new_n629), .A3(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT95), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n325), .A2(new_n448), .A3(new_n517), .A4(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n519), .A2(new_n595), .A3(new_n635), .A4(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT96), .B(G101), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G3));
  NAND2_X1  g454(.A1(new_n590), .A2(new_n187), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n572), .B1(G472), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n642), .A2(new_n635), .A3(new_n517), .ZN(new_n643));
  XOR2_X1   g457(.A(new_n643), .B(KEYINPUT97), .Z(new_n644));
  NAND2_X1  g458(.A1(new_n319), .A2(new_n320), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(KEYINPUT20), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n319), .A2(new_n305), .A3(new_n320), .ZN(new_n647));
  AOI22_X1  g461(.A1(new_n646), .A2(new_n647), .B1(G475), .B2(new_n255), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n187), .A2(G478), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n293), .A2(new_n297), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n296), .B1(new_n299), .B2(new_n282), .ZN(new_n651));
  OAI21_X1  g465(.A(KEYINPUT33), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT33), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n298), .A2(new_n653), .A3(new_n300), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n649), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g469(.A(KEYINPUT98), .B1(new_n301), .B2(G478), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI211_X1 g471(.A(KEYINPUT98), .B(new_n649), .C1(new_n652), .C2(new_n654), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n648), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n426), .A2(new_n440), .A3(new_n442), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n442), .B1(new_n426), .B2(new_n440), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n339), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n644), .A2(new_n660), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT34), .B(G104), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G6));
  XOR2_X1   g482(.A(new_n301), .B(new_n303), .Z(new_n669));
  NAND4_X1  g483(.A1(new_n644), .A2(new_n669), .A3(new_n648), .A4(new_n665), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT35), .B(G107), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G9));
  NAND2_X1  g486(.A1(new_n641), .A2(G472), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n591), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n610), .B(KEYINPUT99), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n615), .A2(KEYINPUT36), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n626), .B1(new_n677), .B2(new_n628), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n519), .A2(new_n680), .A3(new_n637), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT37), .B(G110), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT100), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n681), .B(new_n683), .ZN(G12));
  INV_X1    g498(.A(new_n451), .ZN(new_n685));
  AOI211_X1 g499(.A(G469), .B(G902), .C1(new_n506), .C2(new_n510), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n514), .A2(new_n497), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n499), .A2(new_n508), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n512), .B1(new_n689), .B2(new_n187), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n685), .B1(new_n686), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n691), .A2(new_n679), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n595), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n336), .B1(new_n662), .B2(new_n663), .ZN(new_n694));
  OAI211_X1 g508(.A(new_n669), .B(new_n256), .C1(new_n321), .C2(new_n323), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n330), .B(KEYINPUT102), .Z(new_n696));
  NOR2_X1   g510(.A1(new_n203), .A2(G900), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n697), .A2(G902), .A3(new_n328), .ZN(new_n698));
  XOR2_X1   g512(.A(new_n698), .B(KEYINPUT101), .Z(new_n699));
  NAND2_X1  g513(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n694), .A2(new_n695), .A3(new_n701), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n693), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n259), .ZN(G30));
  NAND2_X1  g518(.A1(new_n446), .A2(new_n447), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT38), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n648), .A2(new_n304), .ZN(new_n707));
  AND4_X1   g521(.A1(new_n336), .A2(new_n706), .A3(new_n679), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n700), .B(KEYINPUT39), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n517), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(KEYINPUT40), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n710), .A2(KEYINPUT40), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n708), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT104), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n592), .B1(new_n591), .B2(new_n593), .ZN(new_n715));
  AOI211_X1 g529(.A(KEYINPUT72), .B(KEYINPUT32), .C1(new_n590), .C2(new_n520), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n559), .B1(new_n547), .B2(new_n546), .ZN(new_n718));
  AOI21_X1  g532(.A(G902), .B1(new_n718), .B2(new_n577), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n719), .B1(new_n551), .B2(new_n561), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(G472), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT103), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n720), .A2(KEYINPUT103), .A3(G472), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n725), .B1(KEYINPUT32), .B2(new_n572), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n714), .B1(new_n717), .B2(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n726), .A2(new_n714), .A3(new_n573), .A4(new_n594), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n713), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(new_n193), .ZN(G45));
  OAI21_X1  g546(.A(new_n256), .B1(new_n321), .B2(new_n323), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n657), .A2(new_n658), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n734), .A3(new_n700), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n694), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n693), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(new_n227), .ZN(G48));
  OR2_X1    g552(.A1(new_n631), .A2(new_n634), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n739), .B1(new_n717), .B2(new_n586), .ZN(new_n740));
  INV_X1    g554(.A(new_n511), .ZN(new_n741));
  OAI21_X1  g555(.A(G469), .B1(new_n741), .B2(G902), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n685), .A3(new_n513), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n744), .A2(new_n660), .A3(new_n665), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n740), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(KEYINPUT41), .B(G113), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G15));
  NOR4_X1   g562(.A1(new_n743), .A2(new_n664), .A3(new_n339), .A4(new_n695), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n740), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G116), .ZN(G18));
  NOR3_X1   g565(.A1(new_n743), .A2(new_n694), .A3(new_n679), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n752), .A2(new_n595), .A3(new_n325), .A4(new_n334), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G119), .ZN(G21));
  INV_X1    g568(.A(KEYINPUT105), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n673), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n641), .A2(KEYINPUT105), .A3(G472), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n580), .A2(new_n561), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n563), .A2(new_n758), .ZN(new_n759));
  AOI22_X1  g573(.A1(new_n756), .A2(new_n757), .B1(new_n520), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n626), .A2(new_n630), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n743), .A2(new_n694), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n648), .A2(new_n304), .A3(new_n335), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n760), .A2(new_n762), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G122), .ZN(G24));
  NAND2_X1  g580(.A1(new_n756), .A2(new_n757), .ZN(new_n767));
  INV_X1    g581(.A(new_n735), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n759), .A2(new_n520), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n752), .A2(new_n767), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G125), .ZN(G27));
  NAND3_X1  g585(.A1(new_n446), .A2(new_n447), .A3(new_n336), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n735), .A2(new_n691), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n591), .A2(new_n593), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n761), .B1(new_n586), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n773), .A2(new_n775), .A3(KEYINPUT42), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n773), .A2(new_n595), .A3(new_n635), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT42), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(KEYINPUT106), .A3(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT106), .B1(new_n777), .B2(new_n778), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n776), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G131), .ZN(G33));
  NOR2_X1   g597(.A1(new_n691), .A2(new_n772), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT107), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n648), .A2(new_n785), .A3(new_n669), .A4(new_n700), .ZN(new_n786));
  OAI21_X1  g600(.A(KEYINPUT107), .B1(new_n695), .B2(new_n701), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n784), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT108), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n740), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n595), .A2(new_n635), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n784), .A2(new_n786), .A3(new_n787), .ZN(new_n792));
  OAI21_X1  g606(.A(KEYINPUT108), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G134), .ZN(G36));
  NOR2_X1   g609(.A1(new_n659), .A2(new_n733), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT43), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(KEYINPUT43), .B1(new_n659), .B2(new_n733), .ZN(new_n799));
  AND4_X1   g613(.A1(new_n674), .A2(new_n798), .A3(new_n678), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(KEYINPUT44), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT109), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n800), .A2(KEYINPUT44), .ZN(new_n803));
  INV_X1    g617(.A(new_n772), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT45), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n512), .B1(new_n689), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n806), .B1(new_n805), .B2(new_n689), .ZN(new_n807));
  NAND2_X1  g621(.A1(G469), .A2(G902), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT46), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n686), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n807), .A2(KEYINPUT46), .A3(new_n808), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n451), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n813), .A2(new_n709), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n803), .A2(new_n804), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n802), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G137), .ZN(G39));
  NAND2_X1  g631(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n813), .A2(new_n818), .ZN(new_n819));
  XOR2_X1   g633(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n820));
  OAI21_X1  g634(.A(new_n819), .B1(new_n813), .B2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  NOR4_X1   g636(.A1(new_n595), .A2(new_n635), .A3(new_n735), .A4(new_n772), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(G140), .ZN(G42));
  AND2_X1   g639(.A1(new_n742), .A2(new_n513), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT49), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XOR2_X1   g642(.A(new_n828), .B(KEYINPUT111), .Z(new_n829));
  NOR2_X1   g643(.A1(new_n826), .A2(new_n827), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n796), .A2(new_n762), .A3(new_n685), .A4(new_n336), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n830), .A2(new_n831), .A3(new_n706), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n829), .A2(new_n832), .A3(new_n730), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n739), .A2(new_n691), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n695), .B1(new_n648), .B2(new_n659), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n835), .A2(new_n642), .A3(new_n448), .A4(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n638), .A2(new_n837), .A3(new_n681), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n772), .A2(new_n324), .A3(new_n701), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n595), .A2(new_n692), .A3(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT112), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n595), .A2(KEYINPUT112), .A3(new_n692), .A4(new_n839), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n838), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n595), .B(new_n692), .C1(new_n702), .C2(new_n736), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n770), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n694), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n678), .A2(new_n701), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n707), .A2(new_n847), .A3(new_n517), .A4(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n572), .A2(KEYINPUT32), .ZN(new_n850));
  INV_X1    g664(.A(new_n725), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n573), .A2(new_n594), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(KEYINPUT104), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n849), .B1(new_n853), .B2(new_n728), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT52), .B1(new_n846), .B2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n849), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n856), .B1(new_n727), .B2(new_n729), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT52), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n857), .A2(new_n858), .A3(new_n770), .A4(new_n845), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n760), .A2(new_n678), .ZN(new_n860));
  AOI22_X1  g674(.A1(new_n790), .A2(new_n793), .B1(new_n860), .B2(new_n773), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n844), .A2(new_n855), .A3(new_n859), .A4(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n740), .B1(new_n745), .B2(new_n749), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n863), .A2(new_n753), .A3(new_n765), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n782), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n834), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n859), .A2(new_n855), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n836), .A2(new_n448), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n643), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n426), .A2(new_n440), .A3(new_n444), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n444), .B1(new_n426), .B2(new_n440), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n338), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n873), .A2(new_n324), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n636), .B1(new_n874), .B2(new_n517), .ZN(new_n875));
  INV_X1    g689(.A(new_n637), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n870), .B1(new_n877), .B2(new_n740), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n842), .A2(new_n843), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n878), .A2(new_n879), .A3(new_n681), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n760), .A2(new_n678), .A3(new_n773), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n789), .B1(new_n740), .B2(new_n788), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n791), .A2(new_n792), .A3(KEYINPUT108), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n777), .A2(new_n778), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT106), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n779), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n864), .B1(new_n889), .B2(new_n776), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n868), .A2(new_n885), .A3(new_n890), .A4(KEYINPUT53), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n867), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT54), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n859), .A2(KEYINPUT53), .A3(new_n855), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT113), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n895), .B1(new_n880), .B2(new_n884), .ZN(new_n896));
  INV_X1    g710(.A(new_n838), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n861), .A2(KEYINPUT113), .A3(new_n897), .A4(new_n879), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n894), .A2(new_n896), .A3(new_n890), .A4(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT54), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n867), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n893), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n744), .A2(KEYINPUT117), .A3(new_n804), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT117), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n904), .B1(new_n743), .B2(new_n772), .ZN(new_n905));
  AOI211_X1 g719(.A(new_n739), .B(new_n330), .C1(new_n903), .C2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(new_n660), .A3(new_n730), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n903), .A2(new_n905), .ZN(new_n908));
  INV_X1    g722(.A(new_n696), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n798), .A2(new_n909), .A3(new_n799), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n908), .A2(new_n911), .A3(new_n775), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT121), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT48), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n907), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n913), .A2(KEYINPUT48), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n912), .A2(new_n916), .A3(new_n914), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n760), .A2(new_n762), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n918), .A2(new_n910), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n763), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n327), .B(KEYINPUT120), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n917), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n915), .A2(new_n922), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n860), .A2(new_n911), .A3(new_n908), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT116), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT50), .ZN(new_n926));
  INV_X1    g740(.A(new_n919), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n705), .B(KEYINPUT38), .Z(new_n928));
  NAND3_X1  g742(.A1(new_n928), .A2(new_n337), .A3(new_n744), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n925), .B(new_n926), .C1(new_n927), .C2(new_n929), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n929), .A2(new_n918), .A3(new_n910), .ZN(new_n931));
  OAI21_X1  g745(.A(KEYINPUT50), .B1(new_n931), .B2(KEYINPUT116), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n924), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n648), .A2(new_n659), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n906), .A2(new_n730), .A3(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT118), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n933), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n826), .A2(new_n451), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n821), .A2(KEYINPUT119), .A3(new_n940), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n918), .A2(new_n772), .A3(new_n910), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(KEYINPUT119), .B1(new_n821), .B2(new_n940), .ZN(new_n944));
  OAI21_X1  g758(.A(KEYINPUT51), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n923), .B1(new_n939), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT51), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n821), .A2(KEYINPUT114), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n940), .B(KEYINPUT115), .Z(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n821), .A2(KEYINPUT114), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n942), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n952), .A2(new_n933), .A3(new_n938), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n946), .B1(new_n947), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n902), .A2(KEYINPUT122), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n326), .A2(new_n203), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(KEYINPUT122), .B1(new_n902), .B2(new_n954), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n833), .B1(new_n957), .B2(new_n958), .ZN(G75));
  AOI21_X1  g773(.A(new_n187), .B1(new_n867), .B2(new_n899), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT56), .B1(new_n960), .B2(G210), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n436), .A2(new_n439), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(new_n437), .Z(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT55), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n961), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n203), .A2(G952), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  OR3_X1    g783(.A1(new_n961), .A2(KEYINPUT123), .A3(new_n965), .ZN(new_n970));
  OAI21_X1  g784(.A(KEYINPUT123), .B1(new_n961), .B2(new_n965), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(G51));
  AOI211_X1 g786(.A(new_n187), .B(new_n807), .C1(new_n867), .C2(new_n899), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n808), .B(KEYINPUT57), .Z(new_n974));
  AND3_X1   g788(.A1(new_n867), .A2(new_n899), .A3(new_n900), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n900), .B1(new_n867), .B2(new_n899), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n973), .B1(new_n977), .B2(new_n511), .ZN(new_n978));
  OAI21_X1  g792(.A(KEYINPUT124), .B1(new_n978), .B2(new_n967), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT124), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n867), .A2(new_n899), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(KEYINPUT54), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n901), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n741), .B1(new_n983), .B2(new_n974), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n980), .B(new_n968), .C1(new_n984), .C2(new_n973), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n979), .A2(new_n985), .ZN(G54));
  AND2_X1   g800(.A1(KEYINPUT58), .A2(G475), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n960), .A2(new_n319), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n319), .B1(new_n960), .B2(new_n987), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n988), .A2(new_n989), .A3(new_n967), .ZN(G60));
  NAND2_X1  g804(.A1(new_n652), .A2(new_n654), .ZN(new_n991));
  INV_X1    g805(.A(new_n902), .ZN(new_n992));
  NAND2_X1  g806(.A1(G478), .A2(G902), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT59), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n991), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n983), .A2(new_n991), .A3(new_n994), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n968), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n995), .A2(new_n997), .ZN(G63));
  XNOR2_X1  g812(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n295), .A2(new_n187), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n981), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(new_n627), .ZN(new_n1003));
  OAI211_X1 g817(.A(new_n1003), .B(new_n968), .C1(new_n677), .C2(new_n1002), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT61), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1004), .B(new_n1005), .ZN(G66));
  OAI21_X1  g820(.A(G953), .B1(new_n331), .B2(new_n401), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n864), .A2(new_n838), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1007), .B1(new_n1008), .B2(G953), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n962), .B1(G898), .B2(new_n203), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1009), .B(new_n1010), .ZN(G69));
  NAND2_X1  g825(.A1(new_n538), .A2(new_n543), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1012), .B(new_n313), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT62), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1014), .B1(new_n731), .B2(new_n846), .ZN(new_n1015));
  INV_X1    g829(.A(new_n846), .ZN(new_n1016));
  OAI211_X1 g830(.A(KEYINPUT62), .B(new_n1016), .C1(new_n713), .C2(new_n730), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  AOI22_X1  g832(.A1(new_n802), .A2(new_n815), .B1(new_n822), .B2(new_n823), .ZN(new_n1019));
  INV_X1    g833(.A(new_n710), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n740), .A2(new_n1020), .A3(new_n804), .A4(new_n836), .ZN(new_n1021));
  AND3_X1   g835(.A1(new_n1018), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n1013), .B1(new_n1022), .B2(G953), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n707), .A2(new_n847), .ZN(new_n1024));
  INV_X1    g838(.A(new_n1024), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n814), .A2(new_n775), .A3(new_n1025), .ZN(new_n1026));
  AND3_X1   g840(.A1(new_n1026), .A2(new_n794), .A3(new_n1016), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1019), .A2(new_n782), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n697), .B1(new_n1028), .B2(new_n203), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1023), .B1(new_n1029), .B2(new_n1013), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n203), .B1(G227), .B2(G900), .ZN(new_n1031));
  XOR2_X1   g845(.A(new_n1031), .B(KEYINPUT126), .Z(new_n1032));
  XNOR2_X1  g846(.A(new_n1030), .B(new_n1032), .ZN(G72));
  NAND2_X1  g847(.A1(G472), .A2(G902), .ZN(new_n1034));
  XOR2_X1   g848(.A(new_n1034), .B(KEYINPUT63), .Z(new_n1035));
  INV_X1    g849(.A(new_n1008), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1035), .B1(new_n1028), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n967), .B1(new_n1037), .B2(new_n583), .ZN(new_n1038));
  NOR2_X1   g852(.A1(new_n551), .A2(new_n561), .ZN(new_n1039));
  INV_X1    g853(.A(new_n1035), .ZN(new_n1040));
  NOR3_X1   g854(.A1(new_n1039), .A2(new_n583), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n892), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n1018), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1043));
  OAI21_X1  g857(.A(new_n1035), .B1(new_n1043), .B2(new_n1036), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1044), .A2(new_n1039), .ZN(new_n1045));
  NAND3_X1  g859(.A1(new_n1038), .A2(new_n1042), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g860(.A(KEYINPUT127), .ZN(new_n1047));
  XNOR2_X1  g861(.A(new_n1046), .B(new_n1047), .ZN(G57));
endmodule


