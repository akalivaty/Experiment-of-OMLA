//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  INV_X1    g0012(.A(KEYINPUT64), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n213), .B1(G1), .B2(G13), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(KEYINPUT64), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n207), .ZN(new_n218));
  INV_X1    g0018(.A(new_n201), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n212), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT65), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n209), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n230));
  OR2_X1    g0030(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n222), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT66), .Z(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G226), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT70), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT69), .B(G50), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XOR2_X1   g0049(.A(G107), .B(G116), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G33), .ZN(new_n256));
  AND2_X1   g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G232), .A3(G1698), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n257), .A2(G226), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G97), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G41), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n263), .B1(new_n214), .B2(new_n216), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n268));
  NAND2_X1  g0068(.A1(KEYINPUT72), .A2(G1), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(KEYINPUT72), .A2(G1), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G41), .A2(G45), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n268), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G238), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(KEYINPUT71), .A3(new_n206), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT71), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(new_n273), .B2(G1), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n263), .A2(G1), .A3(G13), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n277), .A2(new_n279), .A3(G274), .A4(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n276), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(KEYINPUT13), .B1(new_n267), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT13), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n266), .A2(new_n284), .A3(new_n281), .A4(new_n276), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G200), .ZN(new_n287));
  OR2_X1    g0087(.A1(KEYINPUT72), .A2(G1), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n288), .A2(G13), .A3(G20), .A4(new_n269), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n215), .A2(KEYINPUT64), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n213), .A2(G1), .A3(G13), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  NOR3_X1   g0095(.A1(new_n270), .A2(new_n271), .A3(new_n207), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n295), .A2(G68), .A3(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(G20), .A2(G33), .ZN(new_n299));
  INV_X1    g0099(.A(G68), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n299), .A2(G50), .B1(G20), .B2(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n253), .A2(G20), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n302), .B(KEYINPUT73), .ZN(new_n303));
  INV_X1    g0103(.A(G77), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n301), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n294), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT11), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n298), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(KEYINPUT11), .B1(new_n305), .B2(new_n294), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n289), .A2(G68), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT12), .ZN(new_n311));
  NOR3_X1   g0111(.A1(new_n308), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n283), .A2(G190), .A3(new_n285), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n287), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT14), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n286), .B2(G169), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n283), .A2(G179), .A3(new_n285), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n286), .A2(new_n316), .A3(G169), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n312), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n315), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT10), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT75), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G200), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n257), .A2(G222), .A3(new_n259), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n257), .A2(G223), .A3(G1698), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n328), .B(new_n329), .C1(new_n304), .C2(new_n257), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n265), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n275), .A2(G226), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n332), .A2(new_n281), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n327), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n331), .A2(new_n333), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n334), .B1(new_n336), .B2(G190), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n299), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT8), .B(G58), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n338), .B1(new_n303), .B2(new_n339), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n340), .A2(new_n294), .B1(new_n202), .B2(new_n290), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n295), .A2(G50), .A3(new_n297), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT9), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n337), .A2(new_n345), .ZN(new_n346));
  OAI22_X1  g0146(.A1(new_n343), .A2(new_n344), .B1(KEYINPUT75), .B2(new_n324), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n326), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n347), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n349), .A2(new_n337), .A3(new_n325), .A4(new_n345), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n335), .A2(G179), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT74), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT74), .ZN(new_n353));
  INV_X1    g0153(.A(G169), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n353), .B1(new_n335), .B2(new_n354), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n352), .B(new_n343), .C1(new_n351), .C2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n339), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n357), .A2(new_n299), .B1(G20), .B2(G77), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT15), .B(G87), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n302), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n362), .A2(new_n294), .B1(new_n304), .B2(new_n290), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n295), .A2(G77), .A3(new_n297), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n257), .A2(G232), .A3(new_n259), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n257), .A2(G238), .A3(G1698), .ZN(new_n367));
  INV_X1    g0167(.A(G107), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n366), .B(new_n367), .C1(new_n368), .C2(new_n257), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n265), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n275), .A2(G244), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n281), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n365), .B1(new_n373), .B2(G190), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(G200), .ZN(new_n375));
  INV_X1    g0175(.A(G179), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n372), .A2(new_n354), .B1(new_n364), .B2(new_n363), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n374), .A2(new_n375), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AND4_X1   g0179(.A1(new_n348), .A2(new_n350), .A3(new_n356), .A4(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n275), .A2(G232), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n381), .A2(new_n281), .ZN(new_n382));
  MUX2_X1   g0182(.A(G223), .B(G226), .S(G1698), .Z(new_n383));
  NAND2_X1  g0183(.A1(new_n255), .A2(KEYINPUT76), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT76), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT3), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(new_n386), .A3(G33), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n383), .A2(new_n387), .A3(new_n254), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT77), .ZN(new_n389));
  INV_X1    g0189(.A(G87), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n253), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n388), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n265), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n389), .B1(new_n388), .B2(new_n392), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n382), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G200), .ZN(new_n397));
  INV_X1    g0197(.A(G58), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n398), .A2(new_n300), .ZN(new_n399));
  OAI21_X1  g0199(.A(G20), .B1(new_n399), .B2(new_n201), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n299), .A2(G159), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n387), .A2(new_n254), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT7), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(new_n405), .A3(new_n207), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(G68), .ZN(new_n407));
  AOI21_X1  g0207(.A(G20), .B1(new_n387), .B2(new_n254), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n408), .A2(new_n405), .ZN(new_n409));
  OAI211_X1 g0209(.A(KEYINPUT16), .B(new_n403), .C1(new_n407), .C2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT16), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n405), .A2(G20), .ZN(new_n412));
  AOI21_X1  g0212(.A(G33), .B1(new_n384), .B2(new_n386), .ZN(new_n413));
  INV_X1    g0213(.A(new_n256), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n405), .B1(new_n257), .B2(G20), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n300), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n411), .B1(new_n417), .B2(new_n402), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n410), .A2(new_n418), .A3(new_n294), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n296), .A2(new_n339), .ZN(new_n420));
  AND3_X1   g0220(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n420), .A2(new_n421), .B1(new_n290), .B2(new_n339), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n382), .B(G190), .C1(new_n395), .C2(new_n394), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n397), .A2(new_n419), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT17), .ZN(new_n425));
  XNOR2_X1  g0225(.A(new_n424), .B(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n419), .A2(new_n422), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n382), .B(G179), .C1(new_n395), .C2(new_n394), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n381), .A2(new_n281), .ZN(new_n429));
  INV_X1    g0229(.A(new_n254), .ZN(new_n430));
  XNOR2_X1  g0230(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n430), .B1(new_n431), .B2(G33), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n391), .B1(new_n432), .B2(new_n383), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n264), .B1(new_n433), .B2(new_n389), .ZN(new_n434));
  INV_X1    g0234(.A(new_n395), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n429), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n428), .B1(new_n436), .B2(new_n354), .ZN(new_n437));
  AND3_X1   g0237(.A1(new_n427), .A2(KEYINPUT18), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT18), .B1(new_n427), .B2(new_n437), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n426), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n323), .A2(new_n380), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT78), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n323), .A2(new_n380), .A3(KEYINPUT78), .A4(new_n441), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AND2_X1   g0246(.A1(KEYINPUT5), .A2(G41), .ZN(new_n447));
  NOR2_X1   g0247(.A1(KEYINPUT5), .A2(G41), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G45), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n270), .A2(new_n271), .A3(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n450), .A2(new_n452), .A3(G274), .A4(new_n280), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n288), .A2(G45), .A3(new_n269), .ZN(new_n454));
  OAI211_X1 g0254(.A(G270), .B(new_n280), .C1(new_n454), .C2(new_n449), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  MUX2_X1   g0257(.A(G257), .B(G264), .S(G1698), .Z(new_n458));
  NAND3_X1  g0258(.A1(new_n458), .A2(new_n387), .A3(new_n254), .ZN(new_n459));
  INV_X1    g0259(.A(G303), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n460), .B1(new_n254), .B2(new_n256), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT82), .B1(new_n463), .B2(new_n265), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT82), .ZN(new_n465));
  AOI211_X1 g0265(.A(new_n465), .B(new_n264), .C1(new_n459), .C2(new_n462), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n457), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n289), .A2(G116), .ZN(new_n468));
  AOI21_X1  g0268(.A(G20), .B1(G33), .B2(G283), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n253), .A2(G97), .ZN(new_n470));
  INV_X1    g0270(.A(G116), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n469), .A2(new_n470), .B1(G20), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n294), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT20), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n472), .A2(new_n294), .A3(KEYINPUT20), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n468), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n288), .A2(KEYINPUT79), .A3(G33), .A4(new_n269), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n288), .A2(G33), .A3(new_n269), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT79), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n295), .A2(G116), .A3(new_n478), .A4(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n354), .B1(new_n477), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n467), .A2(KEYINPUT21), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n461), .B1(new_n432), .B2(new_n458), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n465), .B1(new_n485), .B2(new_n264), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n463), .A2(new_n265), .A3(KEYINPUT82), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n477), .A2(new_n482), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n488), .A2(new_n489), .A3(G179), .A4(new_n457), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n484), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT83), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT21), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n456), .B1(new_n486), .B2(new_n487), .ZN(new_n495));
  INV_X1    g0295(.A(new_n476), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT20), .B1(new_n472), .B2(new_n294), .ZN(new_n497));
  OAI22_X1  g0297(.A1(new_n496), .A2(new_n497), .B1(G116), .B2(new_n289), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n481), .A2(new_n421), .A3(new_n289), .A4(new_n478), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n499), .A2(new_n471), .ZN(new_n500));
  OAI21_X1  g0300(.A(G169), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n494), .B1(new_n495), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT84), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n467), .A2(new_n483), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(KEYINPUT84), .A3(new_n494), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n484), .A2(KEYINPUT83), .A3(new_n490), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n489), .B1(new_n467), .B2(G200), .ZN(new_n509));
  INV_X1    g0309(.A(G190), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n509), .B1(new_n510), .B2(new_n467), .ZN(new_n511));
  AND4_X1   g0311(.A1(new_n493), .A2(new_n507), .A3(new_n508), .A4(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n432), .A2(KEYINPUT22), .A3(new_n207), .A4(G87), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT22), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n254), .A2(new_n256), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n207), .A2(G87), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT23), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n207), .B2(G107), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n368), .A2(KEYINPUT23), .A3(G20), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n519), .A2(new_n520), .B1(new_n302), .B2(G116), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n513), .A2(new_n517), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT24), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT24), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n513), .A2(new_n517), .A3(new_n524), .A4(new_n521), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n421), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n368), .B1(KEYINPUT85), .B2(KEYINPUT25), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n289), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n529));
  XOR2_X1   g0329(.A(new_n528), .B(new_n529), .Z(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n368), .B2(new_n499), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  AND2_X1   g0333(.A1(G257), .A2(G1698), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n387), .A2(KEYINPUT86), .A3(new_n254), .A4(new_n534), .ZN(new_n535));
  XNOR2_X1  g0335(.A(KEYINPUT87), .B(G294), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G33), .ZN(new_n537));
  INV_X1    g0337(.A(G250), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n538), .A2(G1698), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n387), .A2(new_n254), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n535), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT86), .B1(new_n432), .B2(new_n534), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n265), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(G264), .B(new_n280), .C1(new_n454), .C2(new_n449), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT88), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT88), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n543), .A2(new_n547), .A3(new_n544), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n453), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n327), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n543), .A2(new_n510), .A3(new_n453), .A4(new_n544), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n533), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n546), .A2(G179), .A3(new_n453), .A4(new_n548), .ZN(new_n553));
  INV_X1    g0353(.A(new_n453), .ZN(new_n554));
  OAI21_X1  g0354(.A(G169), .B1(new_n545), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n532), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G116), .ZN(new_n558));
  OR2_X1    g0358(.A1(G238), .A2(G1698), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(G244), .B2(new_n259), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n558), .B1(new_n404), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n265), .ZN(new_n562));
  INV_X1    g0362(.A(G274), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n288), .A2(G45), .A3(new_n563), .A4(new_n269), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n280), .B(new_n564), .C1(new_n452), .C2(G250), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT80), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n268), .B1(new_n454), .B2(new_n538), .ZN(new_n568));
  AOI21_X1  g0368(.A(KEYINPUT80), .B1(new_n568), .B2(new_n564), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n562), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n570), .A2(KEYINPUT81), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT81), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n565), .A2(new_n566), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n568), .A2(KEYINPUT80), .A3(new_n564), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n572), .B1(new_n575), .B2(new_n562), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n354), .B1(new_n571), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n570), .A2(KEYINPUT81), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n575), .A2(new_n572), .A3(new_n562), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n578), .A2(new_n376), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n432), .A2(new_n207), .A3(G68), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT19), .B1(new_n302), .B2(G97), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT19), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n207), .B1(new_n261), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(G97), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n390), .A2(new_n585), .A3(new_n368), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n582), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n588), .A2(new_n294), .B1(new_n290), .B2(new_n359), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(new_n359), .B2(new_n499), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n577), .A2(new_n580), .A3(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(G200), .B1(new_n571), .B2(new_n576), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n578), .A2(G190), .A3(new_n579), .ZN(new_n593));
  OR2_X1    g0393(.A1(new_n499), .A2(new_n390), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n368), .B1(new_n415), .B2(new_n416), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n299), .A2(G77), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT6), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n599), .A2(new_n585), .A3(G107), .ZN(new_n600));
  XNOR2_X1  g0400(.A(G97), .B(G107), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n600), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n598), .B1(new_n602), .B2(new_n207), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n294), .B1(new_n597), .B2(new_n603), .ZN(new_n604));
  MUX2_X1   g0404(.A(new_n289), .B(new_n499), .S(G97), .Z(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI211_X1 g0406(.A(G257), .B(new_n280), .C1(new_n454), .C2(new_n449), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n453), .A2(new_n607), .ZN(new_n608));
  AND2_X1   g0408(.A1(KEYINPUT4), .A2(G244), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n254), .A2(new_n256), .A3(new_n609), .A4(new_n259), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n254), .A2(new_n256), .A3(G250), .A4(G1698), .ZN(new_n611));
  NAND2_X1  g0411(.A1(G33), .A2(G283), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT4), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n387), .A2(G244), .A3(new_n259), .A4(new_n254), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n608), .B(new_n376), .C1(new_n616), .C2(new_n264), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n614), .ZN(new_n618));
  INV_X1    g0418(.A(new_n613), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n264), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n453), .A2(new_n607), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n354), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n606), .A2(new_n617), .A3(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(G200), .B1(new_n620), .B2(new_n621), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n608), .B(G190), .C1(new_n616), .C2(new_n264), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n624), .A2(new_n625), .A3(new_n604), .A4(new_n605), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n591), .A2(new_n596), .A3(new_n627), .ZN(new_n628));
  AND4_X1   g0428(.A1(new_n446), .A2(new_n512), .A3(new_n557), .A4(new_n628), .ZN(G372));
  AND2_X1   g0429(.A1(new_n484), .A2(new_n490), .ZN(new_n630));
  AOI21_X1  g0430(.A(KEYINPUT84), .B1(new_n505), .B2(new_n494), .ZN(new_n631));
  AOI211_X1 g0431(.A(new_n503), .B(KEYINPUT21), .C1(new_n467), .C2(new_n483), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT89), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n553), .A2(new_n555), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n533), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n507), .A2(KEYINPUT89), .A3(new_n630), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n635), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n570), .A2(new_n354), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n580), .A2(new_n590), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n570), .A2(G200), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n593), .A2(new_n595), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n627), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n552), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n641), .ZN(new_n647));
  INV_X1    g0447(.A(new_n623), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n641), .A2(new_n643), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g0451(.A(KEYINPUT90), .B(KEYINPUT26), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n591), .A2(new_n596), .A3(new_n648), .A4(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n647), .B1(new_n651), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n646), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n446), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n320), .A2(new_n319), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n322), .B1(new_n658), .B2(new_n317), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n377), .A2(new_n378), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n314), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n426), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT18), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT91), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n427), .A2(new_n665), .A3(new_n437), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n665), .B1(new_n427), .B2(new_n437), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n664), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n427), .A2(new_n437), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT91), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n427), .A2(new_n437), .A3(new_n665), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(KEYINPUT18), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n348), .B(new_n350), .C1(new_n663), .C2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n356), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n657), .A2(new_n677), .ZN(G369));
  INV_X1    g0478(.A(G330), .ZN(new_n679));
  INV_X1    g0479(.A(new_n489), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n207), .A2(G13), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n272), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT92), .ZN(new_n684));
  INV_X1    g0484(.A(G213), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n685), .B1(new_n682), .B2(KEYINPUT27), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(G343), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n512), .B1(new_n680), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n635), .A2(new_n638), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n689), .A2(new_n680), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n679), .B1(new_n690), .B2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n532), .A2(new_n689), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT93), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n557), .ZN(new_n698));
  INV_X1    g0498(.A(new_n689), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n556), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n694), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n556), .A2(new_n689), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n507), .A2(new_n493), .A3(new_n508), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n689), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n698), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n702), .A2(new_n703), .A3(new_n706), .ZN(G399));
  INV_X1    g0507(.A(new_n210), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G41), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n586), .A2(G116), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(G1), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n220), .B2(new_n710), .ZN(new_n713));
  XOR2_X1   g0513(.A(KEYINPUT94), .B(KEYINPUT28), .Z(new_n714));
  XNOR2_X1  g0514(.A(new_n713), .B(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT29), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n656), .A2(new_n716), .A3(new_n689), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n512), .A2(new_n557), .A3(new_n628), .A4(new_n689), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  AOI211_X1 g0519(.A(new_n376), .B(new_n456), .C1(new_n486), .C2(new_n487), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n608), .B1(new_n616), .B2(new_n264), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n720), .A2(new_n578), .A3(new_n579), .A4(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n546), .A2(new_n548), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n719), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n571), .A2(new_n576), .A3(new_n721), .ZN(new_n726));
  INV_X1    g0526(.A(new_n548), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n547), .B1(new_n543), .B2(new_n544), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n726), .A2(new_n729), .A3(KEYINPUT30), .A4(new_n720), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n721), .A2(new_n570), .A3(new_n376), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n549), .A2(new_n467), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n725), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n699), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT31), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n733), .A2(KEYINPUT31), .A3(new_n699), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n718), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G330), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n637), .A2(new_n493), .A3(new_n507), .A4(new_n508), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n647), .B1(new_n645), .B2(new_n740), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n641), .A2(new_n643), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT95), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n742), .A2(new_n743), .A3(KEYINPUT26), .A4(new_n648), .ZN(new_n744));
  OAI21_X1  g0544(.A(KEYINPUT95), .B1(new_n649), .B2(new_n650), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n591), .A2(new_n596), .A3(new_n648), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(new_n652), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n744), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n699), .B1(new_n741), .B2(new_n748), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n717), .B(new_n739), .C1(new_n716), .C2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n715), .B1(new_n751), .B2(G1), .ZN(G364));
  INV_X1    g0552(.A(new_n694), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n690), .A2(new_n693), .A3(new_n679), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n206), .B1(new_n681), .B2(G45), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n709), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n753), .A2(new_n754), .A3(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G13), .A2(G33), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n690), .A2(new_n693), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G179), .A2(G200), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n207), .B1(new_n764), .B2(G190), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n765), .A2(KEYINPUT99), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(KEYINPUT99), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n585), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G190), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n510), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n772), .A2(G68), .B1(new_n773), .B2(G50), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n207), .A2(G190), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(new_n764), .ZN(new_n776));
  INV_X1    g0576(.A(G159), .ZN(new_n777));
  OAI21_X1  g0577(.A(KEYINPUT32), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OR3_X1    g0578(.A1(new_n776), .A2(KEYINPUT32), .A3(new_n777), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n770), .A2(new_n774), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n376), .A2(G200), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT98), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n781), .B(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n775), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n368), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n783), .A2(new_n207), .A3(new_n510), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n390), .ZN(new_n790));
  NOR4_X1   g0590(.A1(new_n207), .A2(new_n376), .A3(G190), .A4(G200), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR4_X1   g0592(.A1(new_n207), .A2(new_n376), .A3(new_n510), .A4(G200), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n257), .B1(new_n792), .B2(new_n304), .C1(new_n794), .C2(new_n398), .ZN(new_n795));
  NOR4_X1   g0595(.A1(new_n780), .A2(new_n787), .A3(new_n790), .A4(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n536), .ZN(new_n797));
  INV_X1    g0597(.A(new_n773), .ZN(new_n798));
  INV_X1    g0598(.A(G326), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n768), .A2(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT100), .ZN(new_n801));
  INV_X1    g0601(.A(new_n776), .ZN(new_n802));
  AOI22_X1  g0602(.A1(G329), .A2(new_n802), .B1(new_n793), .B2(G322), .ZN(new_n803));
  INV_X1    g0603(.A(G311), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n803), .B(new_n515), .C1(new_n804), .C2(new_n792), .ZN(new_n805));
  INV_X1    g0605(.A(G283), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n789), .A2(new_n460), .B1(new_n786), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(KEYINPUT33), .B(G317), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n805), .B(new_n807), .C1(new_n772), .C2(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n796), .B1(new_n801), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n217), .B1(G20), .B2(new_n354), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n757), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n811), .A2(new_n762), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT97), .Z(new_n815));
  NOR2_X1   g0615(.A1(new_n708), .A2(new_n515), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(G355), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(G116), .B2(new_n210), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n248), .A2(G45), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n432), .B(new_n708), .C1(new_n451), .C2(new_n221), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n818), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n815), .B1(new_n821), .B2(KEYINPUT96), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(KEYINPUT96), .B2(new_n821), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n813), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n763), .A2(new_n824), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n759), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(G396));
  NAND2_X1  g0627(.A1(new_n656), .A2(new_n689), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n699), .A2(new_n365), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n374), .A2(new_n375), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n661), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n699), .A2(new_n660), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n828), .B(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n757), .B1(new_n834), .B2(new_n739), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n739), .B2(new_n834), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n811), .A2(new_n760), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n758), .B1(new_n837), .B2(new_n304), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n789), .A2(new_n368), .B1(new_n786), .B2(new_n390), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n802), .A2(G311), .B1(new_n791), .B2(G116), .ZN(new_n840));
  INV_X1    g0640(.A(G294), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n840), .B(new_n515), .C1(new_n841), .C2(new_n794), .ZN(new_n842));
  INV_X1    g0642(.A(new_n772), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n843), .A2(new_n806), .B1(new_n798), .B2(new_n460), .ZN(new_n844));
  NOR4_X1   g0644(.A1(new_n839), .A2(new_n842), .A3(new_n844), .A4(new_n769), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n793), .A2(G143), .B1(new_n791), .B2(G159), .ZN(new_n846));
  INV_X1    g0646(.A(G150), .ZN(new_n847));
  INV_X1    g0647(.A(G137), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n846), .B1(new_n843), .B2(new_n847), .C1(new_n848), .C2(new_n798), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT34), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n849), .A2(new_n850), .ZN(new_n852));
  INV_X1    g0652(.A(G132), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n432), .B1(new_n853), .B2(new_n776), .C1(new_n768), .C2(new_n398), .ZN(new_n854));
  NOR3_X1   g0654(.A1(new_n851), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n785), .A2(G68), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n789), .B2(new_n202), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT101), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n845), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n833), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n838), .B1(new_n812), .B2(new_n859), .C1(new_n860), .C2(new_n761), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n836), .A2(new_n861), .ZN(G384));
  INV_X1    g0662(.A(new_n602), .ZN(new_n863));
  OR2_X1    g0663(.A1(new_n863), .A2(KEYINPUT35), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(KEYINPUT35), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n864), .A2(G116), .A3(new_n218), .A4(new_n865), .ZN(new_n866));
  XOR2_X1   g0666(.A(new_n866), .B(KEYINPUT36), .Z(new_n867));
  OR3_X1    g0667(.A1(new_n220), .A2(new_n304), .A3(new_n399), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n202), .A2(G68), .ZN(new_n869));
  AOI211_X1 g0669(.A(G13), .B(new_n272), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n272), .A2(new_n681), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n410), .A2(new_n294), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n300), .B1(new_n408), .B2(new_n405), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT7), .B1(new_n432), .B2(G20), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n402), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n876), .A2(KEYINPUT16), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n422), .B1(new_n873), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n688), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(new_n426), .B2(new_n440), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n879), .A2(new_n424), .ZN(new_n882));
  INV_X1    g0682(.A(new_n437), .ZN(new_n883));
  INV_X1    g0683(.A(new_n422), .ZN(new_n884));
  OR2_X1    g0684(.A1(new_n876), .A2(KEYINPUT16), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n421), .B1(new_n876), .B2(KEYINPUT16), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT37), .B1(new_n882), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT37), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n424), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n427), .B1(new_n437), .B2(new_n688), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n881), .A2(new_n894), .A3(KEYINPUT38), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n427), .A2(new_n688), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n424), .B(KEYINPUT17), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n896), .B1(new_n673), .B2(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(KEYINPUT102), .B(new_n424), .C1(new_n666), .C2(new_n667), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n896), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n670), .A2(new_n671), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT102), .B1(new_n901), .B2(new_n424), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT37), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n898), .B1(new_n903), .B2(new_n893), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n895), .B1(new_n904), .B2(KEYINPUT38), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n659), .B(new_n314), .C1(new_n312), .C2(new_n689), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n322), .B(new_n699), .C1(new_n321), .C2(new_n315), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n833), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n738), .A2(new_n908), .A3(KEYINPUT40), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n905), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT38), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n669), .A2(new_n664), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n427), .A2(new_n437), .A3(KEYINPUT18), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n879), .B1(new_n897), .B2(new_n915), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n879), .B(new_n424), .C1(new_n883), .C2(new_n887), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n917), .A2(KEYINPUT37), .B1(new_n891), .B2(new_n892), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n912), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n895), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n920), .A2(new_n738), .A3(new_n908), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT40), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n911), .A2(new_n923), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n446), .A2(new_n738), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n926), .A2(new_n927), .A3(new_n679), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n920), .A2(KEYINPUT39), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n903), .A2(new_n893), .ZN(new_n930));
  INV_X1    g0730(.A(new_n898), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT38), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT39), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n895), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n929), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n321), .A2(new_n322), .A3(new_n689), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n906), .A2(new_n907), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n656), .A2(new_n689), .A3(new_n860), .ZN(new_n941));
  INV_X1    g0741(.A(new_n832), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n943), .A2(new_n920), .B1(new_n674), .B2(new_n687), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n938), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n717), .B1(new_n716), .B2(new_n749), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n676), .B1(new_n946), .B2(new_n446), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n945), .B(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n872), .B1(new_n928), .B2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT103), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n949), .A2(new_n950), .B1(new_n948), .B2(new_n928), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n949), .A2(new_n950), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n871), .B1(new_n951), .B2(new_n952), .ZN(G367));
  OAI21_X1  g0753(.A(new_n814), .B1(new_n210), .B2(new_n359), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n708), .A2(new_n432), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n954), .B1(new_n242), .B2(new_n955), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n257), .B1(new_n776), .B2(new_n848), .C1(new_n794), .C2(new_n847), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(G143), .B2(new_n773), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n791), .A2(G50), .B1(G159), .B2(new_n772), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT109), .ZN(new_n960));
  INV_X1    g0760(.A(new_n768), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(G68), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n788), .A2(G58), .B1(new_n785), .B2(G77), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n958), .A2(new_n960), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n785), .A2(G97), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n802), .A2(G317), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n793), .A2(G303), .B1(new_n791), .B2(G283), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n404), .B1(new_n798), .B2(new_n804), .C1(new_n797), .C2(new_n843), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n789), .A2(new_n471), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n970), .B1(KEYINPUT46), .B2(new_n971), .C1(new_n368), .C2(new_n768), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n788), .A2(KEYINPUT46), .A3(G116), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT108), .Z(new_n974));
  OAI21_X1  g0774(.A(new_n964), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT47), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n758), .B(new_n956), .C1(new_n976), .C2(new_n811), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n689), .A2(new_n595), .ZN(new_n978));
  MUX2_X1   g0778(.A(new_n742), .B(new_n647), .S(new_n978), .Z(new_n979));
  INV_X1    g0779(.A(new_n762), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n699), .A2(new_n606), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n627), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n699), .A2(new_n648), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n703), .B(new_n986), .C1(new_n698), .C2(new_n705), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT45), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n987), .B(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n703), .B1(new_n698), .B2(new_n705), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT105), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT44), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n986), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n991), .A2(new_n992), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n994), .A2(new_n995), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n989), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n702), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n989), .A2(new_n996), .A3(new_n702), .A4(new_n997), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n698), .A2(new_n700), .A3(new_n705), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1003), .A2(KEYINPUT106), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(KEYINPUT106), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1004), .A2(new_n706), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n694), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1004), .A2(new_n753), .A3(new_n706), .A4(new_n1005), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n751), .ZN(new_n1010));
  OAI21_X1  g0810(.A(KEYINPUT107), .B1(new_n1002), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n750), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT107), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1012), .A2(new_n1000), .A3(new_n1013), .A4(new_n1001), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n751), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n709), .B(KEYINPUT41), .Z(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n756), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n986), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n706), .A2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT42), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n623), .B1(new_n984), .B2(new_n637), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n689), .ZN(new_n1024));
  AND2_X1   g0824(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n979), .B(KEYINPUT43), .ZN(new_n1026));
  OAI21_X1  g0826(.A(KEYINPUT104), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n979), .A2(KEYINPUT43), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1026), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT104), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1027), .A2(new_n1029), .A3(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n702), .A2(new_n1020), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1027), .A2(new_n1034), .A3(new_n1029), .A4(new_n1032), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n982), .B1(new_n1019), .B2(new_n1038), .ZN(G387));
  OAI21_X1  g0839(.A(new_n404), .B1(new_n799), .B2(new_n776), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n793), .A2(G317), .B1(new_n791), .B2(G303), .ZN(new_n1041));
  INV_X1    g0841(.A(G322), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1041), .B1(new_n843), .B2(new_n804), .C1(new_n1042), .C2(new_n798), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT48), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n806), .B2(new_n768), .C1(new_n797), .C2(new_n789), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT49), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n1040), .B(new_n1049), .C1(G116), .C2(new_n785), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n788), .A2(G77), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n404), .B1(G150), .B2(new_n802), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1051), .A2(new_n965), .A3(new_n1052), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT110), .Z(new_n1054));
  NOR2_X1   g0854(.A1(new_n768), .A2(new_n359), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n793), .A2(G50), .B1(new_n791), .B2(G68), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1056), .B1(new_n843), .B2(new_n339), .C1(new_n777), .C2(new_n798), .ZN(new_n1057));
  NOR3_X1   g0857(.A1(new_n1054), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n811), .B1(new_n1050), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n711), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n816), .A2(new_n1060), .B1(new_n368), .B2(new_n708), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n238), .A2(G45), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n357), .A2(new_n202), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT50), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n711), .B(new_n451), .C1(new_n300), .C2(new_n304), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n955), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1061), .B1(new_n1062), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n758), .B1(new_n1067), .B2(new_n815), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1059), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n701), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1069), .B1(new_n1070), .B2(new_n762), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n1009), .B2(new_n756), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1010), .A2(new_n709), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1009), .A2(new_n751), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1072), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT111), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g0877(.A(KEYINPUT111), .B(new_n1072), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(G393));
  OAI21_X1  g0879(.A(new_n814), .B1(new_n585), .B2(new_n210), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n251), .B2(new_n955), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n515), .B1(new_n1042), .B2(new_n776), .C1(new_n792), .C2(new_n841), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n789), .A2(new_n806), .B1(new_n786), .B2(new_n368), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1082), .B(new_n1083), .C1(G303), .C2(new_n772), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n793), .A2(G311), .B1(G317), .B2(new_n773), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT52), .Z(new_n1086));
  OAI211_X1 g0886(.A(new_n1084), .B(new_n1086), .C1(new_n471), .C2(new_n768), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT114), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n788), .A2(G68), .B1(G143), .B2(new_n802), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT113), .Z(new_n1091));
  OAI221_X1 g0891(.A(new_n432), .B1(new_n843), .B2(new_n202), .C1(new_n792), .C2(new_n339), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n768), .A2(new_n304), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1092), .B(new_n1093), .C1(G87), .C2(new_n785), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n793), .A2(G159), .B1(G150), .B2(new_n773), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1095), .B(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1091), .A2(new_n1094), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1089), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n758), .B(new_n1081), .C1(new_n1100), .C2(new_n811), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n980), .B2(new_n986), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n1002), .B2(new_n755), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n710), .B1(new_n1002), .B2(new_n1010), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1103), .B1(new_n1015), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(G390));
  AND3_X1   g0906(.A1(new_n733), .A2(KEYINPUT31), .A3(new_n699), .ZN(new_n1107));
  AOI21_X1  g0907(.A(KEYINPUT31), .B1(new_n733), .B2(new_n699), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n679), .B1(new_n1109), .B2(new_n718), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n446), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(KEYINPUT115), .B1(new_n947), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n741), .A2(new_n748), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n716), .B1(new_n1113), .B2(new_n689), .ZN(new_n1114));
  AOI211_X1 g0914(.A(KEYINPUT29), .B(new_n699), .C1(new_n646), .C2(new_n655), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n446), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1116), .A2(KEYINPUT115), .A3(new_n677), .A4(new_n1111), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1112), .A2(new_n1118), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n699), .B(new_n831), .C1(new_n741), .C2(new_n748), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n939), .B1(new_n1120), .B2(new_n832), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1121), .A2(new_n905), .A3(new_n936), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n941), .A2(new_n942), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n937), .B1(new_n1123), .B2(new_n939), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1122), .B1(new_n1124), .B2(new_n935), .ZN(new_n1125));
  AND4_X1   g0925(.A1(G330), .A2(new_n738), .A3(new_n860), .A4(new_n939), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n933), .B(new_n895), .C1(new_n904), .C2(KEYINPUT38), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1128), .B(new_n929), .C1(new_n943), .C2(new_n937), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1110), .A2(new_n860), .A3(new_n939), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1129), .A2(new_n1130), .A3(new_n1122), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n939), .B1(new_n1110), .B2(new_n860), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1123), .B1(new_n1132), .B2(new_n1126), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n940), .B1(new_n739), .B2(new_n833), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1120), .A2(new_n832), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1134), .A2(new_n1135), .A3(new_n1130), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1119), .A2(new_n1127), .A3(new_n1131), .A4(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1116), .A2(new_n677), .A3(new_n1111), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT115), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1141), .A2(new_n1137), .A3(new_n1117), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n1129), .A2(new_n1130), .A3(new_n1122), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1130), .B1(new_n1129), .B2(new_n1122), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1138), .A2(new_n709), .A3(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1127), .A2(new_n756), .A3(new_n1131), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT116), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1128), .A2(new_n760), .A3(new_n929), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n772), .A2(G137), .B1(new_n773), .B2(G128), .ZN(new_n1150));
  XOR2_X1   g0950(.A(KEYINPUT54), .B(G143), .Z(new_n1151));
  AOI21_X1  g0951(.A(new_n515), .B1(new_n791), .B2(new_n1151), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(G125), .A2(new_n802), .B1(new_n793), .B2(G132), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n1150), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n1154), .B1(new_n202), .B2(new_n786), .C1(new_n777), .C2(new_n768), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n788), .A2(G150), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT53), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n794), .A2(new_n471), .B1(new_n776), .B2(new_n841), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n515), .B1(new_n792), .B2(new_n585), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n843), .A2(new_n368), .B1(new_n798), .B2(new_n806), .ZN(new_n1160));
  NOR3_X1   g0960(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1161), .B(new_n856), .C1(new_n390), .C2(new_n789), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n1155), .A2(new_n1157), .B1(new_n1162), .B2(new_n1093), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n811), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n758), .B1(new_n837), .B2(new_n339), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1149), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n1147), .A2(new_n1148), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1148), .B1(new_n1147), .B2(new_n1166), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1146), .B1(new_n1167), .B2(new_n1168), .ZN(G378));
  XOR2_X1   g0969(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n348), .A2(new_n350), .A3(new_n356), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n688), .A2(new_n343), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT119), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1176), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1171), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(KEYINPUT119), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1182), .A2(new_n1170), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1180), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n760), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n837), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n757), .B1(new_n1187), .B2(G50), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n793), .A2(G128), .B1(new_n791), .B2(G137), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n843), .B2(new_n853), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n788), .B2(new_n1151), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n961), .A2(G150), .B1(G125), .B2(new_n773), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT118), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1191), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  OR2_X1    g0996(.A1(new_n1196), .A2(KEYINPUT59), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(KEYINPUT59), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n785), .A2(G159), .ZN(new_n1199));
  AOI211_X1 g0999(.A(G33), .B(G41), .C1(new_n802), .C2(G124), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n431), .A2(new_n253), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n202), .B1(new_n1202), .B2(G41), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n432), .B1(new_n772), .B2(G97), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n962), .B(new_n1204), .C1(new_n471), .C2(new_n798), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n786), .A2(new_n398), .ZN(new_n1206));
  AOI21_X1  g1006(.A(G41), .B1(new_n360), .B2(new_n791), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(G283), .A2(new_n802), .B1(new_n793), .B2(G107), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1051), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(new_n1205), .A2(new_n1206), .A3(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1203), .B1(new_n1210), .B2(KEYINPUT58), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n1211), .A2(KEYINPUT117), .B1(KEYINPUT58), .B2(new_n1210), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1201), .B(new_n1212), .C1(KEYINPUT117), .C2(new_n1211), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1188), .B1(new_n1213), .B2(new_n811), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1186), .A2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n679), .B1(new_n921), .B2(new_n922), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n911), .A2(new_n1216), .A3(new_n1185), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1185), .B1(new_n911), .B2(new_n1216), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n945), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1180), .A2(new_n1184), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n923), .A2(G330), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n893), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n424), .B1(new_n666), .B2(new_n667), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT102), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1225), .A2(new_n896), .A3(new_n899), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1222), .B1(new_n1226), .B2(KEYINPUT37), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n912), .B1(new_n1227), .B2(new_n898), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n909), .B1(new_n1228), .B2(new_n895), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1220), .B1(new_n1221), .B2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n911), .A2(new_n1185), .A3(new_n1216), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1230), .A2(new_n938), .A3(new_n944), .A4(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1219), .A2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1215), .B1(new_n1233), .B2(new_n755), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT57), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1141), .A2(new_n1117), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1236), .B1(new_n1237), .B2(new_n1137), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1235), .B1(new_n1238), .B2(new_n1233), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1127), .A2(new_n1131), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1119), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1219), .A2(new_n1232), .A3(KEYINPUT57), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n710), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1234), .B1(new_n1239), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(G375));
  NOR2_X1   g1046(.A1(new_n939), .A2(new_n761), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT121), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n789), .A2(new_n585), .B1(new_n786), .B2(new_n304), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(G303), .A2(new_n802), .B1(new_n793), .B2(G283), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n257), .B1(G107), .B2(new_n791), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n772), .A2(G116), .B1(new_n773), .B2(G294), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1250), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1249), .A2(new_n1253), .A3(new_n1055), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(G128), .A2(new_n802), .B1(new_n793), .B2(G137), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n1151), .A2(new_n772), .B1(G132), .B2(new_n773), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1255), .A2(new_n432), .A3(new_n1256), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n1257), .B(new_n1206), .C1(G159), .C2(new_n788), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n768), .A2(new_n202), .B1(new_n847), .B2(new_n792), .ZN(new_n1259));
  XOR2_X1   g1059(.A(new_n1259), .B(KEYINPUT122), .Z(new_n1260));
  AOI21_X1  g1060(.A(new_n1254), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1261));
  OAI221_X1 g1061(.A(new_n757), .B1(G68), .B2(new_n1187), .C1(new_n1261), .C2(new_n812), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1248), .A2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(new_n1137), .B2(new_n756), .ZN(new_n1264));
  XOR2_X1   g1064(.A(new_n1017), .B(KEYINPUT120), .Z(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1142), .A2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1137), .B1(new_n1141), .B2(new_n1117), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1264), .B1(new_n1267), .B2(new_n1268), .ZN(G381));
  INV_X1    g1069(.A(new_n1166), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1270), .B1(new_n1237), .B2(new_n756), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1145), .A2(new_n709), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1240), .A2(new_n1142), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1271), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT123), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1146), .A2(KEYINPUT123), .A3(new_n1271), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1245), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(G393), .A2(G396), .ZN(new_n1280));
  INV_X1    g1080(.A(G384), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1280), .A2(new_n1281), .A3(new_n1105), .ZN(new_n1282));
  OR4_X1    g1082(.A1(G387), .A2(new_n1279), .A3(G381), .A4(new_n1282), .ZN(G407));
  OAI211_X1 g1083(.A(G407), .B(G213), .C1(G343), .C2(new_n1279), .ZN(G409));
  AOI21_X1  g1084(.A(new_n826), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1280), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(G387), .A2(new_n1105), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1038), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n750), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n755), .B1(new_n1290), .B2(new_n1017), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(new_n982), .A3(G390), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1288), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT124), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1287), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  AOI211_X1 g1096(.A(KEYINPUT124), .B(new_n1286), .C1(new_n1288), .C2(new_n1293), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT125), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1268), .B1(KEYINPUT60), .B2(new_n1142), .ZN(new_n1301));
  OAI211_X1 g1101(.A(new_n1241), .B(KEYINPUT60), .C1(new_n1112), .C2(new_n1118), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n709), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1264), .B1(new_n1301), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1281), .ZN(new_n1305));
  OAI211_X1 g1105(.A(G384), .B(new_n1264), .C1(new_n1301), .C2(new_n1303), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n685), .A2(G343), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(G2897), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1305), .A2(new_n1306), .A3(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1308), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1233), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1242), .A2(new_n1312), .A3(new_n1266), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1234), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  AOI22_X1  g1115(.A1(new_n1278), .A2(new_n1315), .B1(new_n1245), .B2(G378), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1311), .B1(new_n1316), .B2(new_n1307), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT61), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1300), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  AND3_X1   g1119(.A1(new_n1146), .A2(KEYINPUT123), .A3(new_n1271), .ZN(new_n1320));
  AOI21_X1  g1120(.A(KEYINPUT123), .B1(new_n1146), .B2(new_n1271), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1315), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(KEYINPUT57), .B1(new_n1242), .B2(new_n1312), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1219), .A2(new_n1232), .A3(KEYINPUT57), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n709), .B1(new_n1238), .B2(new_n1324), .ZN(new_n1325));
  OAI211_X1 g1125(.A(G378), .B(new_n1314), .C1(new_n1323), .C2(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1307), .B1(new_n1322), .B2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1308), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1268), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1142), .A2(KEYINPUT60), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1331), .A2(new_n709), .A3(new_n1302), .ZN(new_n1332));
  AOI21_X1  g1132(.A(G384), .B1(new_n1332), .B2(new_n1264), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1306), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1328), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1305), .A2(new_n1306), .A3(new_n1308), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  OAI211_X1 g1137(.A(new_n1300), .B(new_n1318), .C1(new_n1327), .C2(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1338), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1319), .A2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT62), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1342));
  AOI211_X1 g1142(.A(new_n1307), .B(new_n1342), .C1(new_n1322), .C2(new_n1326), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT126), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1341), .B1(new_n1343), .B2(new_n1344), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1342), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1327), .A2(new_n1346), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1347), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1345), .A2(new_n1348), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1299), .B1(new_n1340), .B2(new_n1349), .ZN(new_n1350));
  XNOR2_X1  g1150(.A(new_n1347), .B(KEYINPUT63), .ZN(new_n1351));
  NAND4_X1  g1151(.A1(new_n1351), .A2(new_n1318), .A3(new_n1298), .A4(new_n1317), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1350), .A2(new_n1352), .ZN(G405));
  NOR2_X1   g1153(.A1(new_n1346), .A2(KEYINPUT127), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1354), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1346), .A2(KEYINPUT127), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(G375), .A2(new_n1278), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1356), .A2(new_n1357), .A3(new_n1326), .ZN(new_n1358));
  INV_X1    g1158(.A(new_n1358), .ZN(new_n1359));
  AOI21_X1  g1159(.A(G390), .B1(new_n1292), .B2(new_n982), .ZN(new_n1360));
  INV_X1    g1160(.A(new_n982), .ZN(new_n1361));
  AOI211_X1 g1161(.A(new_n1361), .B(new_n1105), .C1(new_n1289), .C2(new_n1291), .ZN(new_n1362));
  OAI21_X1  g1162(.A(new_n1295), .B1(new_n1360), .B2(new_n1362), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1363), .A2(new_n1286), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1294), .A2(new_n1295), .A3(new_n1287), .ZN(new_n1365));
  INV_X1    g1165(.A(new_n1354), .ZN(new_n1366));
  NAND3_X1  g1166(.A1(new_n1364), .A2(new_n1365), .A3(new_n1366), .ZN(new_n1367));
  AND3_X1   g1167(.A1(new_n1355), .A2(new_n1359), .A3(new_n1367), .ZN(new_n1368));
  AOI21_X1  g1168(.A(new_n1359), .B1(new_n1355), .B2(new_n1367), .ZN(new_n1369));
  NOR2_X1   g1169(.A1(new_n1368), .A2(new_n1369), .ZN(G402));
endmodule


