

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U550 ( .A1(n539), .A2(n538), .ZN(G160) );
  BUF_X1 U551 ( .A(n896), .Z(n518) );
  NOR2_X1 U552 ( .A1(G2105), .A2(n524), .ZN(n896) );
  NOR2_X1 U553 ( .A1(n695), .A2(n933), .ZN(n690) );
  NOR2_X1 U554 ( .A1(n645), .A2(G651), .ZN(n647) );
  AND2_X1 U555 ( .A1(n834), .A2(n833), .ZN(n836) );
  NOR2_X1 U556 ( .A1(n528), .A2(n527), .ZN(G164) );
  INV_X1 U557 ( .A(G2104), .ZN(n524) );
  NAND2_X1 U558 ( .A1(n518), .A2(G102), .ZN(n522) );
  NOR2_X1 U559 ( .A1(G2104), .A2(G2105), .ZN(n519) );
  XOR2_X1 U560 ( .A(KEYINPUT17), .B(n519), .Z(n520) );
  XNOR2_X1 U561 ( .A(KEYINPUT68), .B(n520), .ZN(n747) );
  NAND2_X1 U562 ( .A1(G138), .A2(n747), .ZN(n521) );
  NAND2_X1 U563 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U564 ( .A(KEYINPUT88), .B(n523), .ZN(n528) );
  AND2_X1 U565 ( .A1(n524), .A2(G2105), .ZN(n902) );
  NAND2_X1 U566 ( .A1(G126), .A2(n902), .ZN(n526) );
  AND2_X1 U567 ( .A1(G2104), .A2(G2105), .ZN(n900) );
  NAND2_X1 U568 ( .A1(G114), .A2(n900), .ZN(n525) );
  NAND2_X1 U569 ( .A1(n526), .A2(n525), .ZN(n527) );
  NAND2_X1 U570 ( .A1(n900), .A2(G113), .ZN(n530) );
  NAND2_X1 U571 ( .A1(G137), .A2(n747), .ZN(n529) );
  NAND2_X1 U572 ( .A1(n530), .A2(n529), .ZN(n539) );
  NAND2_X1 U573 ( .A1(G101), .A2(n896), .ZN(n531) );
  XNOR2_X1 U574 ( .A(n531), .B(KEYINPUT23), .ZN(n533) );
  INV_X1 U575 ( .A(KEYINPUT66), .ZN(n532) );
  XNOR2_X1 U576 ( .A(n533), .B(n532), .ZN(n535) );
  NAND2_X1 U577 ( .A1(G125), .A2(n902), .ZN(n534) );
  NAND2_X1 U578 ( .A1(n535), .A2(n534), .ZN(n537) );
  INV_X1 U579 ( .A(KEYINPUT67), .ZN(n536) );
  XNOR2_X1 U580 ( .A(n537), .B(n536), .ZN(n538) );
  AND2_X1 U581 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U582 ( .A(G57), .ZN(G237) );
  INV_X1 U583 ( .A(G132), .ZN(G219) );
  INV_X1 U584 ( .A(G82), .ZN(G220) );
  NOR2_X1 U585 ( .A1(G543), .A2(G651), .ZN(n636) );
  NAND2_X1 U586 ( .A1(G88), .A2(n636), .ZN(n541) );
  XOR2_X1 U587 ( .A(KEYINPUT0), .B(G543), .Z(n645) );
  XNOR2_X1 U588 ( .A(KEYINPUT69), .B(G651), .ZN(n542) );
  NOR2_X1 U589 ( .A1(n645), .A2(n542), .ZN(n639) );
  NAND2_X1 U590 ( .A1(G75), .A2(n639), .ZN(n540) );
  NAND2_X1 U591 ( .A1(n541), .A2(n540), .ZN(n547) );
  NAND2_X1 U592 ( .A1(n647), .A2(G50), .ZN(n545) );
  NOR2_X1 U593 ( .A1(G543), .A2(n542), .ZN(n543) );
  XOR2_X1 U594 ( .A(KEYINPUT1), .B(n543), .Z(n651) );
  NAND2_X1 U595 ( .A1(G62), .A2(n651), .ZN(n544) );
  NAND2_X1 U596 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U597 ( .A1(n547), .A2(n546), .ZN(G166) );
  NAND2_X1 U598 ( .A1(n647), .A2(G52), .ZN(n549) );
  NAND2_X1 U599 ( .A1(G64), .A2(n651), .ZN(n548) );
  NAND2_X1 U600 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U601 ( .A(KEYINPUT71), .B(n550), .Z(n556) );
  NAND2_X1 U602 ( .A1(n636), .A2(G90), .ZN(n551) );
  XNOR2_X1 U603 ( .A(n551), .B(KEYINPUT72), .ZN(n553) );
  NAND2_X1 U604 ( .A1(G77), .A2(n639), .ZN(n552) );
  NAND2_X1 U605 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U606 ( .A(KEYINPUT9), .B(n554), .Z(n555) );
  NOR2_X1 U607 ( .A1(n556), .A2(n555), .ZN(G171) );
  XNOR2_X1 U608 ( .A(KEYINPUT76), .B(KEYINPUT7), .ZN(n568) );
  NAND2_X1 U609 ( .A1(n636), .A2(G89), .ZN(n557) );
  XNOR2_X1 U610 ( .A(n557), .B(KEYINPUT4), .ZN(n559) );
  NAND2_X1 U611 ( .A1(G76), .A2(n639), .ZN(n558) );
  NAND2_X1 U612 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U613 ( .A(n560), .B(KEYINPUT5), .ZN(n566) );
  XNOR2_X1 U614 ( .A(KEYINPUT6), .B(KEYINPUT75), .ZN(n564) );
  NAND2_X1 U615 ( .A1(n647), .A2(G51), .ZN(n562) );
  NAND2_X1 U616 ( .A1(G63), .A2(n651), .ZN(n561) );
  NAND2_X1 U617 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U618 ( .A(n564), .B(n563), .ZN(n565) );
  NAND2_X1 U619 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U620 ( .A(n568), .B(n567), .ZN(G168) );
  XNOR2_X1 U621 ( .A(KEYINPUT77), .B(KEYINPUT8), .ZN(n569) );
  XNOR2_X1 U622 ( .A(n569), .B(G168), .ZN(G286) );
  NAND2_X1 U623 ( .A1(G7), .A2(G661), .ZN(n570) );
  XNOR2_X1 U624 ( .A(n570), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U625 ( .A(G223), .ZN(n837) );
  NAND2_X1 U626 ( .A1(n837), .A2(G567), .ZN(n571) );
  XNOR2_X1 U627 ( .A(n571), .B(KEYINPUT11), .ZN(n572) );
  XNOR2_X1 U628 ( .A(KEYINPUT73), .B(n572), .ZN(G234) );
  NAND2_X1 U629 ( .A1(n651), .A2(G56), .ZN(n573) );
  XOR2_X1 U630 ( .A(KEYINPUT14), .B(n573), .Z(n579) );
  NAND2_X1 U631 ( .A1(n636), .A2(G81), .ZN(n574) );
  XNOR2_X1 U632 ( .A(n574), .B(KEYINPUT12), .ZN(n576) );
  NAND2_X1 U633 ( .A1(G68), .A2(n639), .ZN(n575) );
  NAND2_X1 U634 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U635 ( .A(KEYINPUT13), .B(n577), .Z(n578) );
  NOR2_X1 U636 ( .A1(n579), .A2(n578), .ZN(n581) );
  NAND2_X1 U637 ( .A1(n647), .A2(G43), .ZN(n580) );
  NAND2_X1 U638 ( .A1(n581), .A2(n580), .ZN(n934) );
  INV_X1 U639 ( .A(G860), .ZN(n600) );
  OR2_X1 U640 ( .A1(n934), .A2(n600), .ZN(G153) );
  INV_X1 U641 ( .A(G171), .ZN(G301) );
  NAND2_X1 U642 ( .A1(G868), .A2(G301), .ZN(n591) );
  NAND2_X1 U643 ( .A1(G79), .A2(n639), .ZN(n588) );
  NAND2_X1 U644 ( .A1(G92), .A2(n636), .ZN(n583) );
  NAND2_X1 U645 ( .A1(G54), .A2(n647), .ZN(n582) );
  NAND2_X1 U646 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U647 ( .A1(n651), .A2(G66), .ZN(n584) );
  XOR2_X1 U648 ( .A(KEYINPUT74), .B(n584), .Z(n585) );
  NOR2_X1 U649 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U650 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U651 ( .A(KEYINPUT15), .B(n589), .Z(n933) );
  INV_X1 U652 ( .A(G868), .ZN(n665) );
  NAND2_X1 U653 ( .A1(n933), .A2(n665), .ZN(n590) );
  NAND2_X1 U654 ( .A1(n591), .A2(n590), .ZN(G284) );
  NAND2_X1 U655 ( .A1(n647), .A2(G53), .ZN(n593) );
  NAND2_X1 U656 ( .A1(G65), .A2(n651), .ZN(n592) );
  NAND2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n597) );
  NAND2_X1 U658 ( .A1(G91), .A2(n636), .ZN(n595) );
  NAND2_X1 U659 ( .A1(G78), .A2(n639), .ZN(n594) );
  NAND2_X1 U660 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U661 ( .A1(n597), .A2(n596), .ZN(n937) );
  INV_X1 U662 ( .A(n937), .ZN(G299) );
  NAND2_X1 U663 ( .A1(G868), .A2(G286), .ZN(n599) );
  NAND2_X1 U664 ( .A1(G299), .A2(n665), .ZN(n598) );
  NAND2_X1 U665 ( .A1(n599), .A2(n598), .ZN(G297) );
  NAND2_X1 U666 ( .A1(G559), .A2(n600), .ZN(n601) );
  XNOR2_X1 U667 ( .A(KEYINPUT78), .B(n601), .ZN(n602) );
  INV_X1 U668 ( .A(n933), .ZN(n918) );
  NAND2_X1 U669 ( .A1(n602), .A2(n918), .ZN(n603) );
  XNOR2_X1 U670 ( .A(KEYINPUT16), .B(n603), .ZN(G148) );
  NOR2_X1 U671 ( .A1(G868), .A2(n934), .ZN(n606) );
  NAND2_X1 U672 ( .A1(G868), .A2(n918), .ZN(n604) );
  NOR2_X1 U673 ( .A1(G559), .A2(n604), .ZN(n605) );
  NOR2_X1 U674 ( .A1(n606), .A2(n605), .ZN(G282) );
  NAND2_X1 U675 ( .A1(G123), .A2(n902), .ZN(n607) );
  XOR2_X1 U676 ( .A(KEYINPUT79), .B(n607), .Z(n608) );
  XNOR2_X1 U677 ( .A(n608), .B(KEYINPUT18), .ZN(n610) );
  NAND2_X1 U678 ( .A1(G99), .A2(n518), .ZN(n609) );
  NAND2_X1 U679 ( .A1(n610), .A2(n609), .ZN(n614) );
  NAND2_X1 U680 ( .A1(n900), .A2(G111), .ZN(n612) );
  BUF_X1 U681 ( .A(n747), .Z(n897) );
  NAND2_X1 U682 ( .A1(G135), .A2(n897), .ZN(n611) );
  NAND2_X1 U683 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U684 ( .A1(n614), .A2(n613), .ZN(n1015) );
  XNOR2_X1 U685 ( .A(n1015), .B(G2096), .ZN(n615) );
  XNOR2_X1 U686 ( .A(n615), .B(KEYINPUT80), .ZN(n617) );
  INV_X1 U687 ( .A(G2100), .ZN(n616) );
  NAND2_X1 U688 ( .A1(n617), .A2(n616), .ZN(G156) );
  NAND2_X1 U689 ( .A1(G93), .A2(n636), .ZN(n619) );
  NAND2_X1 U690 ( .A1(G55), .A2(n647), .ZN(n618) );
  NAND2_X1 U691 ( .A1(n619), .A2(n618), .ZN(n622) );
  NAND2_X1 U692 ( .A1(G80), .A2(n639), .ZN(n620) );
  XNOR2_X1 U693 ( .A(KEYINPUT81), .B(n620), .ZN(n621) );
  NOR2_X1 U694 ( .A1(n622), .A2(n621), .ZN(n624) );
  NAND2_X1 U695 ( .A1(G67), .A2(n651), .ZN(n623) );
  NAND2_X1 U696 ( .A1(n624), .A2(n623), .ZN(n664) );
  NAND2_X1 U697 ( .A1(n918), .A2(G559), .ZN(n662) );
  XNOR2_X1 U698 ( .A(n934), .B(n662), .ZN(n625) );
  NOR2_X1 U699 ( .A1(G860), .A2(n625), .ZN(n626) );
  XOR2_X1 U700 ( .A(n664), .B(n626), .Z(G145) );
  NAND2_X1 U701 ( .A1(n639), .A2(G73), .ZN(n627) );
  XNOR2_X1 U702 ( .A(n627), .B(KEYINPUT2), .ZN(n635) );
  NAND2_X1 U703 ( .A1(n636), .A2(G86), .ZN(n628) );
  XNOR2_X1 U704 ( .A(n628), .B(KEYINPUT86), .ZN(n630) );
  NAND2_X1 U705 ( .A1(G48), .A2(n647), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U707 ( .A1(G61), .A2(n651), .ZN(n631) );
  XNOR2_X1 U708 ( .A(KEYINPUT85), .B(n631), .ZN(n632) );
  NOR2_X1 U709 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U710 ( .A1(n635), .A2(n634), .ZN(G305) );
  NAND2_X1 U711 ( .A1(n636), .A2(G85), .ZN(n638) );
  NAND2_X1 U712 ( .A1(G60), .A2(n651), .ZN(n637) );
  NAND2_X1 U713 ( .A1(n638), .A2(n637), .ZN(n643) );
  NAND2_X1 U714 ( .A1(n647), .A2(G47), .ZN(n641) );
  NAND2_X1 U715 ( .A1(G72), .A2(n639), .ZN(n640) );
  NAND2_X1 U716 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U717 ( .A1(n643), .A2(n642), .ZN(n644) );
  XOR2_X1 U718 ( .A(KEYINPUT70), .B(n644), .Z(G290) );
  NAND2_X1 U719 ( .A1(n645), .A2(G87), .ZN(n646) );
  XNOR2_X1 U720 ( .A(KEYINPUT83), .B(n646), .ZN(n654) );
  NAND2_X1 U721 ( .A1(G49), .A2(n647), .ZN(n649) );
  NAND2_X1 U722 ( .A1(G74), .A2(G651), .ZN(n648) );
  NAND2_X1 U723 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U724 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U725 ( .A(KEYINPUT82), .B(n652), .Z(n653) );
  NOR2_X1 U726 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U727 ( .A(KEYINPUT84), .B(n655), .Z(G288) );
  XOR2_X1 U728 ( .A(G290), .B(G288), .Z(n656) );
  XNOR2_X1 U729 ( .A(G305), .B(n656), .ZN(n657) );
  XNOR2_X1 U730 ( .A(KEYINPUT19), .B(n657), .ZN(n659) );
  XNOR2_X1 U731 ( .A(n934), .B(G166), .ZN(n658) );
  XNOR2_X1 U732 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U733 ( .A(n937), .B(n660), .ZN(n661) );
  XNOR2_X1 U734 ( .A(n661), .B(n664), .ZN(n917) );
  XNOR2_X1 U735 ( .A(n662), .B(n917), .ZN(n663) );
  NAND2_X1 U736 ( .A1(n663), .A2(G868), .ZN(n667) );
  NAND2_X1 U737 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U738 ( .A1(n667), .A2(n666), .ZN(G295) );
  XOR2_X1 U739 ( .A(KEYINPUT21), .B(KEYINPUT87), .Z(n671) );
  NAND2_X1 U740 ( .A1(G2078), .A2(G2084), .ZN(n668) );
  XOR2_X1 U741 ( .A(KEYINPUT20), .B(n668), .Z(n669) );
  NAND2_X1 U742 ( .A1(n669), .A2(G2090), .ZN(n670) );
  XNOR2_X1 U743 ( .A(n671), .B(n670), .ZN(n672) );
  NAND2_X1 U744 ( .A1(G2072), .A2(n672), .ZN(G158) );
  XNOR2_X1 U745 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U746 ( .A1(G220), .A2(G219), .ZN(n673) );
  XOR2_X1 U747 ( .A(KEYINPUT22), .B(n673), .Z(n674) );
  NOR2_X1 U748 ( .A1(G218), .A2(n674), .ZN(n675) );
  NAND2_X1 U749 ( .A1(G96), .A2(n675), .ZN(n841) );
  NAND2_X1 U750 ( .A1(n841), .A2(G2106), .ZN(n679) );
  NAND2_X1 U751 ( .A1(G69), .A2(G120), .ZN(n676) );
  NOR2_X1 U752 ( .A1(G237), .A2(n676), .ZN(n677) );
  NAND2_X1 U753 ( .A1(G108), .A2(n677), .ZN(n842) );
  NAND2_X1 U754 ( .A1(n842), .A2(G567), .ZN(n678) );
  NAND2_X1 U755 ( .A1(n679), .A2(n678), .ZN(n854) );
  NAND2_X1 U756 ( .A1(G661), .A2(G483), .ZN(n680) );
  NOR2_X1 U757 ( .A1(n854), .A2(n680), .ZN(n840) );
  NAND2_X1 U758 ( .A1(n840), .A2(G36), .ZN(G176) );
  INV_X1 U759 ( .A(G166), .ZN(G303) );
  NOR2_X1 U760 ( .A1(G164), .A2(G1384), .ZN(n681) );
  XNOR2_X1 U761 ( .A(KEYINPUT65), .B(n681), .ZN(n763) );
  INV_X1 U762 ( .A(KEYINPUT92), .ZN(n682) );
  AND2_X1 U763 ( .A1(G160), .A2(G40), .ZN(n764) );
  XNOR2_X1 U764 ( .A(n682), .B(n764), .ZN(n683) );
  NOR2_X1 U765 ( .A1(n763), .A2(n683), .ZN(n684) );
  XNOR2_X1 U766 ( .A(n684), .B(KEYINPUT64), .ZN(n687) );
  AND2_X1 U767 ( .A1(G1996), .A2(n687), .ZN(n685) );
  XNOR2_X1 U768 ( .A(n685), .B(KEYINPUT26), .ZN(n686) );
  NOR2_X1 U769 ( .A1(n934), .A2(n686), .ZN(n689) );
  INV_X1 U770 ( .A(n687), .ZN(n729) );
  NAND2_X1 U771 ( .A1(n729), .A2(G1341), .ZN(n688) );
  NAND2_X1 U772 ( .A1(n689), .A2(n688), .ZN(n695) );
  XNOR2_X1 U773 ( .A(n690), .B(KEYINPUT97), .ZN(n694) );
  INV_X1 U774 ( .A(n729), .ZN(n710) );
  NOR2_X1 U775 ( .A1(G1348), .A2(n710), .ZN(n692) );
  NOR2_X1 U776 ( .A1(G2067), .A2(n729), .ZN(n691) );
  NOR2_X1 U777 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U778 ( .A1(n694), .A2(n693), .ZN(n697) );
  NAND2_X1 U779 ( .A1(n695), .A2(n933), .ZN(n696) );
  NAND2_X1 U780 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U781 ( .A(n698), .B(KEYINPUT98), .ZN(n703) );
  NAND2_X1 U782 ( .A1(G2072), .A2(n710), .ZN(n699) );
  XNOR2_X1 U783 ( .A(n699), .B(KEYINPUT27), .ZN(n701) );
  INV_X1 U784 ( .A(G1956), .ZN(n958) );
  NOR2_X1 U785 ( .A1(n710), .A2(n958), .ZN(n700) );
  NOR2_X1 U786 ( .A1(n701), .A2(n700), .ZN(n704) );
  NAND2_X1 U787 ( .A1(n704), .A2(n937), .ZN(n702) );
  NAND2_X1 U788 ( .A1(n703), .A2(n702), .ZN(n708) );
  NOR2_X1 U789 ( .A1(n704), .A2(n937), .ZN(n706) );
  XOR2_X1 U790 ( .A(KEYINPUT96), .B(KEYINPUT28), .Z(n705) );
  XNOR2_X1 U791 ( .A(n706), .B(n705), .ZN(n707) );
  NAND2_X1 U792 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U793 ( .A(KEYINPUT29), .B(n709), .ZN(n715) );
  NOR2_X1 U794 ( .A1(G1961), .A2(n710), .ZN(n712) );
  XOR2_X1 U795 ( .A(KEYINPUT25), .B(G2078), .Z(n983) );
  NOR2_X1 U796 ( .A1(n729), .A2(n983), .ZN(n711) );
  NOR2_X1 U797 ( .A1(n712), .A2(n711), .ZN(n720) );
  NOR2_X1 U798 ( .A1(n720), .A2(G301), .ZN(n713) );
  XOR2_X1 U799 ( .A(KEYINPUT95), .B(n713), .Z(n714) );
  NOR2_X1 U800 ( .A1(n715), .A2(n714), .ZN(n725) );
  NAND2_X1 U801 ( .A1(n729), .A2(G8), .ZN(n802) );
  NOR2_X1 U802 ( .A1(G1966), .A2(n802), .ZN(n743) );
  NOR2_X1 U803 ( .A1(n729), .A2(G2084), .ZN(n716) );
  XNOR2_X1 U804 ( .A(KEYINPUT93), .B(n716), .ZN(n739) );
  NAND2_X1 U805 ( .A1(G8), .A2(n739), .ZN(n717) );
  NOR2_X1 U806 ( .A1(n743), .A2(n717), .ZN(n718) );
  XOR2_X1 U807 ( .A(KEYINPUT30), .B(n718), .Z(n719) );
  NOR2_X1 U808 ( .A1(G168), .A2(n719), .ZN(n722) );
  AND2_X1 U809 ( .A1(G301), .A2(n720), .ZN(n721) );
  NOR2_X1 U810 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U811 ( .A(n723), .B(KEYINPUT31), .ZN(n724) );
  NOR2_X2 U812 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U813 ( .A(n726), .B(KEYINPUT99), .ZN(n744) );
  AND2_X1 U814 ( .A1(G286), .A2(G8), .ZN(n727) );
  NAND2_X1 U815 ( .A1(n744), .A2(n727), .ZN(n736) );
  INV_X1 U816 ( .A(G8), .ZN(n734) );
  NOR2_X1 U817 ( .A1(G1971), .A2(n802), .ZN(n728) );
  XNOR2_X1 U818 ( .A(n728), .B(KEYINPUT100), .ZN(n731) );
  NOR2_X1 U819 ( .A1(n729), .A2(G2090), .ZN(n730) );
  NOR2_X1 U820 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U821 ( .A1(n732), .A2(G303), .ZN(n733) );
  OR2_X1 U822 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U823 ( .A1(n736), .A2(n735), .ZN(n738) );
  INV_X1 U824 ( .A(KEYINPUT32), .ZN(n737) );
  XNOR2_X1 U825 ( .A(n738), .B(n737), .ZN(n820) );
  INV_X1 U826 ( .A(n739), .ZN(n740) );
  NAND2_X1 U827 ( .A1(G8), .A2(n740), .ZN(n741) );
  XOR2_X1 U828 ( .A(KEYINPUT94), .B(n741), .Z(n742) );
  NOR2_X1 U829 ( .A1(n743), .A2(n742), .ZN(n745) );
  NAND2_X1 U830 ( .A1(n745), .A2(n744), .ZN(n816) );
  NAND2_X1 U831 ( .A1(G105), .A2(n518), .ZN(n746) );
  XNOR2_X1 U832 ( .A(n746), .B(KEYINPUT38), .ZN(n754) );
  NAND2_X1 U833 ( .A1(n902), .A2(G129), .ZN(n749) );
  NAND2_X1 U834 ( .A1(G141), .A2(n747), .ZN(n748) );
  NAND2_X1 U835 ( .A1(n749), .A2(n748), .ZN(n752) );
  NAND2_X1 U836 ( .A1(n900), .A2(G117), .ZN(n750) );
  XOR2_X1 U837 ( .A(KEYINPUT90), .B(n750), .Z(n751) );
  NOR2_X1 U838 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U839 ( .A1(n754), .A2(n753), .ZN(n911) );
  NOR2_X1 U840 ( .A1(G1996), .A2(n911), .ZN(n1009) );
  NAND2_X1 U841 ( .A1(n902), .A2(G119), .ZN(n756) );
  NAND2_X1 U842 ( .A1(G131), .A2(n897), .ZN(n755) );
  NAND2_X1 U843 ( .A1(n756), .A2(n755), .ZN(n760) );
  NAND2_X1 U844 ( .A1(G95), .A2(n518), .ZN(n758) );
  NAND2_X1 U845 ( .A1(G107), .A2(n900), .ZN(n757) );
  NAND2_X1 U846 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U847 ( .A1(n760), .A2(n759), .ZN(n892) );
  INV_X1 U848 ( .A(G1991), .ZN(n765) );
  NOR2_X1 U849 ( .A1(n892), .A2(n765), .ZN(n762) );
  AND2_X1 U850 ( .A1(n911), .A2(G1996), .ZN(n761) );
  NOR2_X1 U851 ( .A1(n762), .A2(n761), .ZN(n1007) );
  NAND2_X1 U852 ( .A1(n764), .A2(n763), .ZN(n771) );
  NOR2_X1 U853 ( .A1(n1007), .A2(n771), .ZN(n824) );
  NOR2_X1 U854 ( .A1(G1986), .A2(G290), .ZN(n767) );
  AND2_X1 U855 ( .A1(n765), .A2(n892), .ZN(n766) );
  XNOR2_X1 U856 ( .A(KEYINPUT102), .B(n766), .ZN(n1017) );
  NOR2_X1 U857 ( .A1(n767), .A2(n1017), .ZN(n768) );
  NOR2_X1 U858 ( .A1(n824), .A2(n768), .ZN(n769) );
  NOR2_X1 U859 ( .A1(n1009), .A2(n769), .ZN(n770) );
  XNOR2_X1 U860 ( .A(KEYINPUT39), .B(n770), .ZN(n782) );
  INV_X1 U861 ( .A(n771), .ZN(n828) );
  XNOR2_X1 U862 ( .A(G2067), .B(KEYINPUT37), .ZN(n783) );
  NAND2_X1 U863 ( .A1(n518), .A2(G104), .ZN(n772) );
  XOR2_X1 U864 ( .A(KEYINPUT89), .B(n772), .Z(n774) );
  NAND2_X1 U865 ( .A1(G140), .A2(n897), .ZN(n773) );
  NAND2_X1 U866 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U867 ( .A(KEYINPUT34), .B(n775), .ZN(n780) );
  NAND2_X1 U868 ( .A1(G128), .A2(n902), .ZN(n777) );
  NAND2_X1 U869 ( .A1(G116), .A2(n900), .ZN(n776) );
  NAND2_X1 U870 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U871 ( .A(KEYINPUT35), .B(n778), .Z(n779) );
  NOR2_X1 U872 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U873 ( .A(KEYINPUT36), .B(n781), .ZN(n914) );
  NOR2_X1 U874 ( .A1(n783), .A2(n914), .ZN(n1016) );
  NAND2_X1 U875 ( .A1(n828), .A2(n1016), .ZN(n826) );
  NAND2_X1 U876 ( .A1(n782), .A2(n826), .ZN(n784) );
  NAND2_X1 U877 ( .A1(n783), .A2(n914), .ZN(n1006) );
  NAND2_X1 U878 ( .A1(n784), .A2(n1006), .ZN(n785) );
  NAND2_X1 U879 ( .A1(n785), .A2(n828), .ZN(n823) );
  NOR2_X1 U880 ( .A1(G1981), .A2(G305), .ZN(n786) );
  XNOR2_X1 U881 ( .A(KEYINPUT24), .B(n786), .ZN(n787) );
  INV_X1 U882 ( .A(n802), .ZN(n797) );
  NAND2_X1 U883 ( .A1(n787), .A2(n797), .ZN(n788) );
  AND2_X1 U884 ( .A1(n823), .A2(n788), .ZN(n793) );
  INV_X1 U885 ( .A(n793), .ZN(n789) );
  OR2_X1 U886 ( .A1(n789), .A2(n802), .ZN(n791) );
  AND2_X1 U887 ( .A1(n816), .A2(n791), .ZN(n790) );
  AND2_X1 U888 ( .A1(n820), .A2(n790), .ZN(n813) );
  INV_X1 U889 ( .A(n791), .ZN(n796) );
  NOR2_X1 U890 ( .A1(G2090), .A2(G303), .ZN(n792) );
  NAND2_X1 U891 ( .A1(G8), .A2(n792), .ZN(n794) );
  AND2_X1 U892 ( .A1(n794), .A2(n793), .ZN(n795) );
  OR2_X1 U893 ( .A1(n796), .A2(n795), .ZN(n811) );
  XNOR2_X1 U894 ( .A(G1981), .B(G305), .ZN(n930) );
  INV_X1 U895 ( .A(n930), .ZN(n801) );
  INV_X1 U896 ( .A(KEYINPUT33), .ZN(n806) );
  NOR2_X1 U897 ( .A1(G1976), .A2(G288), .ZN(n944) );
  NAND2_X1 U898 ( .A1(n797), .A2(n944), .ZN(n798) );
  NOR2_X1 U899 ( .A1(n806), .A2(n798), .ZN(n799) );
  XNOR2_X1 U900 ( .A(n799), .B(KEYINPUT101), .ZN(n800) );
  AND2_X1 U901 ( .A1(n801), .A2(n800), .ZN(n817) );
  INV_X1 U902 ( .A(n817), .ZN(n809) );
  NAND2_X1 U903 ( .A1(G1976), .A2(G288), .ZN(n938) );
  INV_X1 U904 ( .A(n938), .ZN(n803) );
  OR2_X1 U905 ( .A1(n803), .A2(n802), .ZN(n814) );
  INV_X1 U906 ( .A(G1971), .ZN(n967) );
  AND2_X1 U907 ( .A1(G166), .A2(n967), .ZN(n804) );
  NOR2_X1 U908 ( .A1(n804), .A2(n944), .ZN(n805) );
  OR2_X1 U909 ( .A1(n814), .A2(n805), .ZN(n807) );
  AND2_X1 U910 ( .A1(n807), .A2(n806), .ZN(n808) );
  OR2_X1 U911 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U912 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U913 ( .A1(n813), .A2(n812), .ZN(n822) );
  INV_X1 U914 ( .A(n814), .ZN(n815) );
  AND2_X1 U915 ( .A1(n816), .A2(n815), .ZN(n818) );
  AND2_X1 U916 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U917 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U918 ( .A1(n822), .A2(n821), .ZN(n834) );
  INV_X1 U919 ( .A(n823), .ZN(n832) );
  INV_X1 U920 ( .A(n824), .ZN(n825) );
  NAND2_X1 U921 ( .A1(n826), .A2(n825), .ZN(n827) );
  XOR2_X1 U922 ( .A(KEYINPUT91), .B(n827), .Z(n830) );
  XNOR2_X1 U923 ( .A(G1986), .B(G290), .ZN(n946) );
  AND2_X1 U924 ( .A1(n946), .A2(n828), .ZN(n829) );
  NOR2_X1 U925 ( .A1(n830), .A2(n829), .ZN(n831) );
  OR2_X1 U926 ( .A1(n832), .A2(n831), .ZN(n833) );
  XOR2_X1 U927 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n835) );
  XNOR2_X1 U928 ( .A(n836), .B(n835), .ZN(G329) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n837), .ZN(G217) );
  AND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U931 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U933 ( .A1(n840), .A2(n839), .ZN(G188) );
  XOR2_X1 U934 ( .A(G96), .B(KEYINPUT106), .Z(G221) );
  INV_X1 U936 ( .A(G120), .ZN(G236) );
  INV_X1 U937 ( .A(G69), .ZN(G235) );
  NOR2_X1 U938 ( .A1(n842), .A2(n841), .ZN(G325) );
  INV_X1 U939 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U940 ( .A(KEYINPUT104), .B(G2454), .ZN(n851) );
  XNOR2_X1 U941 ( .A(G2430), .B(G2435), .ZN(n849) );
  XOR2_X1 U942 ( .A(G2451), .B(G2427), .Z(n844) );
  XNOR2_X1 U943 ( .A(G2438), .B(G2446), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U945 ( .A(n845), .B(G2443), .Z(n847) );
  XNOR2_X1 U946 ( .A(G1341), .B(G1348), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U949 ( .A(n851), .B(n850), .ZN(n852) );
  NAND2_X1 U950 ( .A1(n852), .A2(G14), .ZN(n853) );
  XNOR2_X1 U951 ( .A(KEYINPUT105), .B(n853), .ZN(G401) );
  INV_X1 U952 ( .A(n854), .ZN(G319) );
  XNOR2_X1 U953 ( .A(G1991), .B(KEYINPUT41), .ZN(n864) );
  XOR2_X1 U954 ( .A(G1981), .B(G1961), .Z(n856) );
  XNOR2_X1 U955 ( .A(G1996), .B(G1966), .ZN(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U957 ( .A(G1976), .B(G1971), .Z(n858) );
  XNOR2_X1 U958 ( .A(G1986), .B(G1956), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U960 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U961 ( .A(KEYINPUT108), .B(G2474), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n862), .B(n861), .ZN(n863) );
  XNOR2_X1 U963 ( .A(n864), .B(n863), .ZN(G229) );
  XOR2_X1 U964 ( .A(G2678), .B(G2090), .Z(n866) );
  XNOR2_X1 U965 ( .A(G2067), .B(G2084), .ZN(n865) );
  XNOR2_X1 U966 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U967 ( .A(n867), .B(G2096), .Z(n869) );
  XNOR2_X1 U968 ( .A(G2078), .B(G2072), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n869), .B(n868), .ZN(n873) );
  XOR2_X1 U970 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n871) );
  XNOR2_X1 U971 ( .A(KEYINPUT42), .B(G2100), .ZN(n870) );
  XNOR2_X1 U972 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U973 ( .A(n873), .B(n872), .Z(G227) );
  NAND2_X1 U974 ( .A1(G124), .A2(n902), .ZN(n874) );
  XOR2_X1 U975 ( .A(KEYINPUT44), .B(n874), .Z(n875) );
  XNOR2_X1 U976 ( .A(n875), .B(KEYINPUT109), .ZN(n877) );
  NAND2_X1 U977 ( .A1(G136), .A2(n897), .ZN(n876) );
  NAND2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n881) );
  NAND2_X1 U979 ( .A1(G100), .A2(n518), .ZN(n879) );
  NAND2_X1 U980 ( .A1(G112), .A2(n900), .ZN(n878) );
  NAND2_X1 U981 ( .A1(n879), .A2(n878), .ZN(n880) );
  NOR2_X1 U982 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U983 ( .A(KEYINPUT110), .B(n882), .ZN(G162) );
  NAND2_X1 U984 ( .A1(n518), .A2(G106), .ZN(n884) );
  NAND2_X1 U985 ( .A1(G142), .A2(n897), .ZN(n883) );
  NAND2_X1 U986 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U987 ( .A(n885), .B(KEYINPUT45), .ZN(n890) );
  NAND2_X1 U988 ( .A1(G130), .A2(n902), .ZN(n887) );
  NAND2_X1 U989 ( .A1(G118), .A2(n900), .ZN(n886) );
  NAND2_X1 U990 ( .A1(n887), .A2(n886), .ZN(n888) );
  XNOR2_X1 U991 ( .A(KEYINPUT111), .B(n888), .ZN(n889) );
  NAND2_X1 U992 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U993 ( .A(n891), .B(G162), .ZN(n895) );
  XNOR2_X1 U994 ( .A(n892), .B(KEYINPUT48), .ZN(n893) );
  XNOR2_X1 U995 ( .A(n893), .B(KEYINPUT46), .ZN(n894) );
  XNOR2_X1 U996 ( .A(n895), .B(n894), .ZN(n909) );
  NAND2_X1 U997 ( .A1(n518), .A2(G103), .ZN(n899) );
  NAND2_X1 U998 ( .A1(G139), .A2(n897), .ZN(n898) );
  NAND2_X1 U999 ( .A1(n899), .A2(n898), .ZN(n907) );
  NAND2_X1 U1000 ( .A1(n900), .A2(G115), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(n901), .B(KEYINPUT112), .ZN(n904) );
  NAND2_X1 U1002 ( .A1(G127), .A2(n902), .ZN(n903) );
  NAND2_X1 U1003 ( .A1(n904), .A2(n903), .ZN(n905) );
  XOR2_X1 U1004 ( .A(KEYINPUT47), .B(n905), .Z(n906) );
  NOR2_X1 U1005 ( .A1(n907), .A2(n906), .ZN(n1021) );
  XNOR2_X1 U1006 ( .A(G160), .B(n1021), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1008 ( .A(n910), .B(n1015), .Z(n913) );
  XOR2_X1 U1009 ( .A(G164), .B(n911), .Z(n912) );
  XNOR2_X1 U1010 ( .A(n913), .B(n912), .ZN(n915) );
  XNOR2_X1 U1011 ( .A(n915), .B(n914), .ZN(n916) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n916), .ZN(G395) );
  XNOR2_X1 U1013 ( .A(n917), .B(KEYINPUT113), .ZN(n920) );
  XNOR2_X1 U1014 ( .A(G171), .B(n918), .ZN(n919) );
  XNOR2_X1 U1015 ( .A(n920), .B(n919), .ZN(n921) );
  XNOR2_X1 U1016 ( .A(n921), .B(G286), .ZN(n922) );
  NOR2_X1 U1017 ( .A1(G37), .A2(n922), .ZN(G397) );
  NOR2_X1 U1018 ( .A1(G229), .A2(G227), .ZN(n923) );
  XOR2_X1 U1019 ( .A(KEYINPUT49), .B(n923), .Z(n924) );
  NAND2_X1 U1020 ( .A1(G319), .A2(n924), .ZN(n925) );
  NOR2_X1 U1021 ( .A1(G401), .A2(n925), .ZN(n926) );
  XNOR2_X1 U1022 ( .A(KEYINPUT114), .B(n926), .ZN(n928) );
  NOR2_X1 U1023 ( .A1(G395), .A2(G397), .ZN(n927) );
  NAND2_X1 U1024 ( .A1(n928), .A2(n927), .ZN(G225) );
  INV_X1 U1025 ( .A(G225), .ZN(G308) );
  INV_X1 U1026 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1027 ( .A(G16), .B(KEYINPUT56), .ZN(n955) );
  XOR2_X1 U1028 ( .A(G1966), .B(KEYINPUT122), .Z(n929) );
  XNOR2_X1 U1029 ( .A(G168), .B(n929), .ZN(n931) );
  NOR2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1031 ( .A(KEYINPUT57), .B(n932), .Z(n953) );
  XNOR2_X1 U1032 ( .A(G1348), .B(n933), .ZN(n936) );
  XNOR2_X1 U1033 ( .A(G1341), .B(n934), .ZN(n935) );
  NOR2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n943) );
  XNOR2_X1 U1035 ( .A(n937), .B(G1956), .ZN(n939) );
  NAND2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n941) );
  XNOR2_X1 U1037 ( .A(G1971), .B(G303), .ZN(n940) );
  NOR2_X1 U1038 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n950) );
  XNOR2_X1 U1040 ( .A(n944), .B(KEYINPUT123), .ZN(n948) );
  XNOR2_X1 U1041 ( .A(G1961), .B(G301), .ZN(n945) );
  NOR2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1045 ( .A(KEYINPUT124), .B(n951), .ZN(n952) );
  NAND2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1047 ( .A1(n955), .A2(n954), .ZN(n1036) );
  XOR2_X1 U1048 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n978) );
  XNOR2_X1 U1049 ( .A(G1966), .B(G21), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(G1961), .B(G5), .ZN(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n976) );
  XNOR2_X1 U1052 ( .A(G20), .B(n958), .ZN(n962) );
  XNOR2_X1 U1053 ( .A(G1341), .B(G19), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(G1981), .B(G6), .ZN(n959) );
  NOR2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n965) );
  XOR2_X1 U1057 ( .A(KEYINPUT59), .B(G1348), .Z(n963) );
  XNOR2_X1 U1058 ( .A(G4), .B(n963), .ZN(n964) );
  NOR2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1060 ( .A(KEYINPUT60), .B(n966), .Z(n974) );
  XOR2_X1 U1061 ( .A(G1986), .B(G24), .Z(n969) );
  XNOR2_X1 U1062 ( .A(n967), .B(G22), .ZN(n968) );
  NAND2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n971) );
  XNOR2_X1 U1064 ( .A(G23), .B(G1976), .ZN(n970) );
  NOR2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n972) );
  XOR2_X1 U1066 ( .A(KEYINPUT58), .B(n972), .Z(n973) );
  NOR2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1069 ( .A(n978), .B(n977), .ZN(n979) );
  XNOR2_X1 U1070 ( .A(n979), .B(KEYINPUT61), .ZN(n980) );
  NOR2_X1 U1071 ( .A1(G16), .A2(n980), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(KEYINPUT127), .B(n981), .ZN(n982) );
  NAND2_X1 U1073 ( .A1(n982), .A2(G11), .ZN(n1034) );
  XNOR2_X1 U1074 ( .A(n983), .B(G27), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(n984), .B(KEYINPUT119), .ZN(n988) );
  XNOR2_X1 U1076 ( .A(G1996), .B(G32), .ZN(n986) );
  XNOR2_X1 U1077 ( .A(G33), .B(G2072), .ZN(n985) );
  NOR2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n991) );
  XNOR2_X1 U1080 ( .A(KEYINPUT118), .B(G2067), .ZN(n989) );
  XNOR2_X1 U1081 ( .A(G26), .B(n989), .ZN(n990) );
  NOR2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1083 ( .A(KEYINPUT120), .B(n992), .ZN(n993) );
  NAND2_X1 U1084 ( .A1(n993), .A2(G28), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(G25), .B(G1991), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1087 ( .A(KEYINPUT53), .B(n996), .Z(n1000) );
  XNOR2_X1 U1088 ( .A(KEYINPUT54), .B(G34), .ZN(n997) );
  XNOR2_X1 U1089 ( .A(n997), .B(KEYINPUT121), .ZN(n998) );
  XNOR2_X1 U1090 ( .A(G2084), .B(n998), .ZN(n999) );
  NAND2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(G35), .B(G2090), .ZN(n1001) );
  NOR2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(G29), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1095 ( .A(KEYINPUT55), .B(KEYINPUT117), .Z(n1004) );
  XNOR2_X1 U1096 ( .A(n1005), .B(n1004), .ZN(n1032) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1012) );
  XOR2_X1 U1098 ( .A(G2090), .B(G162), .Z(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(n1010), .B(KEYINPUT51), .ZN(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1028) );
  XNOR2_X1 U1102 ( .A(G2084), .B(G160), .ZN(n1013) );
  XNOR2_X1 U1103 ( .A(KEYINPUT115), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(KEYINPUT116), .B(n1020), .ZN(n1026) );
  XOR2_X1 U1108 ( .A(G2072), .B(n1021), .Z(n1023) );
  XOR2_X1 U1109 ( .A(G164), .B(G2078), .Z(n1022) );
  NOR2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1111 ( .A(KEYINPUT50), .B(n1024), .Z(n1025) );
  NOR2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1114 ( .A(KEYINPUT52), .B(n1029), .ZN(n1030) );
  NAND2_X1 U1115 ( .A1(G29), .A2(n1030), .ZN(n1031) );
  NAND2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NOR2_X1 U1117 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1118 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XOR2_X1 U1119 ( .A(KEYINPUT62), .B(n1037), .Z(G311) );
  INV_X1 U1120 ( .A(G311), .ZN(G150) );
endmodule

