//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 0 1 1 0 1 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0 1 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND3_X1  g0009(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  AOI21_X1  g0011(.A(KEYINPUT64), .B1(G1), .B2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n209), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT65), .ZN(new_n219));
  XNOR2_X1  g0019(.A(KEYINPUT66), .B(G244), .ZN(new_n220));
  AND2_X1   g0020(.A1(new_n220), .A2(G77), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G107), .A2(G264), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n206), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT1), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n219), .A2(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT67), .ZN(new_n240));
  XOR2_X1   g0040(.A(G58), .B(G77), .Z(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  INV_X1    g0046(.A(G58), .ZN(new_n247));
  OAI21_X1  g0047(.A(KEYINPUT69), .B1(new_n247), .B2(KEYINPUT8), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT69), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT8), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n249), .A2(new_n250), .A3(G58), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n247), .A2(KEYINPUT8), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n248), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n214), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G1), .A2(G13), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT64), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n262), .A2(new_n210), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT70), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT68), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(KEYINPUT68), .A2(G1), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n269), .A2(G13), .A3(G20), .A4(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(G50), .ZN(new_n272));
  AND3_X1   g0072(.A1(new_n262), .A2(new_n210), .A3(new_n263), .ZN(new_n273));
  AND2_X1   g0073(.A1(KEYINPUT68), .A2(G1), .ZN(new_n274));
  NOR2_X1   g0074(.A1(KEYINPUT68), .A2(G1), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G20), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n272), .B1(new_n279), .B2(G50), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n266), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n265), .A2(KEYINPUT70), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT3), .B(G33), .ZN(new_n286));
  INV_X1    g0086(.A(G1698), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(G222), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(G223), .A3(G1698), .ZN(new_n289));
  INV_X1    g0089(.A(G77), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n288), .B(new_n289), .C1(new_n290), .C2(new_n286), .ZN(new_n291));
  AND2_X1   g0091(.A1(G33), .A2(G41), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n213), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(G274), .B1(new_n292), .B2(new_n260), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G41), .A2(G45), .ZN(new_n296));
  NOR3_X1   g0096(.A1(new_n295), .A2(G1), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n296), .ZN(new_n298));
  AND2_X1   g0098(.A1(G1), .A2(G13), .ZN(new_n299));
  NAND2_X1  g0099(.A1(G33), .A2(G41), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n276), .A2(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n297), .B1(G226), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n294), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G179), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n294), .A2(new_n302), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n285), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  OR3_X1    g0108(.A1(new_n281), .A2(KEYINPUT9), .A3(new_n283), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT9), .B1(new_n281), .B2(new_n283), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G190), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n303), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n313), .B1(G200), .B2(new_n303), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT10), .ZN(new_n315));
  AND3_X1   g0115(.A1(new_n311), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n315), .B1(new_n311), .B2(new_n314), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n308), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n271), .ZN(new_n320));
  INV_X1    g0120(.A(G68), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT12), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n320), .A2(KEYINPUT12), .A3(new_n321), .ZN(new_n323));
  AOI211_X1 g0123(.A(new_n322), .B(new_n323), .C1(G68), .C2(new_n279), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n257), .A2(G50), .ZN(new_n325));
  OAI221_X1 g0125(.A(new_n325), .B1(new_n214), .B2(G68), .C1(new_n290), .C2(new_n254), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n264), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n327), .B(KEYINPUT11), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT14), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n297), .B1(G238), .B2(new_n301), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n286), .A2(G232), .A3(G1698), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n286), .A2(G226), .A3(new_n287), .ZN(new_n333));
  NAND2_X1  g0133(.A1(G33), .A2(G97), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n293), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT13), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n331), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n337), .B1(new_n331), .B2(new_n336), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n330), .B(G169), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n331), .A2(new_n336), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT13), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n343), .A2(G179), .A3(new_n338), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n338), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n330), .B1(new_n346), .B2(G169), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n329), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n299), .A2(new_n300), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n269), .A2(new_n270), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n220), .B(new_n349), .C1(new_n350), .C2(new_n296), .ZN(new_n351));
  INV_X1    g0151(.A(G274), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(new_n299), .B2(new_n300), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n353), .A2(new_n268), .A3(new_n298), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT71), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT71), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n351), .A2(new_n357), .A3(new_n354), .ZN(new_n358));
  INV_X1    g0158(.A(G33), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(KEYINPUT3), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT3), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(G33), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n360), .A2(new_n362), .A3(G232), .A4(new_n287), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n360), .A2(new_n362), .A3(G238), .A4(G1698), .ZN(new_n364));
  INV_X1    g0164(.A(G107), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n363), .B(new_n364), .C1(new_n365), .C2(new_n286), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n293), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n356), .A2(new_n358), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT72), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n355), .A2(KEYINPUT71), .B1(new_n366), .B2(new_n293), .ZN(new_n371));
  AOI21_X1  g0171(.A(KEYINPUT72), .B1(new_n371), .B2(new_n358), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n306), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n368), .A2(new_n369), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n371), .A2(KEYINPUT72), .A3(new_n358), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n374), .A2(new_n304), .A3(new_n375), .ZN(new_n376));
  XNOR2_X1  g0176(.A(KEYINPUT15), .B(G87), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n255), .ZN(new_n379));
  OAI21_X1  g0179(.A(KEYINPUT74), .B1(new_n214), .B2(new_n290), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n257), .A2(KEYINPUT73), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n257), .A2(KEYINPUT73), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n250), .A2(G58), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n252), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n382), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT74), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n381), .B(new_n386), .C1(new_n387), .C2(new_n379), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n264), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n271), .A2(G77), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n279), .B2(G77), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n373), .A2(new_n376), .A3(new_n392), .ZN(new_n393));
  AND2_X1   g0193(.A1(new_n348), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT16), .ZN(new_n395));
  AND2_X1   g0195(.A1(G58), .A2(G68), .ZN(new_n396));
  OAI21_X1  g0196(.A(G20), .B1(new_n396), .B2(new_n201), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT75), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI211_X1 g0199(.A(KEYINPUT75), .B(G20), .C1(new_n396), .C2(new_n201), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n257), .A2(G159), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT7), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(new_n286), .B2(G20), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n360), .A2(new_n362), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n406), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n321), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n395), .B1(new_n403), .B2(new_n408), .ZN(new_n409));
  NOR3_X1   g0209(.A1(new_n286), .A2(new_n404), .A3(G20), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT7), .B1(new_n406), .B2(new_n214), .ZN(new_n411));
  OAI21_X1  g0211(.A(G68), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n399), .A2(new_n400), .B1(G159), .B2(new_n257), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(KEYINPUT16), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n409), .A2(new_n264), .A3(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n320), .A2(new_n253), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(new_n253), .B2(new_n278), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n349), .B1(new_n350), .B2(new_n296), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n354), .B1(new_n420), .B2(new_n231), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n286), .A2(G226), .A3(G1698), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n286), .A2(G223), .A3(new_n287), .ZN(new_n423));
  NAND2_X1  g0223(.A1(G33), .A2(G87), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT76), .ZN(new_n425));
  XNOR2_X1  g0225(.A(new_n424), .B(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n422), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n421), .B1(new_n293), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(G179), .ZN(new_n429));
  INV_X1    g0229(.A(new_n421), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n427), .A2(new_n293), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(G169), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n419), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT18), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT18), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n419), .A2(new_n434), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n430), .A2(new_n431), .A3(new_n312), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(new_n428), .B2(G200), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n440), .A2(new_n415), .A3(new_n418), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT17), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n440), .A2(new_n415), .A3(KEYINPUT17), .A4(new_n418), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n436), .A2(new_n438), .A3(new_n443), .A4(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(G190), .B1(new_n370), .B2(new_n372), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n374), .A2(G200), .A3(new_n375), .ZN(new_n448));
  INV_X1    g0248(.A(new_n392), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n346), .A2(new_n312), .ZN(new_n452));
  INV_X1    g0252(.A(G200), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n453), .B1(new_n343), .B2(new_n338), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n452), .A2(new_n329), .A3(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n319), .A2(new_n394), .A3(new_n446), .A4(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  AND3_X1   g0258(.A1(new_n365), .A2(KEYINPUT23), .A3(G20), .ZN(new_n459));
  AOI21_X1  g0259(.A(KEYINPUT23), .B1(new_n365), .B2(G20), .ZN(new_n460));
  INV_X1    g0260(.A(G116), .ZN(new_n461));
  OAI22_X1  g0261(.A1(new_n459), .A2(new_n460), .B1(new_n461), .B2(new_n254), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n360), .A2(new_n362), .A3(new_n214), .A4(G87), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT22), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT22), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n286), .A2(new_n465), .A3(new_n214), .A4(G87), .ZN(new_n466));
  AOI211_X1 g0266(.A(KEYINPUT24), .B(new_n462), .C1(new_n464), .C2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT24), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n464), .A2(new_n466), .ZN(new_n469));
  INV_X1    g0269(.A(new_n462), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n264), .B1(new_n467), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n269), .A2(G33), .A3(new_n270), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n273), .A2(new_n271), .A3(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(new_n365), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT25), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n476), .B1(new_n271), .B2(G107), .ZN(new_n477));
  NOR3_X1   g0277(.A1(new_n271), .A2(new_n476), .A3(G107), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT90), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(KEYINPUT90), .B(new_n476), .C1(new_n271), .C2(G107), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n475), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n472), .A2(KEYINPUT91), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(KEYINPUT91), .B1(new_n472), .B2(new_n482), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n360), .A2(new_n362), .A3(G257), .A4(G1698), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n360), .A2(new_n362), .A3(G250), .A4(new_n287), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G294), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n293), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT5), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT80), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n491), .B1(new_n492), .B2(G41), .ZN(new_n493));
  INV_X1    g0293(.A(G41), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n494), .A2(KEYINPUT80), .A3(KEYINPUT5), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n269), .A2(G45), .A3(new_n270), .ZN(new_n497));
  OAI211_X1 g0297(.A(G264), .B(new_n349), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(G45), .ZN(new_n499));
  NOR3_X1   g0299(.A1(new_n274), .A2(new_n275), .A3(new_n499), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n500), .A2(new_n353), .A3(new_n493), .A4(new_n495), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n490), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n502), .A2(new_n306), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(G169), .B2(new_n502), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n496), .A2(new_n349), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n497), .A2(new_n349), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n508), .A2(G264), .B1(new_n489), .B2(new_n293), .ZN(new_n509));
  AOI21_X1  g0309(.A(G200), .B1(new_n509), .B2(new_n501), .ZN(new_n510));
  AND4_X1   g0310(.A1(new_n312), .A2(new_n490), .A3(new_n498), .A4(new_n501), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n472), .B(new_n482), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT92), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n502), .A2(new_n453), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(G190), .B2(new_n502), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n516), .A2(KEYINPUT92), .A3(new_n472), .A4(new_n482), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n485), .A2(new_n505), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n360), .A2(new_n362), .A3(G264), .A4(G1698), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n360), .A2(new_n362), .A3(G257), .A4(new_n287), .ZN(new_n520));
  XOR2_X1   g0320(.A(KEYINPUT87), .B(G303), .Z(new_n521));
  OAI211_X1 g0321(.A(new_n519), .B(new_n520), .C1(new_n521), .C2(new_n286), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n293), .ZN(new_n523));
  OAI211_X1 g0323(.A(G270), .B(new_n349), .C1(new_n496), .C2(new_n497), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(new_n501), .A3(new_n524), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n273), .A2(G116), .A3(new_n271), .A4(new_n473), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n320), .A2(new_n461), .ZN(new_n527));
  AOI21_X1  g0327(.A(G20), .B1(G33), .B2(G283), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n359), .A2(G97), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n528), .A2(new_n529), .B1(G20), .B2(new_n461), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n530), .A2(new_n264), .A3(KEYINPUT20), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT20), .B1(new_n530), .B2(new_n264), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n526), .B(new_n527), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n525), .A2(G169), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(KEYINPUT88), .A2(KEYINPUT21), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n522), .A2(new_n293), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n524), .A2(new_n501), .ZN(new_n538));
  OAI21_X1  g0338(.A(G200), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n533), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n524), .A2(new_n501), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n541), .A2(G190), .A3(new_n523), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n533), .A2(G179), .A3(new_n523), .A4(new_n541), .ZN(new_n544));
  INV_X1    g0344(.A(new_n535), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n525), .A2(new_n533), .A3(G169), .A4(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n536), .A2(new_n543), .A3(new_n544), .A4(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT89), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n546), .A2(new_n544), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT89), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n549), .A2(new_n550), .A3(new_n536), .A4(new_n543), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n501), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n553), .B1(G257), .B2(new_n508), .ZN(new_n554));
  INV_X1    g0354(.A(G244), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n555), .A2(G1698), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n556), .A2(new_n360), .A3(new_n362), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT4), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT4), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n286), .A2(new_n559), .A3(new_n556), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n360), .A2(new_n362), .A3(G250), .A4(G1698), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G33), .A2(G283), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n561), .A2(KEYINPUT79), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n293), .ZN(new_n566));
  AOI21_X1  g0366(.A(KEYINPUT79), .B1(new_n561), .B2(new_n564), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n554), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(KEYINPUT82), .B1(new_n568), .B2(G179), .ZN(new_n569));
  XOR2_X1   g0369(.A(G97), .B(G107), .Z(new_n570));
  XNOR2_X1  g0370(.A(KEYINPUT77), .B(KEYINPUT6), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n571), .A2(KEYINPUT78), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n571), .A2(G97), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n570), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n570), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n571), .A2(KEYINPUT78), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n574), .A2(G20), .A3(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(G107), .B1(new_n410), .B2(new_n411), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n257), .A2(G77), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n264), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(G97), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n320), .A2(new_n583), .ZN(new_n584));
  OR2_X1    g0384(.A1(new_n474), .A2(new_n583), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n582), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n508), .A2(G257), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n501), .ZN(new_n588));
  INV_X1    g0388(.A(new_n293), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n562), .A2(new_n563), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n590), .B1(new_n558), .B2(new_n560), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n589), .B1(new_n591), .B2(KEYINPUT79), .ZN(new_n592));
  INV_X1    g0392(.A(new_n567), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n588), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT82), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n594), .A2(new_n595), .A3(new_n306), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n568), .A2(new_n304), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n569), .A2(new_n586), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n312), .B(new_n554), .C1(new_n566), .C2(new_n567), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n594), .B2(G200), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT81), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n585), .A2(new_n584), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n574), .A2(new_n577), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n580), .B(new_n579), .C1(new_n603), .C2(new_n214), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n602), .B1(new_n604), .B2(new_n264), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n600), .A2(new_n601), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n601), .B1(new_n600), .B2(new_n605), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n598), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT85), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT83), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n295), .B2(new_n497), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n500), .A2(KEYINPUT83), .A3(new_n353), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n276), .A2(G45), .B1(new_n299), .B2(new_n300), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n611), .A2(new_n612), .B1(new_n613), .B2(G250), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n360), .A2(new_n362), .A3(G244), .A4(G1698), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n360), .A2(new_n362), .A3(G238), .A4(new_n287), .ZN(new_n616));
  NAND2_X1  g0416(.A1(G33), .A2(G116), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n293), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n453), .B1(new_n614), .B2(new_n619), .ZN(new_n620));
  NOR3_X1   g0420(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n621));
  INV_X1    g0421(.A(new_n334), .ZN(new_n622));
  AND2_X1   g0422(.A1(KEYINPUT84), .A2(KEYINPUT19), .ZN(new_n623));
  NOR2_X1   g0423(.A1(KEYINPUT84), .A2(KEYINPUT19), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n621), .B1(new_n625), .B2(new_n214), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n360), .A2(new_n362), .A3(new_n214), .A4(G68), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n214), .A2(G33), .A3(G97), .ZN(new_n628));
  OR2_X1    g0428(.A1(KEYINPUT84), .A2(KEYINPUT19), .ZN(new_n629));
  NAND2_X1  g0429(.A1(KEYINPUT84), .A2(KEYINPUT19), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n264), .B1(new_n626), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n320), .A2(new_n377), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n273), .A2(G87), .A3(new_n271), .A4(new_n473), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n609), .B1(new_n620), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n497), .A2(G250), .A3(new_n349), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n295), .A2(new_n497), .A3(new_n610), .ZN(new_n639));
  AOI21_X1  g0439(.A(KEYINPUT83), .B1(new_n500), .B2(new_n353), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n618), .A2(new_n293), .ZN(new_n642));
  OAI21_X1  g0442(.A(G200), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(new_n644), .A3(KEYINPUT85), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n614), .A2(G190), .A3(new_n619), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n637), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n611), .A2(new_n612), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n648), .A2(new_n619), .A3(new_n638), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n304), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n633), .B(new_n634), .C1(new_n377), .C2(new_n474), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n650), .B(new_n651), .C1(G179), .C2(new_n649), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(KEYINPUT86), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT86), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n647), .A2(new_n655), .A3(new_n652), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n608), .A2(new_n657), .ZN(new_n658));
  AND4_X1   g0458(.A1(new_n458), .A2(new_n518), .A3(new_n552), .A4(new_n658), .ZN(G372));
  INV_X1    g0459(.A(KEYINPUT26), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n643), .A2(new_n644), .A3(new_n646), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n652), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n660), .B1(new_n598), .B2(new_n662), .ZN(new_n663));
  AND4_X1   g0463(.A1(new_n596), .A2(new_n569), .A3(new_n586), .A4(new_n597), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n654), .A2(new_n664), .A3(new_n656), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n663), .B1(new_n665), .B2(new_n660), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n600), .A2(new_n605), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT81), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n600), .A2(new_n601), .A3(new_n605), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n472), .A2(new_n482), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(new_n504), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n549), .A2(new_n536), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n662), .B1(new_n514), .B2(new_n517), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n670), .A2(new_n598), .A3(new_n674), .A4(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n666), .A2(new_n652), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n458), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n394), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n348), .A2(new_n455), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n679), .A2(new_n443), .A3(new_n444), .A4(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n436), .A2(new_n438), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n316), .A2(new_n317), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n678), .A2(new_n308), .A3(new_n687), .ZN(G369));
  AND2_X1   g0488(.A1(new_n214), .A2(G13), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n276), .A2(new_n689), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(G213), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(G343), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(new_n540), .ZN(new_n697));
  MUX2_X1   g0497(.A(new_n552), .B(new_n673), .S(new_n697), .Z(new_n698));
  AND2_X1   g0498(.A1(new_n698), .A2(G330), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n485), .A2(new_n505), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n695), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n485), .A2(new_n695), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n518), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n699), .A2(new_n705), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n706), .A2(KEYINPUT93), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(KEYINPUT93), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n673), .A2(new_n696), .ZN(new_n710));
  XOR2_X1   g0510(.A(new_n710), .B(KEYINPUT94), .Z(new_n711));
  AND2_X1   g0511(.A1(new_n711), .A2(new_n705), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n672), .A2(new_n696), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n709), .A2(new_n715), .ZN(G399));
  INV_X1    g0516(.A(new_n207), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(G41), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n621), .A2(new_n461), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n719), .A2(G1), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(new_n217), .B2(new_n719), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT28), .ZN(new_n723));
  OAI211_X1 g0523(.A(new_n675), .B(new_n598), .C1(new_n606), .C2(new_n607), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n673), .B1(new_n485), .B2(new_n505), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n652), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n598), .A2(new_n660), .A3(new_n662), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n727), .B1(new_n665), .B2(new_n660), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n696), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(KEYINPUT29), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT30), .ZN(new_n731));
  INV_X1    g0531(.A(new_n525), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n641), .A2(new_n642), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n732), .A2(new_n733), .A3(G179), .A4(new_n509), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n731), .B1(new_n734), .B2(new_n568), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n509), .A2(new_n619), .A3(new_n614), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n525), .A2(new_n306), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n594), .A2(KEYINPUT30), .A3(new_n736), .A4(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n732), .A2(G179), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n739), .A2(new_n568), .A3(new_n502), .A4(new_n649), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n735), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  AND3_X1   g0541(.A1(new_n741), .A2(KEYINPUT31), .A3(new_n695), .ZN(new_n742));
  AOI21_X1  g0542(.A(KEYINPUT31), .B1(new_n741), .B2(new_n695), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n670), .A2(new_n656), .A3(new_n654), .A4(new_n598), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n518), .A2(new_n552), .A3(new_n696), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G330), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT29), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n677), .A2(new_n749), .A3(new_n696), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n730), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n723), .B1(new_n752), .B2(G1), .ZN(G364));
  AOI21_X1  g0553(.A(new_n268), .B1(new_n689), .B2(G45), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n718), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n699), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n757), .B1(G330), .B2(new_n698), .ZN(new_n758));
  INV_X1    g0558(.A(new_n756), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n213), .B1(G20), .B2(new_n304), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n760), .A2(KEYINPUT96), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(KEYINPUT96), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n214), .A2(G179), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n765), .A2(G190), .A3(G200), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n767), .A2(KEYINPUT98), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(KEYINPUT98), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G303), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n406), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  XOR2_X1   g0572(.A(new_n772), .B(KEYINPUT99), .Z(new_n773));
  NOR2_X1   g0573(.A1(new_n214), .A2(new_n306), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G190), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G200), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G322), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n775), .A2(new_n453), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G326), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n777), .A2(new_n778), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n453), .A2(G190), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n774), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G317), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(KEYINPUT33), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n786), .A2(KEYINPUT33), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n785), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G283), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n765), .A2(new_n783), .ZN(new_n791));
  INV_X1    g0591(.A(G311), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G190), .A2(G200), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n774), .A2(new_n793), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n789), .B1(new_n790), .B2(new_n791), .C1(new_n792), .C2(new_n794), .ZN(new_n795));
  AND3_X1   g0595(.A1(new_n306), .A2(new_n453), .A3(KEYINPUT97), .ZN(new_n796));
  AOI21_X1  g0596(.A(KEYINPUT97), .B1(new_n306), .B2(new_n453), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR3_X1   g0598(.A1(new_n798), .A2(new_n214), .A3(G190), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n782), .B(new_n795), .C1(G329), .C2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G294), .ZN(new_n801));
  INV_X1    g0601(.A(new_n798), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n214), .B1(new_n802), .B2(G190), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n773), .B(new_n800), .C1(new_n801), .C2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n794), .ZN(new_n805));
  INV_X1    g0605(.A(new_n791), .ZN(new_n806));
  AOI22_X1  g0606(.A1(G77), .A2(new_n805), .B1(new_n806), .B2(G107), .ZN(new_n807));
  INV_X1    g0607(.A(G87), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n807), .B1(new_n808), .B2(new_n766), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n286), .B1(new_n321), .B2(new_n784), .C1(new_n780), .C2(new_n202), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n809), .B(new_n810), .C1(G58), .C2(new_n776), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n799), .A2(G159), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n812), .B(KEYINPUT32), .Z(new_n813));
  INV_X1    g0613(.A(new_n803), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G97), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n811), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n764), .B1(new_n804), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(G13), .A2(G33), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n214), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT95), .Z(new_n820));
  NAND2_X1  g0620(.A1(new_n764), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n286), .A2(G355), .A3(new_n207), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n242), .A2(new_n499), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n717), .A2(new_n286), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(G45), .B2(new_n217), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n823), .B1(G116), .B2(new_n207), .C1(new_n824), .C2(new_n826), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n759), .B(new_n817), .C1(new_n822), .C2(new_n827), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n820), .B(KEYINPUT100), .Z(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n828), .B1(new_n698), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n758), .A2(new_n831), .ZN(G396));
  NAND2_X1  g0632(.A1(new_n392), .A2(new_n695), .ZN(new_n833));
  AND3_X1   g0633(.A1(new_n393), .A2(KEYINPUT101), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n833), .B1(new_n393), .B2(KEYINPUT101), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n450), .B(new_n696), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n677), .A2(new_n837), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n677), .A2(new_n696), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n450), .B1(new_n834), .B2(new_n835), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n838), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n756), .B1(new_n842), .B2(new_n748), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n748), .B2(new_n842), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n763), .A2(new_n818), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n759), .B1(new_n845), .B2(new_n290), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n406), .B1(new_n806), .B2(G68), .ZN(new_n847));
  INV_X1    g0647(.A(new_n799), .ZN(new_n848));
  INV_X1    g0648(.A(G132), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n847), .B1(new_n848), .B2(new_n849), .C1(new_n770), .C2(new_n202), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(G58), .B2(new_n814), .ZN(new_n851));
  AOI22_X1  g0651(.A1(G150), .A2(new_n785), .B1(new_n805), .B2(G159), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n776), .A2(G143), .ZN(new_n853));
  INV_X1    g0653(.A(G137), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n852), .B(new_n853), .C1(new_n854), .C2(new_n780), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT34), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n770), .A2(new_n365), .B1(new_n848), .B2(new_n792), .ZN(new_n857));
  AOI22_X1  g0657(.A1(G116), .A2(new_n805), .B1(new_n806), .B2(G87), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n858), .B(new_n406), .C1(new_n790), .C2(new_n784), .ZN(new_n859));
  OAI22_X1  g0659(.A1(new_n777), .A2(new_n801), .B1(new_n780), .B2(new_n771), .ZN(new_n860));
  NOR3_X1   g0660(.A1(new_n857), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n851), .A2(new_n856), .B1(new_n815), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n818), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n846), .B1(new_n764), .B2(new_n862), .C1(new_n841), .C2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n844), .A2(new_n864), .ZN(G384));
  INV_X1    g0665(.A(KEYINPUT40), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n348), .A2(KEYINPUT102), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n696), .B1(new_n328), .B2(new_n324), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n455), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT102), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n870), .B(new_n329), .C1(new_n345), .C2(new_n347), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n867), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n345), .A2(new_n347), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n868), .B1(new_n873), .B2(new_n455), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n840), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n747), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n414), .A2(new_n264), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT103), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(new_n403), .B2(new_n408), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n412), .A2(KEYINPUT103), .A3(new_n413), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n879), .A2(new_n395), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n417), .B1(new_n877), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n434), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n441), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n882), .A2(new_n693), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT37), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n693), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n419), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT37), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n435), .A2(new_n888), .A3(new_n889), .A4(new_n441), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n445), .A2(new_n885), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n891), .A2(new_n892), .A3(KEYINPUT38), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT38), .B1(new_n891), .B2(new_n892), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n866), .B1(new_n876), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT105), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n875), .B(new_n747), .C1(new_n893), .C2(new_n894), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n899), .A2(KEYINPUT105), .A3(new_n866), .ZN(new_n900));
  INV_X1    g0700(.A(new_n876), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT38), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n435), .A2(new_n888), .A3(new_n441), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT104), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n903), .A2(new_n904), .A3(KEYINPUT37), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n446), .B2(new_n888), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n903), .A2(KEYINPUT37), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n907), .A2(KEYINPUT104), .A3(new_n890), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n902), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n891), .A2(new_n892), .A3(KEYINPUT38), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n866), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n898), .A2(new_n900), .B1(new_n901), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n458), .A2(new_n747), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT106), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n913), .A2(new_n915), .ZN(new_n917));
  INV_X1    g0717(.A(G330), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n872), .A2(new_n874), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n393), .A2(new_n695), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n921), .B1(new_n838), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n893), .B2(new_n894), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT39), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n903), .A2(KEYINPUT37), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n890), .A2(KEYINPUT104), .ZN(new_n927));
  INV_X1    g0727(.A(new_n888), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n926), .A2(new_n927), .B1(new_n445), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT38), .B1(new_n929), .B2(new_n908), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n925), .B1(new_n930), .B2(new_n893), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n867), .A2(new_n871), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n696), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n894), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n935), .A2(new_n911), .A3(KEYINPUT39), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n931), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n682), .A2(new_n693), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n924), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n457), .B1(new_n730), .B2(new_n750), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n687), .A2(new_n308), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n939), .B(new_n942), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n919), .A2(new_n943), .B1(new_n276), .B2(new_n689), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n943), .B2(new_n919), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT35), .ZN(new_n946));
  OAI211_X1 g0746(.A(G116), .B(new_n215), .C1(new_n603), .C2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(new_n946), .B2(new_n603), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT36), .ZN(new_n949));
  OR3_X1    g0749(.A1(new_n217), .A2(new_n396), .A3(new_n290), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n202), .A2(G68), .ZN(new_n951));
  AOI211_X1 g0751(.A(G13), .B(new_n276), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  OR3_X1    g0752(.A1(new_n945), .A2(new_n949), .A3(new_n952), .ZN(G367));
  INV_X1    g0753(.A(new_n608), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n586), .A2(new_n695), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n664), .A2(new_n695), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n712), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT42), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n959), .B(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n954), .A2(new_n701), .A3(new_n955), .ZN(new_n962));
  AOI21_X1  g0762(.A(KEYINPUT107), .B1(new_n962), .B2(new_n598), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n962), .A2(KEYINPUT107), .A3(new_n598), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n964), .A2(new_n696), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n961), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n696), .A2(new_n644), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n969), .A2(new_n652), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n969), .A2(new_n652), .A3(new_n661), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT43), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n967), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n975), .B1(new_n967), .B2(new_n976), .ZN(new_n979));
  INV_X1    g0779(.A(new_n958), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n978), .A2(new_n979), .B1(new_n709), .B2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n979), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n709), .A2(new_n980), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n982), .A2(new_n983), .A3(new_n977), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n718), .B(KEYINPUT41), .Z(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n699), .A2(KEYINPUT109), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n711), .B(new_n705), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n988), .B(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n752), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n715), .A2(new_n958), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(KEYINPUT45), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT108), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT44), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n994), .B(new_n995), .C1(new_n715), .C2(new_n958), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT45), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n715), .A2(new_n997), .A3(new_n958), .ZN(new_n998));
  AND3_X1   g0798(.A1(new_n993), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n709), .A2(KEYINPUT110), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n995), .B1(new_n715), .B2(new_n958), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n980), .B(KEYINPUT44), .C1(new_n712), .C2(new_n714), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1001), .A2(KEYINPUT108), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT110), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n707), .A2(new_n1004), .A3(new_n708), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n999), .A2(new_n1000), .A3(new_n1003), .A4(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1003), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n993), .A2(new_n996), .A3(new_n998), .ZN(new_n1008));
  OAI211_X1 g0808(.A(KEYINPUT110), .B(new_n709), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n991), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n987), .B1(new_n1010), .B2(new_n751), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n985), .B1(new_n1011), .B2(new_n754), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n791), .A2(new_n290), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1013), .A2(new_n406), .ZN(new_n1014));
  INV_X1    g0814(.A(G150), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1014), .B1(new_n1015), .B2(new_n777), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G58), .A2(new_n767), .B1(new_n785), .B2(G159), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(KEYINPUT112), .B(G137), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1017), .B1(new_n202), .B2(new_n794), .C1(new_n848), .C2(new_n1018), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n1016), .B(new_n1019), .C1(G143), .C2(new_n779), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n321), .B2(new_n803), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n770), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1022), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n799), .A2(G317), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n286), .B1(new_n806), .B2(G97), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G283), .A2(new_n805), .B1(new_n785), .B2(G294), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(KEYINPUT46), .B1(new_n767), .B2(G116), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G311), .B2(new_n779), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n521), .B2(new_n777), .C1(new_n803), .C2(new_n365), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1021), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT113), .Z(new_n1032));
  OR2_X1    g0832(.A1(new_n1032), .A2(KEYINPUT47), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(KEYINPUT47), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1033), .A2(new_n763), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n973), .A2(new_n829), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n825), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n237), .A2(new_n1037), .B1(new_n207), .B2(new_n377), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n756), .B1(new_n821), .B2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT111), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1035), .A2(new_n1036), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1012), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(G387));
  NAND3_X1  g0844(.A1(new_n702), .A2(new_n704), .A3(new_n829), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n286), .A2(new_n207), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n1046), .A2(new_n720), .B1(G107), .B2(new_n207), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n234), .A2(new_n499), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n720), .B(new_n499), .C1(new_n321), .C2(new_n290), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n385), .ZN(new_n1050));
  XOR2_X1   g0850(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n1051));
  NOR3_X1   g0851(.A1(new_n1050), .A2(new_n1051), .A3(G50), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1051), .B1(new_n1050), .B2(G50), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1037), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1047), .B1(new_n1048), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n756), .B1(new_n1056), .B2(new_n821), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n290), .A2(new_n766), .B1(new_n794), .B2(new_n321), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n406), .B(new_n1058), .C1(G97), .C2(new_n806), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n814), .A2(new_n378), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G50), .A2(new_n776), .B1(new_n779), .B2(G159), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n799), .A2(G150), .B1(new_n253), .B2(new_n785), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n286), .B1(new_n806), .B2(G116), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n803), .A2(new_n790), .B1(new_n801), .B2(new_n766), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n521), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1066), .A2(new_n805), .B1(new_n785), .B2(G311), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1067), .B1(new_n777), .B2(new_n786), .C1(new_n778), .C2(new_n780), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT48), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1065), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n1069), .B2(new_n1068), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT49), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1064), .B1(new_n781), .B2(new_n848), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1063), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1057), .B1(new_n1075), .B2(new_n763), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n990), .A2(new_n755), .B1(new_n1045), .B2(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n718), .B(KEYINPUT115), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n991), .A2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n990), .A2(new_n752), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1077), .B1(new_n1079), .B2(new_n1080), .ZN(G393));
  NAND2_X1  g0881(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n991), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1006), .A2(new_n1009), .A3(new_n991), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1084), .A2(new_n1078), .A3(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n958), .A2(new_n820), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT116), .Z(new_n1088));
  AOI22_X1  g0888(.A1(new_n245), .A2(new_n825), .B1(G97), .B2(new_n717), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n822), .A2(new_n1089), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G150), .A2(new_n779), .B1(new_n776), .B2(G159), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(KEYINPUT117), .B(KEYINPUT51), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1091), .B(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n290), .B2(new_n803), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n799), .A2(G143), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n406), .B1(new_n806), .B2(G87), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n767), .A2(G68), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n385), .A2(new_n805), .B1(new_n785), .B2(G50), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n406), .B1(new_n791), .B2(new_n365), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n521), .A2(new_n784), .B1(new_n794), .B2(new_n801), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n1100), .B(new_n1101), .C1(G283), .C2(new_n767), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1102), .B1(new_n461), .B2(new_n803), .C1(new_n778), .C2(new_n848), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(G311), .A2(new_n776), .B1(new_n779), .B2(G317), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT52), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n1094), .A2(new_n1099), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n759), .B(new_n1090), .C1(new_n763), .C2(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1082), .A2(new_n755), .B1(new_n1088), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1086), .A2(new_n1108), .ZN(G390));
  AOI21_X1  g0909(.A(new_n934), .B1(new_n910), .B2(new_n911), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n841), .B(new_n696), .C1(new_n726), .C2(new_n728), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n922), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1110), .B1(new_n1113), .B2(new_n921), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n931), .A2(new_n936), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n923), .B2(new_n934), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n747), .A2(G330), .A3(new_n841), .A4(new_n920), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n1114), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1117), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n755), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n845), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n766), .A2(new_n1015), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1123), .B(new_n1124), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(G128), .A2(new_n779), .B1(new_n776), .B2(G132), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(KEYINPUT54), .B(G143), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n794), .A2(new_n1127), .B1(new_n791), .B2(new_n202), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n286), .B1(new_n784), .B2(new_n1018), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1126), .A2(new_n1130), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1125), .B(new_n1131), .C1(G125), .C2(new_n799), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n814), .A2(G159), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n803), .A2(new_n290), .B1(new_n461), .B2(new_n777), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT120), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n770), .A2(new_n808), .B1(new_n848), .B2(new_n801), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(G97), .A2(new_n805), .B1(new_n785), .B2(G107), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n286), .B1(new_n806), .B2(G68), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1137), .B(new_n1138), .C1(new_n790), .C2(new_n780), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1132), .A2(new_n1133), .B1(new_n1135), .B2(new_n1140), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n756), .B1(new_n253), .B2(new_n1122), .C1(new_n1141), .C2(new_n764), .ZN(new_n1142));
  XOR2_X1   g0942(.A(new_n1142), .B(KEYINPUT121), .Z(new_n1143));
  INV_X1    g0943(.A(new_n1115), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1143), .B1(new_n1144), .B2(new_n863), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1119), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1114), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n838), .A2(new_n922), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n518), .A2(new_n552), .A3(new_n696), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n658), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n918), .B1(new_n1151), .B2(new_n744), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n920), .B1(new_n1152), .B2(new_n841), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1117), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1149), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n747), .A2(G330), .A3(new_n841), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n921), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1157), .A2(new_n922), .A3(new_n1111), .A4(new_n1117), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1155), .A2(KEYINPUT118), .A3(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n748), .A2(new_n457), .ZN(new_n1160));
  NOR3_X1   g0960(.A1(new_n940), .A2(new_n941), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT118), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1113), .A2(new_n1162), .A3(new_n1117), .A4(new_n1157), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1159), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1078), .B1(new_n1148), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1164), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1120), .A2(new_n1166), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1121), .B(new_n1145), .C1(new_n1165), .C2(new_n1167), .ZN(G378));
  INV_X1    g0968(.A(KEYINPUT122), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n285), .A2(new_n887), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n318), .A2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n308), .B(new_n1170), .C1(new_n316), .C2(new_n317), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1174), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1169), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1174), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(KEYINPUT122), .A3(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1177), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n918), .B1(new_n901), .B2(new_n912), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n899), .A2(KEYINPUT105), .A3(new_n866), .ZN(new_n1185));
  AOI21_X1  g0985(.A(KEYINPUT105), .B1(new_n899), .B2(new_n866), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1183), .B(new_n1184), .C1(new_n1185), .C2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(KEYINPUT40), .B1(new_n930), .B2(new_n893), .ZN(new_n1188));
  OAI21_X1  g0988(.A(G330), .B1(new_n1188), .B2(new_n876), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n898), .B2(new_n900), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1187), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n939), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1187), .B(new_n939), .C1(new_n1190), .C2(new_n1191), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1161), .B1(new_n1148), .B2(new_n1164), .ZN(new_n1197));
  AOI21_X1  g0997(.A(KEYINPUT57), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1194), .A2(KEYINPUT57), .A3(new_n1195), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1161), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1159), .A2(new_n1163), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1200), .B1(new_n1120), .B2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1078), .B1(new_n1199), .B2(new_n1203), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1198), .A2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n756), .B1(new_n1122), .B2(G50), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n286), .A2(G41), .ZN(new_n1207));
  AOI211_X1 g1007(.A(G50), .B(new_n1207), .C1(new_n359), .C2(new_n494), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1207), .B1(new_n290), .B2(new_n766), .C1(new_n780), .C2(new_n461), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(G107), .B2(new_n776), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n791), .A2(new_n247), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(G97), .B2(new_n785), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n377), .B2(new_n794), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G283), .B2(new_n799), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1210), .B(new_n1214), .C1(new_n321), .C2(new_n803), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT58), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1208), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n785), .A2(G132), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1218), .B1(new_n794), .B2(new_n854), .C1(new_n766), .C2(new_n1127), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(G125), .A2(new_n779), .B1(new_n776), .B2(G128), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1220), .B(new_n1221), .C1(new_n1015), .C2(new_n803), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1222), .A2(KEYINPUT59), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(KEYINPUT59), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n799), .A2(G124), .ZN(new_n1225));
  AOI211_X1 g1025(.A(G33), .B(G41), .C1(new_n806), .C2(G159), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1217), .B1(new_n1216), .B2(new_n1215), .C1(new_n1223), .C2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1206), .B1(new_n1228), .B2(new_n763), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n1183), .B2(new_n863), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n1196), .B2(new_n755), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1205), .A2(new_n1232), .ZN(G375));
  NAND2_X1  g1033(.A1(new_n921), .A2(new_n818), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(KEYINPUT123), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n849), .A2(new_n780), .B1(new_n777), .B2(new_n1018), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n1015), .A2(new_n794), .B1(new_n784), .B2(new_n1127), .ZN(new_n1237));
  NOR4_X1   g1037(.A1(new_n1236), .A2(new_n1237), .A3(new_n406), .A4(new_n1211), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1022), .A2(G159), .B1(G128), .B2(new_n799), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1238), .B(new_n1239), .C1(new_n202), .C2(new_n803), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n777), .A2(new_n790), .B1(new_n780), .B2(new_n801), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n365), .A2(new_n794), .B1(new_n784), .B2(new_n461), .ZN(new_n1242));
  NOR4_X1   g1042(.A1(new_n1241), .A2(new_n1242), .A3(new_n286), .A4(new_n1013), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1022), .A2(G97), .B1(G303), .B2(new_n799), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1243), .A2(new_n1244), .A3(new_n1060), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n764), .B1(new_n1240), .B2(new_n1245), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n759), .B(new_n1246), .C1(new_n321), .C2(new_n845), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1202), .A2(new_n755), .B1(new_n1235), .B2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1201), .A2(new_n1200), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1249), .A2(new_n987), .A3(new_n1164), .ZN(new_n1250));
  AND2_X1   g1050(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(G381));
  OR2_X1    g1052(.A1(G393), .A2(G396), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(G390), .A2(G384), .A3(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1145), .B1(new_n1148), .B2(new_n754), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1078), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(new_n1120), .B2(new_n1166), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1148), .A2(new_n1164), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1255), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1254), .A2(new_n1043), .A3(new_n1259), .A4(new_n1251), .ZN(new_n1260));
  OR2_X1    g1060(.A1(new_n1260), .A2(G375), .ZN(G407));
  NOR2_X1   g1061(.A1(new_n1260), .A2(G375), .ZN(new_n1262));
  INV_X1    g1062(.A(G213), .ZN(new_n1263));
  OR3_X1    g1063(.A1(new_n1263), .A2(KEYINPUT124), .A3(G343), .ZN(new_n1264));
  OAI21_X1  g1064(.A(KEYINPUT124), .B1(new_n1263), .B2(G343), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1266), .B(KEYINPUT125), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(G375), .A2(G378), .A3(new_n1267), .ZN(new_n1268));
  OR4_X1    g1068(.A1(KEYINPUT126), .A2(new_n1262), .A3(new_n1263), .A4(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(G407), .A2(G213), .ZN(new_n1270));
  OAI21_X1  g1070(.A(KEYINPUT126), .B1(new_n1270), .B2(new_n1268), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1269), .A2(new_n1271), .ZN(G409));
  INV_X1    g1072(.A(KEYINPUT61), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1267), .ZN(new_n1274));
  OAI211_X1 g1074(.A(G378), .B(new_n1232), .C1(new_n1198), .C2(new_n1204), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1276));
  NOR3_X1   g1076(.A1(new_n1203), .A2(new_n1276), .A3(new_n986), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1230), .B1(new_n1276), .B2(new_n754), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1259), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1274), .B1(new_n1275), .B2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(G2897), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1267), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT60), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1249), .A2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1161), .B1(new_n1159), .B2(new_n1163), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(KEYINPUT60), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1284), .A2(new_n1078), .A3(new_n1164), .A4(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(G384), .B1(new_n1287), .B2(new_n1248), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1078), .B(new_n1164), .C1(new_n1285), .C2(KEYINPUT60), .ZN(new_n1289));
  AOI211_X1 g1089(.A(new_n1283), .B(new_n1161), .C1(new_n1159), .C2(new_n1163), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1248), .B(G384), .C1(new_n1289), .C2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1282), .B1(new_n1288), .B2(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1248), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1294));
  INV_X1    g1094(.A(G384), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n1296), .B(new_n1291), .C1(new_n1281), .C2(new_n1266), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1293), .A2(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1273), .B1(new_n1280), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(KEYINPUT127), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1275), .A2(new_n1279), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1296), .A2(new_n1291), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1301), .A2(KEYINPUT62), .A3(new_n1267), .A4(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1266), .ZN(new_n1305));
  AOI211_X1 g1105(.A(new_n1305), .B(new_n1302), .C1(new_n1275), .C2(new_n1279), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1304), .B1(new_n1306), .B2(KEYINPUT62), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT127), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1308), .B(new_n1273), .C1(new_n1280), .C2(new_n1298), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1300), .A2(new_n1307), .A3(new_n1309), .ZN(new_n1310));
  AND2_X1   g1110(.A1(new_n1011), .A2(new_n754), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1041), .B(G390), .C1(new_n1311), .C2(new_n985), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1086), .B(new_n1108), .C1(new_n1012), .C2(new_n1042), .ZN(new_n1313));
  XOR2_X1   g1113(.A(G393), .B(G396), .Z(new_n1314));
  AND3_X1   g1114(.A1(new_n1312), .A2(new_n1313), .A3(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1314), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1316));
  OR2_X1    g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1310), .A2(new_n1317), .ZN(new_n1318));
  NOR3_X1   g1118(.A1(new_n1315), .A2(new_n1316), .A3(KEYINPUT61), .ZN(new_n1319));
  OR2_X1    g1119(.A1(new_n1306), .A2(KEYINPUT63), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1280), .A2(KEYINPUT63), .A3(new_n1303), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1301), .A2(new_n1266), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1322), .A2(new_n1297), .A3(new_n1293), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1319), .A2(new_n1320), .A3(new_n1321), .A4(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1318), .A2(new_n1324), .ZN(G405));
  AOI21_X1  g1125(.A(G378), .B1(new_n1205), .B2(new_n1232), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1275), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(new_n1302), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1303), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  XNOR2_X1  g1131(.A(new_n1331), .B(new_n1317), .ZN(G402));
endmodule


