//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 1 1 1 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n801, new_n802, new_n803, new_n804, new_n806, new_n807,
    new_n808, new_n809, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938;
  NOR2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203));
  AOI21_X1  g002(.A(new_n202), .B1(KEYINPUT23), .B2(new_n203), .ZN(new_n204));
  AND2_X1   g003(.A1(new_n202), .A2(KEYINPUT23), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207));
  XOR2_X1   g006(.A(new_n207), .B(KEYINPUT24), .Z(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G183gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n209), .A2(G190gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n206), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n207), .B(KEYINPUT24), .ZN(new_n212));
  INV_X1    g011(.A(G183gat), .ZN(new_n213));
  INV_X1    g012(.A(G190gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(KEYINPUT25), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  AOI22_X1  g015(.A1(new_n211), .A2(KEYINPUT25), .B1(new_n206), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n209), .A2(KEYINPUT27), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT27), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(new_n213), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT28), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(new_n222), .A3(new_n214), .ZN(new_n223));
  XOR2_X1   g022(.A(KEYINPUT27), .B(G183gat), .Z(new_n224));
  OAI21_X1  g023(.A(KEYINPUT28), .B1(new_n224), .B2(G190gat), .ZN(new_n225));
  INV_X1    g024(.A(G169gat), .ZN(new_n226));
  INV_X1    g025(.A(G176gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT26), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT26), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n202), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n203), .A3(new_n231), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n232), .A2(new_n207), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n223), .A2(new_n225), .A3(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G113gat), .B(G120gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n235), .A2(KEYINPUT1), .ZN(new_n236));
  XNOR2_X1  g035(.A(G127gat), .B(G134gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n237), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n239), .B1(KEYINPUT1), .B2(new_n235), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n217), .A2(new_n234), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT65), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n217), .A2(new_n234), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(new_n241), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT65), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n217), .A2(new_n234), .A3(new_n247), .A4(new_n242), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n244), .A2(new_n246), .A3(new_n248), .ZN(new_n249));
  AND2_X1   g048(.A1(G227gat), .A2(G233gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(KEYINPUT32), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT34), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT34), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n251), .A2(KEYINPUT32), .A3(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n249), .A2(new_n250), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n253), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n254), .B1(new_n251), .B2(KEYINPUT32), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT32), .ZN(new_n260));
  AOI211_X1 g059(.A(new_n260), .B(KEYINPUT34), .C1(new_n249), .C2(new_n250), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n256), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT33), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n251), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G15gat), .B(G43gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(G71gat), .B(G99gat), .ZN(new_n266));
  XOR2_X1   g065(.A(new_n265), .B(new_n266), .Z(new_n267));
  NAND2_X1  g066(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n258), .A2(new_n262), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n269), .B1(new_n258), .B2(new_n262), .ZN(new_n271));
  INV_X1    g070(.A(G228gat), .ZN(new_n272));
  INV_X1    g071(.A(G233gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G211gat), .B(G218gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n275), .B(KEYINPUT66), .ZN(new_n276));
  AND2_X1   g075(.A1(G211gat), .A2(G218gat), .ZN(new_n277));
  OR2_X1    g076(.A1(new_n277), .A2(KEYINPUT22), .ZN(new_n278));
  XNOR2_X1  g077(.A(G197gat), .B(G204gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT29), .ZN(new_n282));
  OR2_X1    g081(.A1(new_n275), .A2(KEYINPUT66), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n275), .A2(KEYINPUT66), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n283), .A2(new_n278), .A3(new_n279), .A4(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n281), .A2(new_n282), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT3), .ZN(new_n287));
  XOR2_X1   g086(.A(G141gat), .B(G148gat), .Z(new_n288));
  INV_X1    g087(.A(G155gat), .ZN(new_n289));
  INV_X1    g088(.A(G162gat), .ZN(new_n290));
  OAI21_X1  g089(.A(KEYINPUT2), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G155gat), .B(G162gat), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n288), .A2(new_n291), .A3(new_n293), .ZN(new_n296));
  AOI22_X1  g095(.A1(new_n286), .A2(new_n287), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n295), .A2(new_n287), .A3(new_n296), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(new_n282), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n281), .A2(new_n285), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n274), .B1(new_n298), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n302), .ZN(new_n304));
  INV_X1    g103(.A(new_n274), .ZN(new_n305));
  NOR3_X1   g104(.A1(new_n304), .A2(new_n297), .A3(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(G22gat), .B1(new_n303), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n298), .A2(new_n274), .A3(new_n302), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n305), .B1(new_n304), .B2(new_n297), .ZN(new_n309));
  INV_X1    g108(.A(G22gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G78gat), .B(G106gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(KEYINPUT31), .B(G50gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n313), .B(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT70), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n307), .A2(new_n311), .A3(new_n318), .ZN(new_n319));
  OR2_X1    g118(.A1(new_n307), .A2(KEYINPUT70), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n316), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NOR3_X1   g120(.A1(new_n270), .A2(new_n271), .A3(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G1gat), .B(G29gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n323), .B(G85gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT0), .B(G57gat), .ZN(new_n325));
  XOR2_X1   g124(.A(new_n324), .B(new_n325), .Z(new_n326));
  NAND2_X1  g125(.A1(new_n295), .A2(new_n296), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(new_n241), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n295), .A2(new_n238), .A3(new_n296), .A4(new_n240), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(KEYINPUT69), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G225gat), .A2(G233gat), .ZN(new_n331));
  XOR2_X1   g130(.A(new_n331), .B(KEYINPUT68), .Z(new_n332));
  INV_X1    g131(.A(KEYINPUT69), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n327), .A2(new_n333), .A3(new_n241), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n330), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n327), .A2(KEYINPUT3), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n336), .A2(new_n241), .A3(new_n299), .ZN(new_n337));
  AND2_X1   g136(.A1(new_n329), .A2(KEYINPUT4), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n329), .A2(KEYINPUT4), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n329), .A2(new_n332), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n335), .B(KEYINPUT5), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  OR2_X1    g141(.A1(new_n332), .A2(KEYINPUT5), .ZN(new_n343));
  OR2_X1    g142(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n326), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT6), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n342), .A2(new_n344), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT71), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT71), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n342), .A2(new_n344), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n326), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT6), .ZN(new_n352));
  INV_X1    g151(.A(new_n326), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n352), .B1(new_n347), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n346), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G8gat), .B(G36gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(G64gat), .B(G92gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  AND2_X1   g157(.A1(G226gat), .A2(G233gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n245), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT29), .B1(new_n217), .B2(new_n234), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n360), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n301), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n360), .B(new_n301), .C1(new_n359), .C2(new_n361), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n358), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT30), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n364), .A2(new_n358), .A3(new_n365), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT67), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n364), .A2(new_n365), .ZN(new_n370));
  INV_X1    g169(.A(new_n358), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT30), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n369), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n366), .A2(KEYINPUT67), .A3(KEYINPUT30), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n367), .B(new_n368), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n376), .A2(KEYINPUT35), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n322), .A2(KEYINPUT73), .A3(new_n355), .A4(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n354), .B(new_n345), .ZN(new_n379));
  INV_X1    g178(.A(new_n375), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT67), .B1(new_n366), .B2(KEYINPUT30), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n379), .A2(new_n382), .A3(new_n367), .A4(new_n368), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n257), .B1(new_n253), .B2(new_n255), .ZN(new_n384));
  NOR3_X1   g183(.A1(new_n259), .A2(new_n261), .A3(new_n256), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n268), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AND3_X1   g185(.A1(new_n316), .A2(new_n319), .A3(new_n320), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n258), .A2(new_n262), .A3(new_n269), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT35), .B1(new_n383), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT73), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n386), .A2(new_n387), .A3(new_n355), .A4(new_n388), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT35), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n382), .A2(new_n393), .A3(new_n367), .A4(new_n368), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n391), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n390), .A3(new_n395), .ZN(new_n396));
  AND3_X1   g195(.A1(new_n342), .A2(new_n344), .A3(new_n349), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n349), .B1(new_n342), .B2(new_n344), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n353), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n354), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n399), .A2(new_n400), .B1(KEYINPUT6), .B2(new_n345), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n370), .A2(KEYINPUT72), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT37), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT38), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT37), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n370), .A2(KEYINPUT72), .A3(new_n405), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n403), .A2(new_n404), .A3(new_n358), .A4(new_n406), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n403), .A2(new_n358), .A3(new_n406), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n366), .A2(KEYINPUT38), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n401), .B(new_n407), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n340), .A2(new_n332), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n411), .A2(KEYINPUT39), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n412), .A2(new_n353), .ZN(new_n413));
  AND2_X1   g212(.A1(new_n330), .A2(new_n334), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n411), .B(KEYINPUT39), .C1(new_n332), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT40), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT40), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n413), .A2(new_n418), .A3(new_n415), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n351), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n376), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n410), .A2(new_n421), .A3(new_n387), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n383), .A2(new_n321), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n386), .A2(KEYINPUT36), .A3(new_n388), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT36), .B1(new_n386), .B2(new_n388), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n422), .B(new_n423), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n396), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(G231gat), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n428), .A2(new_n273), .ZN(new_n429));
  NAND2_X1  g228(.A1(G71gat), .A2(G78gat), .ZN(new_n430));
  NOR2_X1   g229(.A1(G71gat), .A2(G78gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n431), .B(KEYINPUT82), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(KEYINPUT83), .ZN(new_n434));
  XNOR2_X1  g233(.A(G57gat), .B(G64gat), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n430), .B(new_n432), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT83), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n433), .B(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT84), .ZN(new_n439));
  INV_X1    g238(.A(G57gat), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n439), .B1(new_n440), .B2(G64gat), .ZN(new_n441));
  INV_X1    g240(.A(G64gat), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n442), .A2(KEYINPUT84), .A3(G57gat), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n441), .B(new_n443), .C1(G57gat), .C2(new_n442), .ZN(new_n444));
  INV_X1    g243(.A(new_n430), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n438), .B(new_n444), .C1(new_n445), .C2(new_n431), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n436), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n447), .A2(KEYINPUT21), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(KEYINPUT21), .ZN(new_n449));
  XNOR2_X1  g248(.A(G15gat), .B(G22gat), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT16), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n450), .B1(new_n451), .B2(G1gat), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n452), .B1(G1gat), .B2(new_n450), .ZN(new_n453));
  INV_X1    g252(.A(G8gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n453), .B(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT85), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n449), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n456), .B1(new_n449), .B2(new_n455), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n448), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n459), .ZN(new_n461));
  INV_X1    g260(.A(new_n448), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n457), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n429), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n460), .A2(new_n463), .A3(new_n429), .ZN(new_n466));
  XNOR2_X1  g265(.A(G183gat), .B(G211gat), .ZN(new_n467));
  XOR2_X1   g266(.A(new_n467), .B(G127gat), .Z(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n465), .A2(new_n466), .A3(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n471), .B(G155gat), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n460), .A2(new_n463), .A3(new_n429), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n468), .B1(new_n473), .B2(new_n464), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n470), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n472), .B1(new_n470), .B2(new_n474), .ZN(new_n476));
  OR2_X1    g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(KEYINPUT86), .B(G134gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(new_n290), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  XOR2_X1   g280(.A(KEYINPUT80), .B(KEYINPUT17), .Z(new_n482));
  INV_X1    g281(.A(KEYINPUT15), .ZN(new_n483));
  INV_X1    g282(.A(G43gat), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n483), .B1(new_n484), .B2(G50gat), .ZN(new_n485));
  INV_X1    g284(.A(G50gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(G43gat), .ZN(new_n487));
  AOI22_X1  g286(.A1(new_n485), .A2(new_n487), .B1(G29gat), .B2(G36gat), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT14), .ZN(new_n489));
  INV_X1    g288(.A(G29gat), .ZN(new_n490));
  INV_X1    g289(.A(G36gat), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT78), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n495));
  NOR2_X1   g294(.A1(G29gat), .A2(G36gat), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n496), .A2(KEYINPUT78), .A3(new_n489), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n484), .A2(KEYINPUT76), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT76), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(G43gat), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n499), .A2(new_n501), .A3(KEYINPUT77), .A4(new_n486), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(new_n483), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT77), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n504), .B1(new_n486), .B2(G43gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(KEYINPUT76), .B(G43gat), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n505), .B1(new_n506), .B2(new_n486), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n488), .B(new_n498), .C1(new_n503), .C2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT79), .ZN(new_n509));
  NAND2_X1  g308(.A1(G29gat), .A2(G36gat), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n489), .A2(new_n490), .A3(new_n491), .A4(KEYINPUT75), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(new_n495), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT75), .B1(new_n496), .B2(new_n489), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n485), .A2(new_n487), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n508), .A2(new_n509), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n509), .B1(new_n508), .B2(new_n516), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n482), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n508), .A2(KEYINPUT17), .A3(new_n516), .ZN(new_n520));
  NAND2_X1  g319(.A1(G85gat), .A2(G92gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT7), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT7), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n523), .A2(G85gat), .A3(G92gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  OR2_X1    g324(.A1(G99gat), .A2(G106gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(G99gat), .A2(G106gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OR2_X1    g327(.A1(G85gat), .A2(G92gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(KEYINPUT8), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n525), .A2(new_n528), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT87), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI22_X1  g332(.A1(new_n522), .A2(new_n524), .B1(KEYINPUT8), .B2(new_n527), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n534), .A2(KEYINPUT87), .A3(new_n528), .A4(new_n529), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n529), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n537), .A2(new_n527), .A3(new_n526), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n519), .A2(new_n520), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n508), .A2(new_n516), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT79), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n508), .A2(new_n509), .A3(new_n516), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n539), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(G190gat), .B(G218gat), .Z(new_n547));
  NAND3_X1  g346(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n540), .A2(new_n546), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n481), .B1(new_n549), .B2(KEYINPUT89), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n540), .A2(new_n546), .A3(new_n548), .ZN(new_n551));
  INV_X1    g350(.A(new_n547), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OR2_X1    g352(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n549), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n555), .A2(KEYINPUT88), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n550), .A2(new_n553), .ZN(new_n557));
  AND3_X1   g356(.A1(new_n554), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n556), .B1(new_n554), .B2(new_n557), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n477), .A2(new_n560), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n427), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G229gat), .A2(G233gat), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n519), .A2(new_n455), .A3(new_n520), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n453), .B(G8gat), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT81), .B1(new_n544), .B2(new_n565), .ZN(new_n566));
  OAI211_X1 g365(.A(KEYINPUT81), .B(new_n565), .C1(new_n517), .C2(new_n518), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n563), .B(new_n564), .C1(new_n566), .C2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT18), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n565), .B1(new_n517), .B2(new_n518), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT81), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(new_n567), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n542), .A2(new_n543), .A3(new_n455), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n563), .B(KEYINPUT13), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n575), .A2(KEYINPUT18), .A3(new_n563), .A4(new_n564), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n571), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT74), .B(KEYINPUT11), .ZN(new_n583));
  XNOR2_X1  g382(.A(G169gat), .B(G197gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G113gat), .B(G141gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT12), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n582), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n571), .A2(new_n580), .A3(new_n588), .A4(new_n581), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n436), .A2(new_n446), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n539), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT10), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n528), .B(KEYINPUT90), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(new_n537), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n536), .A2(new_n598), .A3(new_n446), .A4(new_n436), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n595), .A2(new_n596), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n545), .A2(KEYINPUT10), .A3(new_n447), .ZN(new_n601));
  AOI22_X1  g400(.A1(new_n600), .A2(new_n601), .B1(G230gat), .B2(G233gat), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n595), .A2(new_n599), .ZN(new_n603));
  NAND2_X1  g402(.A1(G230gat), .A2(G233gat), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G120gat), .B(G148gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(G176gat), .B(G204gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  NOR3_X1   g407(.A1(new_n602), .A2(new_n605), .A3(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n608), .B(KEYINPUT91), .Z(new_n611));
  XNOR2_X1  g410(.A(new_n604), .B(KEYINPUT92), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n613), .B1(new_n600), .B2(new_n601), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n611), .B1(new_n605), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n593), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n562), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n618), .A2(new_n379), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT93), .B(G1gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(G1324gat));
  INV_X1    g420(.A(new_n376), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n451), .A2(new_n454), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT42), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n626), .A2(KEYINPUT94), .A3(new_n627), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(KEYINPUT94), .B1(new_n626), .B2(new_n627), .ZN(new_n631));
  OAI221_X1 g430(.A(new_n628), .B1(new_n454), .B2(new_n623), .C1(new_n630), .C2(new_n631), .ZN(G1325gat));
  INV_X1    g431(.A(new_n618), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n424), .A2(new_n425), .ZN(new_n634));
  AND3_X1   g433(.A1(new_n633), .A2(G15gat), .A3(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n270), .A2(new_n271), .ZN(new_n636));
  AOI21_X1  g435(.A(G15gat), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n635), .A2(new_n637), .ZN(G1326gat));
  NOR2_X1   g437(.A1(new_n618), .A2(new_n387), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(G22gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT95), .B(KEYINPUT43), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(G1327gat));
  NAND2_X1  g441(.A1(new_n427), .A2(new_n560), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT44), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n477), .A2(new_n617), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(G29gat), .B1(new_n647), .B2(new_n379), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n643), .A2(new_n645), .ZN(new_n649));
  INV_X1    g448(.A(new_n379), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n649), .A2(new_n490), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT45), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n648), .A2(new_n652), .ZN(G1328gat));
  NAND3_X1  g452(.A1(new_n649), .A2(new_n491), .A3(new_n376), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n654), .B1(KEYINPUT96), .B2(KEYINPUT46), .ZN(new_n655));
  NAND2_X1  g454(.A1(KEYINPUT96), .A2(KEYINPUT46), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n655), .B(new_n656), .Z(new_n657));
  OAI21_X1  g456(.A(G36gat), .B1(new_n647), .B2(new_n622), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(G1329gat));
  INV_X1    g458(.A(new_n634), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n506), .B1(new_n647), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n636), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n662), .A2(new_n506), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n649), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT47), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(G1330gat));
  INV_X1    g466(.A(KEYINPUT48), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n644), .A2(new_n321), .A3(new_n646), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(G50gat), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n649), .A2(new_n486), .A3(new_n321), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n668), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AND3_X1   g471(.A1(new_n669), .A2(KEYINPUT97), .A3(G50gat), .ZN(new_n673));
  AOI22_X1  g472(.A1(new_n669), .A2(G50gat), .B1(KEYINPUT97), .B2(new_n668), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n671), .B(KEYINPUT98), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n672), .B1(new_n675), .B2(new_n676), .ZN(G1331gat));
  AND3_X1   g476(.A1(new_n427), .A2(new_n593), .A3(new_n561), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n616), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n679), .A2(new_n379), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(new_n440), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1332gat));
  AND2_X1   g482(.A1(new_n678), .A2(new_n616), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n622), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n685), .B(KEYINPUT101), .Z(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT102), .ZN(new_n688));
  OR2_X1    g487(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1333gat));
  OAI21_X1  g489(.A(G71gat), .B1(new_n679), .B2(new_n660), .ZN(new_n691));
  XOR2_X1   g490(.A(new_n636), .B(KEYINPUT103), .Z(new_n692));
  OR2_X1    g491(.A1(new_n692), .A2(G71gat), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n691), .B1(new_n679), .B2(new_n693), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n694), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g494(.A1(new_n684), .A2(new_n321), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(G78gat), .ZN(G1335gat));
  INV_X1    g496(.A(KEYINPUT106), .ZN(new_n698));
  INV_X1    g497(.A(new_n616), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n700));
  INV_X1    g499(.A(new_n560), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n701), .B1(new_n396), .B2(new_n426), .ZN(new_n702));
  INV_X1    g501(.A(new_n477), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n703), .A2(new_n592), .ZN(new_n704));
  AOI211_X1 g503(.A(new_n700), .B(KEYINPUT51), .C1(new_n702), .C2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n427), .A2(new_n560), .A3(new_n704), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT51), .ZN(new_n707));
  AOI21_X1  g506(.A(KEYINPUT105), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n427), .A2(KEYINPUT51), .A3(new_n560), .A4(new_n704), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT104), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT104), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n702), .A2(new_n712), .A3(KEYINPUT51), .A4(new_n704), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n699), .B1(new_n709), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(G85gat), .B1(new_n715), .B2(new_n650), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n644), .A2(new_n616), .A3(new_n704), .ZN(new_n717));
  INV_X1    g516(.A(G85gat), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n717), .A2(new_n718), .A3(new_n379), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n698), .B1(new_n716), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n706), .A2(new_n707), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n700), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n706), .A2(KEYINPUT105), .A3(new_n707), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n711), .A2(new_n713), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n616), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n718), .B1(new_n726), .B2(new_n379), .ZN(new_n727));
  OR3_X1    g526(.A1(new_n717), .A2(new_n718), .A3(new_n379), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n727), .A2(KEYINPUT106), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n720), .A2(new_n729), .ZN(G1336gat));
  NAND4_X1  g529(.A1(new_n644), .A2(new_n616), .A3(new_n376), .A4(new_n704), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT52), .B1(new_n731), .B2(G92gat), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n622), .A2(G92gat), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n732), .B1(new_n726), .B2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT52), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT51), .B1(new_n706), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n737), .B2(new_n706), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n699), .B1(new_n739), .B2(new_n714), .ZN(new_n740));
  AOI22_X1  g539(.A1(new_n740), .A2(new_n733), .B1(new_n731), .B2(G92gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n735), .B1(new_n736), .B2(new_n741), .ZN(G1337gat));
  XOR2_X1   g541(.A(KEYINPUT108), .B(G99gat), .Z(new_n743));
  OAI21_X1  g542(.A(new_n743), .B1(new_n717), .B2(new_n660), .ZN(new_n744));
  OR2_X1    g543(.A1(new_n726), .A2(new_n743), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n745), .B2(new_n662), .ZN(G1338gat));
  NAND4_X1  g545(.A1(new_n644), .A2(new_n616), .A3(new_n321), .A4(new_n704), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT53), .B1(new_n747), .B2(G106gat), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n387), .A2(G106gat), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n748), .B1(new_n726), .B2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT53), .ZN(new_n752));
  AOI22_X1  g551(.A1(new_n740), .A2(new_n749), .B1(new_n747), .B2(G106gat), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(G1339gat));
  NOR4_X1   g553(.A1(new_n477), .A2(new_n560), .A3(new_n592), .A4(new_n616), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT55), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT109), .ZN(new_n757));
  AOI211_X1 g556(.A(KEYINPUT54), .B(new_n613), .C1(new_n600), .C2(new_n601), .ZN(new_n758));
  INV_X1    g557(.A(new_n608), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT54), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n614), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n762), .A2(KEYINPUT109), .A3(new_n608), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n600), .A2(new_n601), .A3(new_n613), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n765), .A2(new_n602), .A3(new_n761), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n756), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n766), .B1(new_n760), .B2(new_n763), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n609), .B1(new_n768), .B2(KEYINPUT55), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n592), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n576), .B(new_n578), .C1(new_n566), .C2(new_n568), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT110), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n564), .B1(new_n566), .B2(new_n568), .ZN(new_n773));
  INV_X1    g572(.A(new_n563), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT110), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n575), .A2(new_n776), .A3(new_n576), .A4(new_n578), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n772), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n587), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n779), .A2(new_n591), .A3(new_n616), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n779), .A2(KEYINPUT111), .A3(new_n591), .A4(new_n616), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n770), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n701), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n779), .A2(new_n591), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n560), .A2(new_n769), .A3(new_n767), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n755), .B1(new_n477), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n789), .A2(new_n389), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n790), .A2(new_n650), .A3(new_n622), .ZN(new_n791));
  INV_X1    g590(.A(G113gat), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n791), .A2(new_n792), .A3(new_n593), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n790), .A2(new_n650), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT112), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n790), .A2(new_n796), .A3(new_n650), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n798), .A2(new_n592), .A3(new_n622), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n793), .B1(new_n799), .B2(new_n792), .ZN(G1340gat));
  OAI21_X1  g599(.A(G120gat), .B1(new_n791), .B2(new_n699), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n622), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n699), .A2(G120gat), .ZN(new_n803));
  XOR2_X1   g602(.A(new_n803), .B(KEYINPUT113), .Z(new_n804));
  OAI21_X1  g603(.A(new_n801), .B1(new_n802), .B2(new_n804), .ZN(G1341gat));
  NOR2_X1   g604(.A1(new_n477), .A2(G127gat), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n795), .A2(new_n622), .A3(new_n797), .A4(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(G127gat), .B1(new_n791), .B2(new_n477), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT114), .ZN(G1342gat));
  OAI21_X1  g609(.A(G134gat), .B1(new_n791), .B2(new_n701), .ZN(new_n811));
  INV_X1    g610(.A(G134gat), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n560), .A2(new_n622), .ZN(new_n813));
  XOR2_X1   g612(.A(new_n813), .B(KEYINPUT115), .Z(new_n814));
  NAND4_X1  g613(.A1(new_n795), .A2(new_n812), .A3(new_n797), .A4(new_n814), .ZN(new_n815));
  XOR2_X1   g614(.A(KEYINPUT116), .B(KEYINPUT56), .Z(new_n816));
  AND2_X1   g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n815), .A2(new_n816), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n811), .B1(new_n817), .B2(new_n818), .ZN(G1343gat));
  NOR2_X1   g618(.A1(new_n634), .A2(new_n387), .ZN(new_n820));
  XOR2_X1   g619(.A(new_n820), .B(KEYINPUT118), .Z(new_n821));
  NAND2_X1  g620(.A1(new_n788), .A2(new_n477), .ZN(new_n822));
  INV_X1    g621(.A(new_n755), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n821), .A2(new_n650), .A3(new_n824), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n825), .A2(new_n622), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n593), .A2(G141gat), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n770), .A2(new_n780), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n701), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n829), .A2(new_n701), .A3(KEYINPUT117), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n832), .A2(new_n787), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n755), .B1(new_n834), .B2(new_n477), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT57), .B1(new_n835), .B2(new_n387), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n387), .B1(new_n822), .B2(new_n823), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT57), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n622), .A2(new_n650), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n634), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n836), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(G141gat), .B1(new_n842), .B2(new_n593), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n845), .B1(new_n843), .B2(KEYINPUT119), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n828), .B(new_n843), .C1(KEYINPUT119), .C2(new_n845), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(G1344gat));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n850), .B(G148gat), .C1(new_n842), .C2(new_n699), .ZN(new_n851));
  INV_X1    g650(.A(G148gat), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n634), .A2(new_n699), .A3(new_n840), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n703), .B1(new_n830), .B2(new_n787), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n838), .B(new_n321), .C1(new_n854), .C2(new_n755), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n853), .B(new_n855), .C1(new_n837), .C2(new_n838), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n852), .B1(new_n856), .B2(KEYINPUT120), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT57), .B1(new_n789), .B2(new_n387), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT120), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n858), .A2(new_n859), .A3(new_n853), .A4(new_n855), .ZN(new_n860));
  AOI211_X1 g659(.A(KEYINPUT121), .B(new_n850), .C1(new_n857), .C2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT121), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n856), .A2(KEYINPUT120), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n863), .A2(G148gat), .A3(new_n860), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n862), .B1(new_n864), .B2(KEYINPUT59), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n851), .B1(new_n861), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n826), .A2(new_n852), .A3(new_n616), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(G1345gat));
  NOR3_X1   g667(.A1(new_n842), .A2(new_n289), .A3(new_n477), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n826), .A2(new_n703), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n869), .B1(new_n870), .B2(new_n289), .ZN(G1346gat));
  OAI21_X1  g670(.A(G162gat), .B1(new_n842), .B2(new_n701), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n825), .A2(new_n290), .A3(new_n814), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(G1347gat));
  NOR2_X1   g673(.A1(new_n622), .A2(new_n650), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n790), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(new_n226), .A3(new_n592), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n789), .A2(new_n650), .A3(new_n622), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n692), .A2(new_n321), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n592), .A3(new_n880), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n881), .A2(KEYINPUT122), .A3(G169gat), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT122), .B1(new_n881), .B2(G169gat), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n878), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT123), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n884), .B(new_n885), .ZN(G1348gat));
  AOI21_X1  g685(.A(G176gat), .B1(new_n877), .B2(new_n616), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n879), .A2(new_n880), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n888), .A2(new_n227), .A3(new_n699), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n887), .A2(new_n889), .ZN(G1349gat));
  OAI21_X1  g689(.A(new_n209), .B1(new_n888), .B2(new_n477), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n876), .A2(new_n224), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n891), .B1(new_n892), .B2(new_n477), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g693(.A1(new_n877), .A2(new_n214), .A3(new_n560), .ZN(new_n895));
  OAI21_X1  g694(.A(G190gat), .B1(new_n888), .B2(new_n701), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n896), .A2(KEYINPUT61), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n896), .A2(KEYINPUT61), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n895), .B1(new_n897), .B2(new_n898), .ZN(G1351gat));
  NAND2_X1  g698(.A1(new_n858), .A2(new_n855), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT124), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n900), .B(new_n901), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n634), .A2(new_n650), .A3(new_n622), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n902), .A2(KEYINPUT125), .A3(new_n592), .A4(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(new_n855), .ZN(new_n905));
  INV_X1    g704(.A(new_n837), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n905), .B1(new_n906), .B2(KEYINPUT57), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n901), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n900), .A2(KEYINPUT124), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n908), .A2(new_n909), .A3(new_n592), .A4(new_n903), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT125), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n904), .A2(new_n912), .A3(G197gat), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n879), .A2(new_n820), .ZN(new_n914));
  OR3_X1    g713(.A1(new_n914), .A2(G197gat), .A3(new_n593), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(G1352gat));
  NAND2_X1  g715(.A1(new_n902), .A2(new_n903), .ZN(new_n917));
  OAI21_X1  g716(.A(G204gat), .B1(new_n917), .B2(new_n699), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(KEYINPUT126), .ZN(new_n920));
  INV_X1    g719(.A(G204gat), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n879), .A2(new_n820), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n920), .B1(new_n922), .B2(new_n699), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n919), .A2(KEYINPUT126), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n923), .B(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n918), .A2(new_n925), .ZN(G1353gat));
  OR3_X1    g725(.A1(new_n914), .A2(G211gat), .A3(new_n477), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n907), .A2(KEYINPUT127), .A3(new_n703), .A4(new_n903), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n858), .A2(new_n703), .A3(new_n855), .A4(new_n903), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT127), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n928), .A2(new_n931), .A3(G211gat), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT63), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n932), .A2(new_n933), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n927), .B1(new_n934), .B2(new_n935), .ZN(G1354gat));
  OAI21_X1  g735(.A(G218gat), .B1(new_n917), .B2(new_n701), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n914), .A2(G218gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n701), .B2(new_n938), .ZN(G1355gat));
endmodule


