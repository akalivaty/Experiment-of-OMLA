//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 0 1 0 1 0 1 0 1 0 0 1 1 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 0 1 1 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT11), .B1(new_n192), .B2(G134), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(G134), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(new_n192), .ZN(new_n197));
  NAND2_X1  g011(.A1(KEYINPUT65), .A2(G137), .ZN(new_n198));
  AND2_X1   g012(.A1(KEYINPUT11), .A2(G134), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n197), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  AND3_X1   g015(.A1(new_n195), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n201), .B1(new_n195), .B2(new_n200), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G107), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G104), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT76), .ZN(new_n207));
  INV_X1    g021(.A(G104), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n207), .B1(new_n208), .B2(G107), .ZN(new_n209));
  NOR3_X1   g023(.A1(new_n205), .A2(KEYINPUT76), .A3(G104), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n206), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G101), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G143), .ZN(new_n214));
  INV_X1    g028(.A(G143), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G146), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n214), .B(new_n216), .C1(KEYINPUT1), .C2(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT1), .B1(new_n215), .B2(G146), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n215), .A2(G146), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n213), .A2(G143), .ZN(new_n221));
  OAI211_X1 g035(.A(G128), .B(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G101), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n208), .A2(G107), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n205), .A2(KEYINPUT3), .A3(G104), .ZN(new_n225));
  AOI21_X1  g039(.A(KEYINPUT3), .B1(new_n205), .B2(G104), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n223), .B(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n212), .A2(new_n218), .A3(new_n222), .A4(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT10), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n230), .B1(new_n208), .B2(G107), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n205), .A2(KEYINPUT3), .A3(G104), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n223), .B1(new_n233), .B2(new_n224), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT4), .ZN(new_n235));
  NAND2_X1  g049(.A1(KEYINPUT0), .A2(G128), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(KEYINPUT0), .A2(G128), .ZN(new_n238));
  OAI22_X1  g052(.A1(new_n220), .A2(new_n221), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n214), .A2(new_n216), .A3(new_n236), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n234), .A2(new_n235), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n205), .A2(G104), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n242), .B1(new_n231), .B2(new_n232), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n235), .B1(new_n243), .B2(new_n223), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G101), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  AOI22_X1  g061(.A1(new_n228), .A2(new_n229), .B1(new_n241), .B2(new_n247), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n222), .A2(new_n218), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n249), .A2(KEYINPUT10), .A3(new_n227), .A4(new_n212), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n204), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(KEYINPUT76), .B1(new_n205), .B2(G104), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n207), .A2(new_n208), .A3(G107), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n252), .A2(new_n253), .B1(G104), .B2(new_n205), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n227), .B1(new_n254), .B2(new_n223), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n222), .A2(new_n218), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n229), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n239), .A2(new_n240), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n245), .A2(new_n235), .A3(G101), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n227), .A2(KEYINPUT4), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n258), .B(new_n259), .C1(new_n260), .C2(new_n234), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n257), .A2(new_n261), .A3(new_n250), .A4(new_n204), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(G110), .B(G140), .ZN(new_n264));
  INV_X1    g078(.A(G227), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(G953), .ZN(new_n266));
  XOR2_X1   g080(.A(new_n264), .B(new_n266), .Z(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NOR3_X1   g082(.A1(new_n251), .A2(new_n263), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT77), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n255), .A2(new_n256), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n204), .B1(new_n271), .B2(new_n228), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n270), .B1(new_n272), .B2(KEYINPUT12), .ZN(new_n273));
  INV_X1    g087(.A(new_n204), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n255), .A2(new_n256), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n212), .A2(new_n227), .B1(new_n218), .B2(new_n222), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT12), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n277), .A2(KEYINPUT77), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n272), .A2(KEYINPUT12), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n273), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n262), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n269), .B1(new_n282), .B2(new_n268), .ZN(new_n283));
  OAI21_X1  g097(.A(G469), .B1(new_n283), .B2(G902), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n268), .B1(new_n251), .B2(new_n263), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT79), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n263), .A2(new_n268), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n281), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n257), .A2(new_n261), .A3(new_n250), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n274), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n267), .B1(new_n291), .B2(new_n262), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT79), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n287), .A2(new_n289), .A3(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT68), .B(G902), .ZN(new_n295));
  XNOR2_X1  g109(.A(KEYINPUT78), .B(G469), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n191), .B1(new_n284), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT80), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n298), .B(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G224), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT7), .B1(new_n301), .B2(G953), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n239), .A2(new_n240), .A3(G125), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(G125), .B1(new_n222), .B2(new_n218), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n303), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT82), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n304), .B(new_n302), .C1(new_n306), .C2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G125), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n256), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n311), .A2(KEYINPUT82), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n307), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G113), .ZN(new_n314));
  INV_X1    g128(.A(G116), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n315), .A2(G119), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT5), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n314), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G119), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G116), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n315), .A2(G119), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(KEYINPUT5), .ZN(new_n322));
  XNOR2_X1  g136(.A(G116), .B(G119), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n314), .A2(KEYINPUT2), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT2), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G113), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n318), .A2(new_n322), .B1(new_n323), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n212), .A2(new_n328), .A3(new_n227), .ZN(new_n329));
  XNOR2_X1  g143(.A(G110), .B(G122), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n260), .A2(new_n234), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n320), .A2(new_n321), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(new_n324), .A3(new_n326), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n327), .A2(new_n323), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n259), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n329), .B(new_n330), .C1(new_n331), .C2(new_n336), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n313), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n318), .A2(new_n322), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n334), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT81), .B1(new_n255), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n255), .A2(new_n340), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n255), .A2(new_n340), .A3(KEYINPUT81), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  XOR2_X1   g159(.A(new_n330), .B(KEYINPUT8), .Z(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(G902), .B1(new_n338), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(G210), .B1(G237), .B2(G902), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n329), .B1(new_n331), .B2(new_n336), .ZN(new_n351));
  INV_X1    g165(.A(new_n330), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(KEYINPUT6), .A3(new_n337), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT6), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n351), .A2(new_n355), .A3(new_n352), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n311), .A2(new_n304), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n301), .A2(G953), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n357), .B(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n354), .A2(new_n356), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n349), .A2(new_n350), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n350), .B1(new_n349), .B2(new_n360), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n361), .B1(new_n362), .B2(KEYINPUT83), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT83), .ZN(new_n364));
  AOI211_X1 g178(.A(new_n364), .B(new_n350), .C1(new_n349), .C2(new_n360), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(G214), .B1(G237), .B2(G902), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G478), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n370), .A2(KEYINPUT15), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT13), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n372), .B1(new_n217), .B2(G143), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n217), .A2(G143), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n215), .A2(G128), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n376), .A2(new_n372), .ZN(new_n377));
  OAI21_X1  g191(.A(G134), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G122), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G116), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n315), .A2(G122), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G107), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n380), .A2(new_n381), .A3(new_n205), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n217), .A2(G143), .ZN(new_n386));
  INV_X1    g200(.A(G134), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n376), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n378), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G217), .ZN(new_n390));
  NOR3_X1   g204(.A1(new_n188), .A2(new_n390), .A3(G953), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT87), .ZN(new_n392));
  AOI21_X1  g206(.A(KEYINPUT14), .B1(new_n379), .B2(G116), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n379), .A2(G116), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n381), .A2(KEYINPUT14), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n392), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n205), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n376), .A2(new_n386), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G134), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n388), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n384), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n389), .B(new_n391), .C1(new_n400), .C2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT88), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT14), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n408), .B1(new_n315), .B2(G122), .ZN(new_n409));
  AOI21_X1  g223(.A(KEYINPUT87), .B1(new_n409), .B2(new_n381), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n399), .B1(new_n410), .B2(new_n396), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G107), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(new_n384), .A3(new_n403), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n413), .A2(KEYINPUT88), .A3(new_n389), .A4(new_n391), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n389), .B1(new_n400), .B2(new_n404), .ZN(new_n415));
  INV_X1    g229(.A(new_n391), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n407), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n371), .B1(new_n418), .B2(new_n295), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n295), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT89), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n418), .A2(KEYINPUT89), .A3(new_n295), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n419), .B1(new_n424), .B2(new_n371), .ZN(new_n425));
  INV_X1    g239(.A(G140), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G125), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n310), .A2(G140), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n428), .A3(KEYINPUT16), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT70), .ZN(new_n430));
  XNOR2_X1  g244(.A(G125), .B(G140), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT70), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(new_n432), .A3(KEYINPUT16), .ZN(new_n433));
  OR2_X1    g247(.A1(new_n427), .A2(KEYINPUT16), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n430), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n213), .ZN(new_n436));
  NOR2_X1   g250(.A1(G237), .A2(G953), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(G143), .A3(G214), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(G143), .B1(new_n437), .B2(G214), .ZN(new_n440));
  OAI21_X1  g254(.A(G131), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT17), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n437), .A2(G214), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n215), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(new_n201), .A3(new_n438), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n441), .A2(new_n442), .A3(new_n445), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n430), .A2(new_n433), .A3(G146), .A4(new_n434), .ZN(new_n447));
  OAI211_X1 g261(.A(KEYINPUT17), .B(G131), .C1(new_n439), .C2(new_n440), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n436), .A2(new_n446), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(G113), .B(G122), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n450), .B(new_n208), .ZN(new_n451));
  NAND2_X1  g265(.A1(KEYINPUT18), .A2(G131), .ZN(new_n452));
  XOR2_X1   g266(.A(new_n452), .B(KEYINPUT84), .Z(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(new_n444), .A3(new_n438), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n431), .B(new_n213), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT18), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n454), .B(new_n455), .C1(new_n456), .C2(new_n441), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n449), .A2(new_n451), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n441), .A2(new_n445), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT19), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT85), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n431), .A2(new_n461), .ZN(new_n462));
  OR2_X1    g276(.A1(new_n460), .A2(KEYINPUT85), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n463), .A2(new_n461), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n462), .B1(new_n431), .B2(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n459), .B(new_n447), .C1(new_n465), .C2(G146), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n466), .A2(new_n457), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n458), .B1(new_n467), .B2(new_n451), .ZN(new_n468));
  NOR2_X1   g282(.A1(G475), .A2(G902), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(KEYINPUT20), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT20), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n468), .A2(new_n472), .A3(new_n469), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n449), .A2(new_n451), .A3(new_n457), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n451), .B1(new_n449), .B2(new_n457), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n190), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT86), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT86), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n479), .B(new_n190), .C1(new_n475), .C2(new_n476), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n478), .A2(G475), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n474), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(G952), .ZN(new_n483));
  AOI211_X1 g297(.A(G953), .B(new_n483), .C1(G234), .C2(G237), .ZN(new_n484));
  INV_X1    g298(.A(G953), .ZN(new_n485));
  AOI211_X1 g299(.A(new_n485), .B(new_n295), .C1(G234), .C2(G237), .ZN(new_n486));
  XNOR2_X1  g300(.A(KEYINPUT21), .B(G898), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n425), .A2(new_n482), .A3(new_n488), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n369), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G472), .ZN(new_n491));
  INV_X1    g305(.A(new_n295), .ZN(new_n492));
  INV_X1    g306(.A(new_n335), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n258), .B1(new_n202), .B2(new_n203), .ZN(new_n494));
  AOI21_X1  g308(.A(G134), .B1(new_n197), .B2(new_n198), .ZN(new_n495));
  INV_X1    g309(.A(new_n194), .ZN(new_n496));
  OAI21_X1  g310(.A(G131), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n195), .A2(new_n200), .A3(new_n201), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n497), .A2(new_n498), .A3(new_n218), .A4(new_n222), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n500), .A2(KEYINPUT67), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT67), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n502), .B1(new_n494), .B2(new_n499), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n493), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT28), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n500), .A2(new_n335), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n494), .A2(new_n493), .A3(new_n499), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT28), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n437), .A2(G210), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(KEYINPUT27), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT26), .B(G101), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT29), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n492), .B1(new_n511), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n509), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n506), .A2(new_n515), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT64), .ZN(new_n523));
  AOI21_X1  g337(.A(KEYINPUT30), .B1(new_n500), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT30), .ZN(new_n525));
  AOI211_X1 g339(.A(KEYINPUT64), .B(new_n525), .C1(new_n494), .C2(new_n499), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n335), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n527), .A2(new_n508), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n522), .B(new_n517), .C1(new_n528), .C2(new_n515), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n491), .B1(new_n519), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n527), .A2(new_n515), .A3(new_n508), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT31), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n527), .A2(KEYINPUT31), .A3(new_n515), .A4(new_n508), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n506), .A2(new_n521), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n516), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT32), .ZN(new_n539));
  NOR2_X1   g353(.A1(G472), .A2(G902), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n533), .A2(new_n534), .B1(new_n516), .B2(new_n536), .ZN(new_n542));
  INV_X1    g356(.A(new_n540), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT32), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n530), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n436), .A2(new_n447), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n217), .A2(G119), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n319), .A2(G128), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n547), .A2(new_n548), .A3(KEYINPUT69), .A4(KEYINPUT23), .ZN(new_n549));
  OR2_X1    g363(.A1(KEYINPUT69), .A2(KEYINPUT23), .ZN(new_n550));
  NAND2_X1  g364(.A1(KEYINPUT69), .A2(KEYINPUT23), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n550), .A2(G119), .A3(new_n217), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(G110), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n547), .A2(new_n548), .ZN(new_n555));
  XNOR2_X1  g369(.A(KEYINPUT24), .B(G110), .ZN(new_n556));
  OAI22_X1  g370(.A1(new_n553), .A2(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n546), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n431), .A2(new_n213), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n447), .A2(new_n560), .ZN(new_n561));
  XOR2_X1   g375(.A(KEYINPUT71), .B(G110), .Z(new_n562));
  AOI21_X1  g376(.A(new_n562), .B1(new_n549), .B2(new_n552), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n563), .A2(KEYINPUT72), .B1(new_n555), .B2(new_n556), .ZN(new_n564));
  INV_X1    g378(.A(new_n562), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n553), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT72), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT73), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n561), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n564), .A2(new_n568), .A3(KEYINPUT73), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT74), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n553), .A2(KEYINPUT72), .A3(new_n565), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n555), .A2(new_n556), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n563), .A2(KEYINPUT72), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n570), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n561), .ZN(new_n579));
  AND4_X1   g393(.A1(KEYINPUT74), .A2(new_n578), .A3(new_n572), .A4(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n559), .B1(new_n573), .B2(new_n580), .ZN(new_n581));
  XOR2_X1   g395(.A(KEYINPUT22), .B(G137), .Z(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(KEYINPUT75), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n485), .A2(G221), .A3(G234), .ZN(new_n584));
  XOR2_X1   g398(.A(new_n583), .B(new_n584), .Z(new_n585));
  NAND2_X1  g399(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n585), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n559), .B(new_n587), .C1(new_n573), .C2(new_n580), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n390), .B1(new_n295), .B2(G234), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(G902), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n586), .A2(new_n295), .A3(new_n588), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n593), .A2(KEYINPUT25), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT25), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n586), .A2(new_n595), .A3(new_n295), .A4(new_n588), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n590), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n592), .B1(new_n594), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n545), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n300), .A2(new_n490), .A3(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(G101), .ZN(G3));
  NAND2_X1  g415(.A1(new_n538), .A2(new_n295), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G472), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n538), .A2(new_n540), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n605), .A2(new_n598), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n300), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n350), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n354), .A2(new_n356), .A3(new_n359), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n313), .A2(new_n337), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n346), .B1(new_n343), .B2(new_n344), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n190), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n608), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n368), .B1(new_n613), .B2(new_n361), .ZN(new_n614));
  INV_X1    g428(.A(new_n488), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n422), .A2(new_n370), .A3(new_n423), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT33), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n418), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n417), .A2(KEYINPUT33), .A3(new_n405), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n618), .A2(G478), .A3(new_n295), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n614), .A2(new_n482), .A3(new_n615), .A4(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n607), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT34), .B(G104), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G6));
  OR2_X1    g439(.A1(new_n481), .A2(KEYINPUT90), .ZN(new_n626));
  AOI22_X1  g440(.A1(new_n481), .A2(KEYINPUT90), .B1(new_n471), .B2(new_n473), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n627), .A3(new_n425), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n614), .A2(new_n615), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n300), .A2(new_n606), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT91), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G107), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  INV_X1    g448(.A(new_n605), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n585), .A2(KEYINPUT36), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n581), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n581), .A2(new_n637), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n591), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n641), .B1(new_n594), .B2(new_n597), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n300), .A2(new_n490), .A3(new_n635), .A4(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT37), .B(G110), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G12));
  INV_X1    g459(.A(G900), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n486), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n484), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n626), .A2(new_n627), .A3(new_n425), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT92), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n596), .A2(new_n590), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n593), .A2(KEYINPUT25), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n652), .A2(new_n653), .B1(new_n640), .B2(new_n591), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n545), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n651), .A2(new_n300), .A3(new_n655), .A4(new_n614), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G128), .ZN(G30));
  XNOR2_X1  g471(.A(KEYINPUT93), .B(KEYINPUT38), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n366), .B(new_n658), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n425), .A2(new_n482), .A3(new_n367), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n659), .A2(new_n654), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n516), .B1(new_n527), .B2(new_n508), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT94), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n509), .A2(new_n515), .ZN(new_n664));
  OR3_X1    g478(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n663), .B1(new_n662), .B2(new_n664), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n665), .A2(new_n190), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(G472), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT95), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n541), .A2(new_n544), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n667), .A2(KEYINPUT95), .A3(G472), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n673), .A2(KEYINPUT96), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n673), .A2(KEYINPUT96), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n661), .B(KEYINPUT97), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n649), .B(KEYINPUT39), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n300), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT40), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n300), .A2(KEYINPUT40), .A3(new_n677), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n676), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n673), .B(KEYINPUT96), .ZN(new_n684));
  AOI21_X1  g498(.A(KEYINPUT97), .B1(new_n684), .B2(new_n661), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(new_n215), .ZN(G45));
  NAND3_X1  g501(.A1(new_n621), .A2(new_n482), .A3(new_n649), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n300), .A2(new_n655), .A3(new_n614), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G146), .ZN(G48));
  INV_X1    g505(.A(new_n191), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n292), .B(new_n286), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n492), .B1(new_n693), .B2(new_n289), .ZN(new_n694));
  INV_X1    g508(.A(G469), .ZN(new_n695));
  OAI211_X1 g509(.A(new_n692), .B(new_n297), .C1(new_n694), .C2(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n696), .A2(new_n622), .ZN(new_n697));
  INV_X1    g511(.A(new_n530), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n539), .B1(new_n538), .B2(new_n540), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n542), .A2(KEYINPUT32), .A3(new_n543), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  AOI22_X1  g515(.A1(new_n652), .A2(new_n653), .B1(new_n591), .B2(new_n589), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n697), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT98), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n599), .A2(KEYINPUT98), .A3(new_n697), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT41), .B(G113), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  INV_X1    g523(.A(new_n696), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n701), .A2(new_n702), .A3(new_n630), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G116), .ZN(G18));
  NAND2_X1  g526(.A1(new_n294), .A2(new_n295), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(G469), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n714), .A2(new_n692), .A3(new_n297), .A4(new_n614), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT99), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n489), .A3(new_n655), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G119), .ZN(G21));
  NOR2_X1   g532(.A1(new_n696), .A2(new_n488), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n540), .B(KEYINPUT100), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n506), .A2(new_n510), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n516), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n720), .B1(new_n535), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n723), .B1(new_n602), .B2(G472), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n613), .A2(new_n361), .ZN(new_n725));
  AND4_X1   g539(.A1(new_n425), .A2(new_n725), .A3(new_n482), .A4(new_n367), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n719), .A2(new_n702), .A3(new_n724), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT101), .B(G122), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G24));
  AND3_X1   g543(.A1(new_n642), .A2(new_n724), .A3(KEYINPUT102), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT102), .B1(new_n642), .B2(new_n724), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n716), .B(new_n689), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G125), .ZN(G27));
  NAND2_X1  g547(.A1(new_n284), .A2(new_n297), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT103), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR4_X1   g550(.A1(new_n363), .A2(new_n365), .A3(new_n191), .A4(new_n368), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n284), .A2(KEYINPUT103), .A3(new_n297), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NOR4_X1   g553(.A1(new_n739), .A2(new_n545), .A3(new_n598), .A4(new_n688), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT104), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT105), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n741), .B1(new_n742), .B2(KEYINPUT42), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n743), .B1(new_n742), .B2(KEYINPUT42), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n739), .ZN(new_n746));
  AOI21_X1  g560(.A(KEYINPUT42), .B1(new_n742), .B2(KEYINPUT104), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n746), .A2(new_n599), .A3(new_n689), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n201), .ZN(G33));
  NAND3_X1  g564(.A1(new_n651), .A2(new_n746), .A3(new_n599), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G134), .ZN(G36));
  AND2_X1   g566(.A1(new_n474), .A2(new_n481), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n621), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n754), .A2(KEYINPUT43), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT43), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n756), .B1(new_n753), .B2(new_n621), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n758), .A2(KEYINPUT44), .A3(new_n605), .A4(new_n642), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n363), .A2(new_n368), .A3(new_n365), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n297), .ZN(new_n762));
  OAI21_X1  g576(.A(G469), .B1(new_n283), .B2(KEYINPUT45), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n283), .A2(KEYINPUT45), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT106), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n283), .A2(KEYINPUT106), .A3(KEYINPUT45), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n763), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n695), .A2(new_n190), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n762), .B1(new_n770), .B2(KEYINPUT46), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT46), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n772), .B1(new_n768), .B2(new_n769), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n191), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT44), .ZN(new_n775));
  INV_X1    g589(.A(new_n758), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n605), .A2(new_n642), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n761), .A2(new_n774), .A3(new_n677), .A4(new_n778), .ZN(new_n779));
  XOR2_X1   g593(.A(KEYINPUT107), .B(G137), .Z(new_n780));
  XNOR2_X1  g594(.A(new_n779), .B(new_n780), .ZN(G39));
  INV_X1    g595(.A(new_n760), .ZN(new_n782));
  NOR4_X1   g596(.A1(new_n701), .A2(new_n702), .A3(new_n782), .A4(new_n688), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n774), .A2(KEYINPUT47), .ZN(new_n784));
  INV_X1    g598(.A(new_n769), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n766), .A2(new_n767), .ZN(new_n786));
  OAI211_X1 g600(.A(KEYINPUT46), .B(new_n785), .C1(new_n786), .C2(new_n763), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n787), .A2(new_n297), .A3(new_n773), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n692), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT47), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n783), .B1(new_n784), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  AOI21_X1  g607(.A(new_n695), .B1(new_n294), .B2(new_n295), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n762), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n737), .A2(new_n484), .A3(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n776), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n797), .B1(new_n731), .B2(new_n730), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n674), .A2(new_n675), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n796), .A2(new_n598), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n753), .A2(new_n616), .A3(new_n620), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n798), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AND4_X1   g617(.A1(new_n702), .A2(new_n758), .A3(new_n484), .A4(new_n724), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n659), .A2(new_n367), .A3(new_n696), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n804), .A2(new_n805), .A3(KEYINPUT50), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT115), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n804), .A2(new_n805), .A3(new_n808), .A4(KEYINPUT50), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n804), .A2(new_n805), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n811), .A2(KEYINPUT50), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n803), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n789), .B(new_n790), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n762), .A2(new_n794), .A3(new_n692), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n760), .B(new_n804), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n813), .A2(new_n816), .A3(KEYINPUT51), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n621), .A2(new_n482), .ZN(new_n818));
  OR2_X1    g632(.A1(new_n801), .A2(new_n818), .ZN(new_n819));
  AOI211_X1 g633(.A(new_n483), .B(G953), .C1(new_n804), .C2(new_n716), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT116), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n797), .A2(new_n599), .ZN(new_n822));
  XOR2_X1   g636(.A(new_n822), .B(KEYINPUT48), .Z(new_n823));
  NOR2_X1   g637(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n819), .A2(new_n820), .A3(KEYINPUT116), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n817), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT51), .B1(new_n813), .B2(new_n816), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n726), .A2(new_n692), .A3(new_n649), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n736), .A2(new_n738), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n673), .A2(new_n829), .A3(new_n830), .A4(new_n654), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n831), .A2(KEYINPUT52), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT112), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n732), .A2(new_n833), .A3(new_n656), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n833), .B1(new_n732), .B2(new_n656), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n690), .B(new_n832), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n732), .A2(new_n656), .A3(new_n690), .A4(new_n831), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT98), .B1(new_n599), .B2(new_n697), .ZN(new_n841));
  AND4_X1   g655(.A1(KEYINPUT98), .A2(new_n697), .A3(new_n701), .A4(new_n702), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT99), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n715), .B(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n701), .A2(new_n489), .A3(new_n642), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n711), .B(new_n727), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(KEYINPUT110), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n711), .A2(new_n727), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT110), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n707), .A2(new_n849), .A3(new_n850), .A4(new_n717), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n425), .A2(KEYINPUT111), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n425), .A2(KEYINPUT111), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n818), .B1(new_n854), .B2(new_n482), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n369), .A2(new_n615), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n300), .A2(new_n855), .A3(new_n857), .A4(new_n606), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n858), .A2(new_n643), .A3(new_n600), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n848), .A2(new_n851), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n688), .A2(new_n191), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(new_n736), .A3(new_n738), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n642), .A2(new_n724), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT102), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n642), .A2(new_n724), .A3(KEYINPUT102), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n862), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n626), .A2(new_n627), .A3(new_n649), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n298), .A2(new_n299), .ZN(new_n869));
  AOI211_X1 g683(.A(KEYINPUT80), .B(new_n191), .C1(new_n284), .C2(new_n297), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n854), .B(new_n868), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n701), .A2(new_n642), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n760), .B1(new_n867), .B2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(new_n745), .A3(new_n748), .A4(new_n751), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n860), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT53), .B1(new_n840), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n837), .B(KEYINPUT52), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n830), .B(new_n861), .C1(new_n730), .C2(new_n731), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n300), .A2(new_n655), .A3(new_n854), .A4(new_n868), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n782), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n748), .B(new_n751), .C1(new_n740), .C2(new_n744), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n883), .A2(new_n848), .A3(new_n851), .A4(new_n859), .ZN(new_n884));
  XOR2_X1   g698(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n885));
  NOR3_X1   g699(.A1(new_n878), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(KEYINPUT54), .B1(new_n877), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n885), .B1(new_n878), .B2(new_n884), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n843), .A2(new_n847), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n883), .A2(new_n890), .A3(new_n859), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n840), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g707(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n888), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n887), .A2(new_n895), .ZN(new_n896));
  OAI22_X1  g710(.A1(new_n828), .A2(new_n896), .B1(G952), .B2(G953), .ZN(new_n897));
  NOR4_X1   g711(.A1(new_n598), .A2(new_n191), .A3(new_n368), .A4(new_n754), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n899), .A2(KEYINPUT108), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(KEYINPUT108), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n795), .B(KEYINPUT49), .Z(new_n902));
  NOR2_X1   g716(.A1(new_n902), .A2(new_n659), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n900), .A2(new_n799), .A3(new_n901), .A4(new_n903), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT109), .Z(new_n905));
  NAND2_X1  g719(.A1(new_n897), .A2(new_n905), .ZN(G75));
  INV_X1    g720(.A(new_n885), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n837), .B(new_n838), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n907), .B1(new_n876), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n891), .B1(new_n839), .B2(new_n836), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n492), .B(new_n608), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(KEYINPUT117), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n354), .A2(new_n356), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(new_n359), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT55), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT56), .ZN(new_n916));
  AOI22_X1  g730(.A1(new_n912), .A2(new_n915), .B1(new_n916), .B2(new_n911), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT117), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n911), .A2(new_n918), .A3(new_n916), .A4(new_n915), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n485), .A2(G952), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n917), .A2(new_n922), .ZN(G51));
  XOR2_X1   g737(.A(new_n769), .B(KEYINPUT118), .Z(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT57), .ZN(new_n925));
  INV_X1    g739(.A(new_n895), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n894), .B1(new_n888), .B2(new_n893), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n294), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n888), .A2(new_n893), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n930), .A2(new_n492), .A3(new_n768), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n920), .B1(new_n929), .B2(new_n931), .ZN(G54));
  AND2_X1   g746(.A1(KEYINPUT58), .A2(G475), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n492), .B(new_n933), .C1(new_n909), .C2(new_n910), .ZN(new_n934));
  INV_X1    g748(.A(new_n468), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n930), .A2(new_n492), .A3(new_n468), .A4(new_n933), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n936), .A2(new_n921), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(KEYINPUT119), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT119), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n936), .A2(new_n940), .A3(new_n937), .A4(new_n921), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n939), .A2(new_n941), .ZN(G60));
  NAND2_X1  g756(.A1(new_n618), .A2(new_n619), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(G478), .A2(G902), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT59), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n944), .B(new_n946), .C1(new_n926), .C2(new_n927), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n921), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n944), .B1(new_n896), .B2(new_n946), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(G63));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n951));
  NAND2_X1  g765(.A1(G217), .A2(G902), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT60), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n953), .B1(new_n888), .B2(new_n893), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n640), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n921), .B1(new_n954), .B2(new_n589), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n951), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n954), .A2(new_n589), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n959), .A2(KEYINPUT61), .A3(new_n921), .A4(new_n955), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n958), .A2(new_n960), .ZN(G66));
  XNOR2_X1  g775(.A(new_n860), .B(KEYINPUT120), .ZN(new_n962));
  OR3_X1    g776(.A1(new_n962), .A2(KEYINPUT121), .A3(G953), .ZN(new_n963));
  OAI21_X1  g777(.A(KEYINPUT121), .B1(new_n962), .B2(G953), .ZN(new_n964));
  OAI21_X1  g778(.A(G953), .B1(new_n487), .B2(new_n301), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n913), .B1(G898), .B2(new_n485), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(G69));
  OAI21_X1  g782(.A(G953), .B1(new_n265), .B2(new_n646), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n524), .A2(new_n526), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n465), .B(KEYINPUT122), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n970), .B(new_n971), .Z(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(G900), .B2(G953), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n774), .A2(new_n599), .A3(new_n677), .A4(new_n726), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT125), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n745), .A2(new_n976), .A3(new_n748), .A4(new_n751), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n882), .A2(KEYINPUT125), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n792), .A2(new_n975), .A3(new_n977), .A4(new_n978), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n690), .B(new_n779), .C1(new_n834), .C2(new_n835), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(KEYINPUT124), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n732), .A2(new_n656), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(KEYINPUT112), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n732), .A2(new_n833), .A3(new_n656), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT124), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n985), .A2(new_n986), .A3(new_n690), .A4(new_n779), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n979), .B1(new_n981), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n974), .B1(new_n988), .B2(new_n485), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT123), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n969), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n855), .A2(new_n599), .A3(new_n760), .ZN(new_n992));
  OAI211_X1 g806(.A(new_n792), .B(new_n779), .C1(new_n678), .C2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT62), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n690), .B1(new_n834), .B2(new_n835), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n994), .B1(new_n995), .B2(new_n686), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n684), .A2(new_n661), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT97), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n999), .A2(new_n676), .A3(new_n682), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n1000), .A2(KEYINPUT62), .A3(new_n985), .A4(new_n690), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n993), .B1(new_n996), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n972), .B1(new_n1002), .B2(G953), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n981), .A2(new_n987), .ZN(new_n1004));
  INV_X1    g818(.A(new_n979), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1004), .A2(new_n485), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1006), .A2(new_n973), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n991), .B(new_n1008), .ZN(G72));
  NAND2_X1  g823(.A1(new_n1002), .A2(new_n962), .ZN(new_n1010));
  XNOR2_X1  g824(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n491), .A2(new_n190), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1011), .B(new_n1012), .ZN(new_n1013));
  AOI211_X1 g827(.A(new_n516), .B(new_n528), .C1(new_n1010), .C2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n877), .A2(new_n886), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n528), .B(new_n515), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n1013), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n921), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n528), .A2(new_n516), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n988), .A2(new_n962), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1019), .B1(new_n1020), .B2(new_n1013), .ZN(new_n1021));
  NOR3_X1   g835(.A1(new_n1014), .A2(new_n1018), .A3(new_n1021), .ZN(G57));
endmodule


