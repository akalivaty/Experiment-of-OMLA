//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1225, new_n1226, new_n1227, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G77), .A2(G244), .ZN(new_n217));
  INV_X1    g0017(.A(G116), .ZN(new_n218));
  INV_X1    g0018(.A(G270), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n220), .B1(G50), .B2(G226), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  XNOR2_X1  g0022(.A(KEYINPUT64), .B(G68), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n225));
  INV_X1    g0025(.A(G58), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  INV_X1    g0027(.A(G107), .ZN(new_n228));
  INV_X1    g0028(.A(G264), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n225), .B1(new_n226), .B2(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(KEYINPUT65), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n221), .B1(new_n222), .B2(new_n224), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  AND2_X1   g0032(.A1(new_n230), .A2(new_n231), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n208), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n211), .B(new_n216), .C1(new_n234), .C2(KEYINPUT1), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n235), .B1(KEYINPUT1), .B2(new_n234), .ZN(G361));
  XOR2_X1   g0036(.A(G238), .B(G244), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT67), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G226), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n242), .B(new_n246), .ZN(G358));
  XNOR2_X1  g0047(.A(G68), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(new_n226), .ZN(new_n249));
  XOR2_X1   g0049(.A(KEYINPUT68), .B(G50), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n251), .B(new_n254), .Z(G351));
  INV_X1    g0055(.A(G13), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(G1), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G20), .ZN(new_n258));
  INV_X1    g0058(.A(G50), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n214), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n261), .B1(new_n207), .B2(G33), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n262), .B1(G1), .B2(new_n206), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n260), .B1(new_n264), .B2(new_n259), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n265), .B(KEYINPUT71), .ZN(new_n266));
  INV_X1    g0066(.A(new_n262), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT8), .B(G58), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n206), .A2(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n206), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G150), .ZN(new_n273));
  OAI22_X1  g0073(.A1(new_n201), .A2(new_n206), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n267), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n266), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n276), .B(KEYINPUT9), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n271), .A2(KEYINPUT3), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT3), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(G33), .ZN(new_n280));
  OAI21_X1  g0080(.A(KEYINPUT70), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n271), .A2(KEYINPUT3), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT70), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G1698), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(G222), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(G223), .A3(G1698), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n288), .B(new_n289), .C1(new_n202), .C2(new_n286), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n291), .ZN(new_n293));
  INV_X1    g0093(.A(G41), .ZN(new_n294));
  INV_X1    g0094(.A(G45), .ZN(new_n295));
  AOI21_X1  g0095(.A(G1), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT69), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(G41), .A2(G45), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT69), .B1(new_n299), .B2(G1), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n293), .A2(new_n298), .A3(G274), .A4(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n291), .A2(new_n296), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n302), .B1(G226), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n292), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G200), .ZN(new_n306));
  INV_X1    g0106(.A(new_n305), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G190), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n277), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT10), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n276), .B1(new_n307), .B2(G169), .ZN(new_n311));
  INV_X1    g0111(.A(G179), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n311), .B1(new_n312), .B2(new_n307), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(G58), .A2(G68), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n223), .B2(G58), .ZN(new_n317));
  INV_X1    g0117(.A(G159), .ZN(new_n318));
  OAI22_X1  g0118(.A1(new_n317), .A2(new_n206), .B1(new_n318), .B2(new_n272), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n206), .A2(KEYINPUT7), .ZN(new_n320));
  AND2_X1   g0120(.A1(KEYINPUT76), .A2(G33), .ZN(new_n321));
  NOR2_X1   g0121(.A1(KEYINPUT76), .A2(G33), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n279), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n320), .B1(new_n323), .B2(new_n283), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  AND3_X1   g0125(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n284), .B1(new_n282), .B2(new_n283), .ZN(new_n327));
  NOR3_X1   g0127(.A1(new_n326), .A2(new_n327), .A3(G20), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n325), .B1(new_n328), .B2(KEYINPUT7), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n319), .B1(new_n329), .B2(new_n223), .ZN(new_n330));
  XOR2_X1   g0130(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT78), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G68), .ZN(new_n334));
  OR2_X1    g0134(.A1(KEYINPUT76), .A2(G33), .ZN(new_n335));
  NAND2_X1  g0135(.A1(KEYINPUT76), .A2(G33), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(KEYINPUT3), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(G20), .B1(new_n337), .B2(new_n282), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT7), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n334), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n321), .A2(new_n322), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n278), .B1(new_n341), .B2(KEYINPUT3), .ZN(new_n342));
  OAI21_X1  g0142(.A(KEYINPUT7), .B1(new_n342), .B2(G20), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n319), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n262), .B1(new_n344), .B2(KEYINPUT16), .ZN(new_n345));
  INV_X1    g0145(.A(new_n319), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n281), .A2(new_n206), .A3(new_n285), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n324), .B1(new_n347), .B2(new_n339), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n346), .B1(new_n348), .B2(new_n224), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT78), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n349), .A2(new_n350), .A3(new_n331), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n333), .A2(new_n345), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n258), .A2(new_n268), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(new_n264), .B2(new_n268), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n303), .A2(G232), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n301), .A2(new_n355), .ZN(new_n356));
  MUX2_X1   g0156(.A(G223), .B(G226), .S(G1698), .Z(new_n357));
  AOI22_X1  g0157(.A1(new_n342), .A2(new_n357), .B1(G33), .B2(G87), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n356), .B1(new_n293), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G200), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(G190), .B2(new_n359), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n352), .A2(new_n354), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT17), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(KEYINPUT79), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT79), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n352), .A2(new_n367), .A3(new_n354), .A4(new_n362), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n365), .B1(new_n369), .B2(KEYINPUT17), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n359), .A2(G169), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n356), .B(G179), .C1(new_n293), .C2(new_n358), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  AND3_X1   g0174(.A1(new_n349), .A2(new_n350), .A3(new_n331), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n350), .B1(new_n349), .B2(new_n331), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n337), .A2(new_n282), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n377), .A2(new_n339), .A3(new_n206), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(G68), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n338), .A2(new_n339), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n346), .B(KEYINPUT16), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n267), .ZN(new_n382));
  NOR3_X1   g0182(.A1(new_n375), .A2(new_n376), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n354), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n374), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT18), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n373), .B1(new_n352), .B2(new_n354), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT18), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n370), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n223), .A2(new_n206), .ZN(new_n392));
  OAI22_X1  g0192(.A1(new_n272), .A2(new_n259), .B1(new_n269), .B2(new_n202), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n267), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  XNOR2_X1  g0194(.A(new_n394), .B(KEYINPUT11), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n392), .A2(KEYINPUT12), .A3(new_n257), .ZN(new_n396));
  INV_X1    g0196(.A(new_n258), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n396), .B1(KEYINPUT12), .B2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n334), .B1(new_n263), .B2(KEYINPUT12), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  XOR2_X1   g0201(.A(new_n401), .B(KEYINPUT74), .Z(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT13), .ZN(new_n404));
  NOR2_X1   g0204(.A1(G226), .A2(G1698), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n405), .B1(new_n227), .B2(G1698), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n286), .A2(new_n406), .B1(G33), .B2(G97), .ZN(new_n407));
  OR2_X1    g0207(.A1(new_n407), .A2(new_n293), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n302), .B1(G238), .B2(new_n303), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n404), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n408), .A2(new_n404), .A3(new_n409), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(G190), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(G200), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n403), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(G169), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT14), .B1(new_n414), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT75), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n414), .A2(new_n421), .A3(G179), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT14), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n413), .A2(new_n423), .A3(G169), .ZN(new_n424));
  OAI21_X1  g0224(.A(KEYINPUT75), .B1(new_n413), .B2(new_n312), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n420), .A2(new_n422), .A3(new_n424), .A4(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n418), .B1(new_n426), .B2(new_n402), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n326), .A2(new_n327), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n293), .B1(new_n428), .B2(new_n228), .ZN(new_n429));
  NOR2_X1   g0229(.A1(G232), .A2(G1698), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n430), .B1(new_n222), .B2(G1698), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n429), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n302), .B1(G244), .B2(new_n303), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n434), .A2(G179), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n435), .B1(new_n419), .B2(new_n434), .ZN(new_n436));
  XNOR2_X1  g0236(.A(KEYINPUT15), .B(G87), .ZN(new_n437));
  OAI22_X1  g0237(.A1(new_n437), .A2(new_n269), .B1(new_n206), .B2(new_n202), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n268), .A2(new_n272), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n267), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  XOR2_X1   g0240(.A(new_n440), .B(KEYINPUT72), .Z(new_n441));
  NAND2_X1  g0241(.A1(new_n264), .A2(G77), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n441), .B(new_n442), .C1(G77), .C2(new_n258), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n436), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  XNOR2_X1  g0245(.A(new_n443), .B(KEYINPUT73), .ZN(new_n446));
  INV_X1    g0246(.A(G190), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n434), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n448), .B1(G200), .B2(new_n434), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n445), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n427), .A2(new_n450), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n315), .A2(new_n391), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT25), .B1(new_n397), .B2(new_n228), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n397), .A2(KEYINPUT25), .A3(new_n228), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n205), .A2(G33), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n262), .A2(new_n258), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n454), .A2(new_n455), .B1(new_n458), .B2(G107), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  OR3_X1    g0260(.A1(new_n206), .A2(KEYINPUT23), .A3(G107), .ZN(new_n461));
  OAI21_X1  g0261(.A(KEYINPUT23), .B1(new_n206), .B2(G107), .ZN(new_n462));
  INV_X1    g0262(.A(new_n341), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G116), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n461), .B(new_n462), .C1(new_n464), .C2(G20), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n342), .A2(new_n206), .ZN(new_n466));
  INV_X1    g0266(.A(G87), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT22), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n467), .A2(KEYINPUT22), .A3(G20), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n286), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n465), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT24), .ZN(new_n472));
  XNOR2_X1  g0272(.A(new_n471), .B(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n460), .B1(new_n473), .B2(new_n267), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT86), .ZN(new_n476));
  NOR2_X1   g0276(.A1(G250), .A2(G1698), .ZN(new_n477));
  INV_X1    g0277(.A(G257), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n477), .B1(new_n478), .B2(G1698), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n342), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT85), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n463), .A2(G294), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n481), .B1(new_n480), .B2(new_n482), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n483), .A2(new_n484), .A3(new_n293), .ZN(new_n485));
  XNOR2_X1  g0285(.A(KEYINPUT5), .B(G41), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n295), .A2(G1), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n293), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(new_n229), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n476), .B1(new_n485), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n484), .A2(new_n293), .ZN(new_n492));
  INV_X1    g0292(.A(new_n483), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n490), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n494), .A2(KEYINPUT86), .A3(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n293), .A2(G274), .A3(new_n487), .A4(new_n486), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n491), .A2(new_n496), .A3(G179), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n494), .A2(new_n495), .ZN(new_n499));
  INV_X1    g0299(.A(new_n497), .ZN(new_n500));
  OAI21_X1  g0300(.A(G169), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n475), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n491), .A2(new_n496), .A3(new_n497), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n504), .A2(new_n360), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n499), .A2(G190), .A3(new_n500), .ZN(new_n506));
  OAI211_X1 g0306(.A(KEYINPUT87), .B(new_n474), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT87), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n506), .B1(new_n360), .B2(new_n504), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n508), .B1(new_n509), .B2(new_n475), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT84), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT21), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n458), .A2(G116), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n397), .A2(new_n218), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n206), .A2(G116), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n262), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G33), .A2(G283), .ZN(new_n518));
  INV_X1    g0318(.A(G97), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n518), .B(new_n206), .C1(G33), .C2(new_n519), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n517), .A2(KEYINPUT20), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT20), .B1(new_n517), .B2(new_n520), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n514), .B(new_n515), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G169), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n428), .A2(G303), .ZN(new_n525));
  NOR2_X1   g0325(.A1(G257), .A2(G1698), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n526), .B1(new_n229), .B2(G1698), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n342), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n293), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n497), .B1(new_n489), .B2(new_n219), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n512), .B(new_n513), .C1(new_n524), .C2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT83), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(G179), .ZN(new_n534));
  INV_X1    g0334(.A(new_n523), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n531), .A2(new_n523), .A3(KEYINPUT83), .A4(G179), .ZN(new_n537));
  INV_X1    g0337(.A(new_n531), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n512), .A2(new_n513), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n538), .A2(G169), .A3(new_n539), .A4(new_n523), .ZN(new_n540));
  AND4_X1   g0340(.A1(new_n532), .A2(new_n536), .A3(new_n537), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n487), .A2(G274), .ZN(new_n542));
  OAI21_X1  g0342(.A(G250), .B1(new_n295), .B2(G1), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n542), .B1(new_n291), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n342), .A2(G238), .A3(new_n287), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n342), .A2(G244), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n545), .B(new_n464), .C1(new_n546), .C2(new_n287), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n544), .B1(new_n547), .B2(new_n291), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G200), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT82), .ZN(new_n551));
  AOI21_X1  g0351(.A(G20), .B1(G33), .B2(G97), .ZN(new_n552));
  NOR2_X1   g0352(.A1(G97), .A2(G107), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n552), .B1(new_n467), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT19), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G97), .ZN(new_n556));
  OAI22_X1  g0356(.A1(new_n554), .A2(new_n555), .B1(new_n269), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(new_n466), .B2(new_n334), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n558), .A2(new_n267), .B1(new_n397), .B2(new_n437), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n458), .A2(G87), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n550), .A2(new_n551), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n548), .A2(new_n360), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n559), .A2(new_n560), .ZN(new_n563));
  OAI21_X1  g0363(.A(KEYINPUT82), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n548), .A2(G190), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n561), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n523), .B1(new_n538), .B2(G200), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n447), .B2(new_n538), .ZN(new_n568));
  OR2_X1    g0368(.A1(new_n457), .A2(new_n437), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n548), .A2(new_n312), .B1(new_n559), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(G169), .B2(new_n548), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n541), .A2(new_n566), .A3(new_n568), .A4(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n272), .A2(new_n202), .ZN(new_n573));
  XOR2_X1   g0373(.A(new_n573), .B(KEYINPUT80), .Z(new_n574));
  NAND3_X1  g0374(.A1(new_n228), .A2(KEYINPUT6), .A3(G97), .ZN(new_n575));
  XOR2_X1   g0375(.A(G97), .B(G107), .Z(new_n576));
  OAI21_X1  g0376(.A(new_n575), .B1(new_n576), .B2(KEYINPUT6), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n574), .B1(G20), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n329), .A2(G107), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n262), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n397), .A2(new_n519), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n457), .B2(new_n519), .ZN(new_n582));
  OR2_X1    g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n497), .B1(new_n489), .B2(new_n478), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT4), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n546), .B2(G1698), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n286), .A2(KEYINPUT4), .A3(G244), .A4(new_n287), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n286), .A2(G250), .A3(G1698), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .A4(new_n518), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n584), .B1(new_n589), .B2(new_n291), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n590), .A2(new_n419), .ZN(new_n591));
  AOI211_X1 g0391(.A(new_n312), .B(new_n584), .C1(new_n589), .C2(new_n291), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n583), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n590), .A2(G190), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n580), .A2(new_n582), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n594), .B(new_n595), .C1(new_n360), .C2(new_n590), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT81), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n593), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n597), .B1(new_n593), .B2(new_n596), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n572), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  AND4_X1   g0400(.A1(new_n452), .A2(new_n503), .A3(new_n511), .A4(new_n600), .ZN(G372));
  NAND2_X1  g0401(.A1(new_n426), .A2(new_n402), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n418), .B2(new_n444), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n603), .A2(new_n370), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT89), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n352), .A2(new_n354), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT18), .B1(new_n606), .B2(new_n374), .ZN(new_n607));
  AOI211_X1 g0407(.A(new_n386), .B(new_n373), .C1(new_n352), .C2(new_n354), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n605), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n387), .A2(KEYINPUT89), .A3(new_n389), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n310), .B1(new_n604), .B2(new_n612), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n613), .A2(new_n314), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n590), .A2(G179), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n419), .B2(new_n590), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n566), .A2(new_n583), .A3(new_n616), .A4(new_n571), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(KEYINPUT26), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT88), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n595), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n550), .A2(new_n559), .A3(new_n560), .A4(new_n565), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n621), .A2(new_n571), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT26), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n615), .B(KEYINPUT88), .C1(new_n419), .C2(new_n590), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n620), .A2(new_n622), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n618), .A2(new_n625), .A3(new_n571), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n503), .A2(new_n541), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n593), .A2(new_n596), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n628), .A2(new_n622), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n511), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n452), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n614), .A2(new_n632), .ZN(G369));
  NAND2_X1  g0433(.A1(new_n257), .A2(new_n206), .ZN(new_n634));
  OR2_X1    g0434(.A1(new_n634), .A2(KEYINPUT27), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(KEYINPUT27), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(new_n636), .A3(G213), .ZN(new_n637));
  INV_X1    g0437(.A(G343), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n541), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n474), .B1(new_n501), .B2(new_n498), .ZN(new_n642));
  INV_X1    g0442(.A(new_n639), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n474), .A2(new_n643), .ZN(new_n644));
  AOI211_X1 g0444(.A(new_n642), .B(new_n644), .C1(new_n507), .C2(new_n510), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n503), .A2(new_n643), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT90), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n644), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n511), .A2(new_n503), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT90), .ZN(new_n650));
  INV_X1    g0450(.A(new_n646), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n641), .B1(new_n647), .B2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n503), .A2(new_n639), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n647), .A2(new_n652), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n523), .A2(new_n639), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n541), .A2(new_n568), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n541), .B2(new_n657), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G330), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n655), .A2(new_n662), .ZN(G399));
  INV_X1    g0463(.A(new_n209), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(G41), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n553), .A2(new_n467), .A3(new_n218), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n666), .A2(G1), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(new_n212), .B2(new_n666), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT28), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n571), .B1(new_n617), .B2(KEYINPUT26), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n620), .A2(new_n622), .A3(new_n624), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n672), .B1(KEYINPUT26), .B2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT92), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n627), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n511), .A2(new_n629), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n674), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n678), .A2(KEYINPUT29), .A3(new_n643), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n631), .A2(new_n643), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT29), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n600), .A2(new_n503), .A3(new_n511), .A4(new_n643), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT30), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n534), .A2(KEYINPUT91), .ZN(new_n685));
  NOR4_X1   g0485(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT91), .A4(new_n312), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n685), .A2(new_n590), .A3(new_n687), .A4(new_n548), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n491), .A2(new_n496), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n684), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n491), .A2(new_n496), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT91), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n692), .B1(new_n531), .B2(G179), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n693), .A2(new_n686), .A3(new_n549), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n691), .A2(new_n694), .A3(KEYINPUT30), .A4(new_n590), .ZN(new_n695));
  NOR4_X1   g0495(.A1(new_n590), .A2(G179), .A3(new_n531), .A4(new_n548), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n504), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n690), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  AND3_X1   g0498(.A1(new_n698), .A2(KEYINPUT31), .A3(new_n639), .ZN(new_n699));
  AOI21_X1  g0499(.A(KEYINPUT31), .B1(new_n698), .B2(new_n639), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n683), .A2(new_n701), .ZN(new_n702));
  AOI22_X1  g0502(.A1(new_n679), .A2(new_n682), .B1(G330), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n671), .B1(new_n703), .B2(G1), .ZN(G364));
  NOR2_X1   g0504(.A1(new_n256), .A2(G20), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n205), .B1(new_n705), .B2(G45), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n665), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n286), .A2(new_n209), .ZN(new_n709));
  INV_X1    g0509(.A(G355), .ZN(new_n710));
  OAI22_X1  g0510(.A1(new_n709), .A2(new_n710), .B1(G116), .B2(new_n209), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n251), .A2(G45), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n377), .A2(new_n209), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n713), .B1(new_n295), .B2(new_n213), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n711), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(G13), .A2(G33), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(G20), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n214), .B1(G20), .B2(new_n419), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n708), .B1(new_n715), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n206), .A2(new_n447), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n312), .A2(G200), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n206), .A2(G190), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  AOI22_X1  g0529(.A1(G58), .A2(new_n726), .B1(new_n729), .B2(G77), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n312), .A2(new_n360), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n723), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n730), .B1(new_n259), .B2(new_n732), .ZN(new_n733));
  XOR2_X1   g0533(.A(new_n733), .B(KEYINPUT93), .Z(new_n734));
  NAND2_X1  g0534(.A1(new_n731), .A2(new_n727), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n360), .A2(G179), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n723), .A2(new_n736), .ZN(new_n737));
  OAI22_X1  g0537(.A1(new_n334), .A2(new_n735), .B1(new_n737), .B2(new_n467), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n727), .A2(new_n736), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n738), .B1(G107), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G179), .A2(G200), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n727), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n318), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT32), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n206), .B1(new_n742), .B2(G190), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G97), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n741), .A2(new_n745), .A3(new_n286), .A4(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n734), .A2(new_n749), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n750), .A2(KEYINPUT94), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(KEYINPUT94), .ZN(new_n752));
  INV_X1    g0552(.A(G303), .ZN(new_n753));
  INV_X1    g0553(.A(G283), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n737), .A2(new_n753), .B1(new_n739), .B2(new_n754), .ZN(new_n755));
  AOI211_X1 g0555(.A(new_n286), .B(new_n755), .C1(G294), .C2(new_n747), .ZN(new_n756));
  XOR2_X1   g0556(.A(KEYINPUT33), .B(G317), .Z(new_n757));
  INV_X1    g0557(.A(G322), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n757), .A2(new_n735), .B1(new_n725), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT95), .ZN(new_n760));
  INV_X1    g0560(.A(G326), .ZN(new_n761));
  INV_X1    g0561(.A(G311), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n732), .A2(new_n761), .B1(new_n728), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n743), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n763), .B1(G329), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n756), .A2(new_n760), .A3(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n751), .A2(new_n752), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n722), .B1(new_n767), .B2(new_n719), .ZN(new_n768));
  INV_X1    g0568(.A(new_n718), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n768), .B1(new_n659), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n708), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n660), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n659), .A2(G330), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n770), .B1(new_n772), .B2(new_n773), .ZN(G396));
  NOR2_X1   g0574(.A1(new_n444), .A2(new_n643), .ZN(new_n775));
  OR2_X1    g0575(.A1(new_n775), .A2(KEYINPUT97), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(KEYINPUT97), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n443), .A2(new_n639), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n776), .A2(new_n777), .B1(new_n450), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n680), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n639), .B1(new_n626), .B2(new_n630), .ZN(new_n781));
  INV_X1    g0581(.A(new_n779), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n702), .A2(G330), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n708), .B(new_n786), .C1(KEYINPUT98), .C2(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n788), .B1(KEYINPUT98), .B2(new_n787), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n719), .A2(new_n716), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n708), .B1(G77), .B2(new_n791), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT96), .Z(new_n793));
  INV_X1    g0593(.A(new_n719), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n739), .A2(new_n334), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n795), .B1(G132), .B2(new_n764), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(new_n259), .B2(new_n737), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n377), .B(new_n797), .C1(G58), .C2(new_n747), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n735), .A2(new_n273), .ZN(new_n799));
  INV_X1    g0599(.A(G143), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n725), .A2(new_n800), .B1(new_n728), .B2(new_n318), .ZN(new_n801));
  INV_X1    g0601(.A(new_n732), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n799), .B(new_n801), .C1(G137), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(KEYINPUT34), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n803), .A2(KEYINPUT34), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n798), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n739), .A2(new_n467), .ZN(new_n807));
  INV_X1    g0607(.A(G294), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n754), .A2(new_n735), .B1(new_n725), .B2(new_n808), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n807), .B(new_n809), .C1(G311), .C2(new_n764), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n732), .A2(new_n753), .B1(new_n737), .B2(new_n228), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(G116), .B2(new_n729), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n810), .A2(new_n428), .A3(new_n748), .A4(new_n812), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n806), .A2(new_n813), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n793), .B1(new_n794), .B2(new_n814), .C1(new_n782), .C2(new_n717), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n789), .A2(new_n815), .ZN(G384));
  OR2_X1    g0616(.A1(new_n577), .A2(KEYINPUT35), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n577), .A2(KEYINPUT35), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n817), .A2(G116), .A3(new_n215), .A4(new_n818), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT36), .Z(new_n820));
  OAI211_X1 g0620(.A(G77), .B(new_n213), .C1(new_n224), .C2(new_n226), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n259), .A2(G68), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n205), .B(G13), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n369), .ZN(new_n825));
  INV_X1    g0625(.A(new_n637), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n383), .B2(new_n384), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT102), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n606), .A2(KEYINPUT102), .A3(new_n826), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n388), .A2(KEYINPUT37), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n825), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n344), .A2(new_n332), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n354), .B1(new_n382), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(KEYINPUT100), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n373), .A2(new_n637), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT100), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n838), .B(new_n354), .C1(new_n382), .C2(new_n834), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n836), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n366), .A2(new_n368), .A3(new_n840), .ZN(new_n841));
  AND3_X1   g0641(.A1(new_n841), .A2(KEYINPUT101), .A3(KEYINPUT37), .ZN(new_n842));
  AOI21_X1  g0642(.A(KEYINPUT101), .B1(new_n841), .B2(KEYINPUT37), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n833), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(KEYINPUT103), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT103), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n846), .B(new_n833), .C1(new_n842), .C2(new_n843), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n836), .A2(new_n826), .A3(new_n839), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(new_n370), .B2(new_n390), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n848), .A2(KEYINPUT38), .A3(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT38), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n385), .A2(new_n605), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n388), .A2(KEYINPUT89), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n854), .A2(new_n363), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT102), .B1(new_n606), .B2(new_n826), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n828), .B(new_n637), .C1(new_n352), .C2(new_n354), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(KEYINPUT37), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT104), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n825), .A2(new_n831), .A3(new_n861), .A4(new_n832), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT37), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n366), .A2(new_n863), .A3(new_n385), .A4(new_n368), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT104), .B1(new_n859), .B2(new_n864), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n860), .A2(new_n862), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n831), .B1(new_n611), .B2(new_n370), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n853), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n852), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n779), .B1(new_n683), .B2(new_n701), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n427), .B1(new_n403), .B2(new_n643), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT99), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n403), .A2(new_n643), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n426), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n872), .B1(new_n426), .B2(new_n873), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n871), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n870), .A2(new_n877), .A3(KEYINPUT40), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n869), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n870), .A2(new_n877), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n841), .A2(KEYINPUT37), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT101), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n841), .A2(KEYINPUT101), .A3(KEYINPUT37), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n846), .B1(new_n886), .B2(new_n833), .ZN(new_n887));
  INV_X1    g0687(.A(new_n847), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n851), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n853), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n881), .B1(new_n890), .B2(new_n852), .ZN(new_n891));
  OAI211_X1 g0691(.A(G330), .B(new_n880), .C1(new_n891), .C2(KEYINPUT40), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n452), .A2(G330), .A3(new_n702), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n894), .B(KEYINPUT106), .Z(new_n895));
  AOI21_X1  g0695(.A(new_n878), .B1(new_n852), .B2(new_n868), .ZN(new_n896));
  INV_X1    g0696(.A(new_n881), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT38), .B1(new_n848), .B2(new_n851), .ZN(new_n898));
  AOI211_X1 g0698(.A(new_n853), .B(new_n850), .C1(new_n845), .C2(new_n847), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT40), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n896), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n902), .A2(new_n452), .A3(new_n702), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n895), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(KEYINPUT39), .B1(new_n898), .B2(new_n899), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT105), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT39), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n868), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n906), .B1(new_n899), .B2(new_n908), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n852), .A2(KEYINPUT105), .A3(new_n907), .A4(new_n868), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n905), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n602), .A2(new_n639), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n444), .A2(new_n639), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n781), .B2(new_n782), .ZN(new_n915));
  INV_X1    g0715(.A(new_n877), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n898), .B2(new_n899), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n612), .A2(new_n637), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n913), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n679), .A2(new_n682), .A3(new_n452), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n614), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n922), .B(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n904), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n205), .B2(new_n705), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n904), .A2(new_n925), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n824), .B1(new_n927), .B2(new_n928), .ZN(G367));
  OAI221_X1 g0729(.A(new_n720), .B1(new_n209), .B2(new_n437), .C1(new_n246), .C2(new_n713), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n930), .A2(new_n708), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n725), .A2(new_n753), .B1(new_n739), .B2(new_n519), .ZN(new_n932));
  OAI22_X1  g0732(.A1(new_n735), .A2(new_n808), .B1(new_n728), .B2(new_n754), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XOR2_X1   g0734(.A(KEYINPUT111), .B(G311), .Z(new_n935));
  INV_X1    g0735(.A(G317), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n732), .A2(new_n935), .B1(new_n936), .B2(new_n743), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n937), .A2(new_n342), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n737), .A2(new_n218), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n939), .A2(KEYINPUT46), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n939), .A2(KEYINPUT46), .B1(G107), .B2(new_n747), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n934), .A2(new_n938), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  AOI22_X1  g0742(.A1(G143), .A2(new_n802), .B1(new_n726), .B2(G150), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n334), .B2(new_n746), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT112), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(G137), .ZN(new_n947));
  OAI22_X1  g0747(.A1(new_n737), .A2(new_n226), .B1(new_n743), .B2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n735), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n948), .B1(G159), .B2(new_n949), .ZN(new_n950));
  AOI22_X1  g0750(.A1(G50), .A2(new_n729), .B1(new_n740), .B2(G77), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n946), .A2(new_n286), .A3(new_n950), .A4(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n944), .A2(new_n945), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n942), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT47), .Z(new_n955));
  NAND2_X1  g0755(.A1(new_n563), .A2(new_n639), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n622), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n571), .B2(new_n956), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n931), .B1(new_n794), .B2(new_n955), .C1(new_n958), .C2(new_n769), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT109), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n958), .B(KEYINPUT43), .Z(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT107), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT42), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n628), .B1(new_n595), .B2(new_n643), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n620), .A2(new_n624), .A3(new_n639), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n964), .B1(new_n653), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n642), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n639), .B1(new_n969), .B2(new_n593), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n963), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  NOR3_X1   g0771(.A1(new_n645), .A2(KEYINPUT90), .A3(new_n646), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n650), .B1(new_n649), .B2(new_n651), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n640), .B(new_n967), .C1(new_n972), .C2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(KEYINPUT42), .ZN(new_n975));
  INV_X1    g0775(.A(new_n970), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n975), .A2(KEYINPUT107), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n971), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n653), .A2(new_n964), .A3(new_n967), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n962), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n981));
  AOI21_X1  g0781(.A(KEYINPUT107), .B1(new_n975), .B2(new_n976), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n963), .B(new_n970), .C1(new_n974), .C2(KEYINPUT42), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n981), .B(new_n979), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT108), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n978), .A2(KEYINPUT108), .A3(new_n981), .A4(new_n979), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n980), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n967), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n662), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n960), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n988), .A2(new_n990), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n665), .B(KEYINPUT41), .Z(new_n993));
  NOR3_X1   g0793(.A1(new_n972), .A2(new_n973), .A3(new_n640), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n660), .B1(new_n994), .B2(new_n653), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n640), .B1(new_n972), .B2(new_n973), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n647), .A2(new_n652), .A3(new_n641), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n996), .A2(new_n661), .A3(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n995), .A2(new_n703), .A3(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT110), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT44), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n655), .B2(new_n967), .ZN(new_n1003));
  OAI211_X1 g0803(.A(KEYINPUT44), .B(new_n989), .C1(new_n653), .C2(new_n654), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n655), .A2(KEYINPUT45), .A3(new_n967), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n654), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n996), .A2(new_n1007), .A3(new_n967), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT45), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1005), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n662), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1005), .A2(new_n1011), .A3(new_n662), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1001), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n993), .B1(new_n1016), .B2(new_n703), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n991), .B(new_n992), .C1(new_n1017), .C2(new_n707), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n988), .A2(new_n960), .A3(new_n990), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n959), .B1(new_n1018), .B2(new_n1019), .ZN(G387));
  NAND2_X1  g0820(.A1(new_n995), .A2(new_n998), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n707), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n656), .A2(new_n769), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n268), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G50), .A2(new_n726), .B1(new_n949), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n318), .B2(new_n732), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT113), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n737), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(G77), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n273), .B2(new_n743), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1027), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n746), .A2(new_n437), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n334), .A2(new_n728), .B1(new_n739), .B2(new_n519), .ZN(new_n1035));
  NOR4_X1   g0835(.A1(new_n1033), .A2(new_n377), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n739), .A2(new_n218), .B1(new_n743), .B2(new_n761), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G322), .A2(new_n802), .B1(new_n726), .B2(G317), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n935), .A2(new_n735), .B1(new_n728), .B2(new_n753), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n1041), .A2(KEYINPUT48), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1041), .A2(KEYINPUT48), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n737), .A2(new_n808), .B1(new_n746), .B2(new_n754), .ZN(new_n1044));
  NOR3_X1   g0844(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n342), .B(new_n1037), .C1(new_n1045), .C2(KEYINPUT49), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1045), .A2(KEYINPUT49), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1036), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n242), .A2(new_n295), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n1049), .A2(new_n713), .B1(new_n668), .B2(new_n709), .ZN(new_n1050));
  OR3_X1    g0850(.A1(new_n268), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1051));
  OAI21_X1  g0851(.A(KEYINPUT50), .B1(new_n268), .B2(G50), .ZN(new_n1052));
  AOI21_X1  g0852(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1051), .A2(new_n668), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n1050), .A2(new_n1054), .B1(new_n228), .B2(new_n664), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n708), .B1(new_n1048), .B2(new_n794), .C1(new_n1055), .C2(new_n721), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n665), .B(KEYINPUT114), .Z(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n1022), .B2(new_n703), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1023), .B1(new_n1024), .B2(new_n1056), .C1(new_n1001), .C2(new_n1058), .ZN(G393));
  INV_X1    g0859(.A(new_n1057), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1015), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n662), .B1(new_n1005), .B2(new_n1011), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1060), .B1(new_n1063), .B2(new_n1001), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n1001), .B2(new_n1063), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n989), .A2(new_n718), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n720), .B1(new_n519), .B2(new_n209), .C1(new_n254), .C2(new_n713), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n708), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n737), .A2(new_n754), .B1(new_n743), .B2(new_n758), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT115), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n228), .A2(new_n739), .B1(new_n728), .B2(new_n808), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(G303), .B2(new_n949), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n286), .B1(G116), .B2(new_n747), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1070), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n732), .A2(new_n936), .B1(new_n725), .B2(new_n762), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n1075), .B(KEYINPUT52), .Z(new_n1076));
  OAI22_X1  g0876(.A1(new_n732), .A2(new_n273), .B1(new_n725), .B2(new_n318), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT51), .Z(new_n1078));
  OAI22_X1  g0878(.A1(new_n735), .A2(new_n259), .B1(new_n743), .B2(new_n800), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n223), .B2(new_n1029), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n747), .A2(G77), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n807), .B1(new_n1025), .B2(new_n729), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1080), .A2(new_n342), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n1074), .A2(new_n1076), .B1(new_n1078), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1068), .B1(new_n1084), .B2(new_n719), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n1063), .A2(new_n707), .B1(new_n1066), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1065), .A2(new_n1086), .ZN(G390));
  NAND3_X1  g0887(.A1(new_n614), .A2(new_n923), .A3(new_n893), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n702), .A2(G330), .A3(new_n782), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n916), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n870), .A2(new_n877), .A3(G330), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n678), .A2(new_n643), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n914), .B1(new_n1095), .B2(new_n782), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n915), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(KEYINPUT116), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1098), .A2(KEYINPUT116), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1089), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n912), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n915), .B2(new_n916), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n905), .A2(new_n909), .A3(new_n910), .A4(new_n1104), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n869), .B(new_n1103), .C1(new_n1096), .C2(new_n916), .ZN(new_n1106));
  AND3_X1   g0906(.A1(new_n1105), .A2(new_n1092), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1092), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1102), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1092), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1094), .A2(new_n1096), .B1(new_n1098), .B2(KEYINPUT116), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n915), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1093), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT116), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1088), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1105), .A2(new_n1092), .A3(new_n1106), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1112), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1109), .A2(new_n1120), .A3(new_n1057), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n911), .A2(new_n717), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n725), .A2(new_n218), .B1(new_n743), .B2(new_n808), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n795), .B(new_n1123), .C1(G87), .C2(new_n1029), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n735), .A2(new_n228), .B1(new_n728), .B2(new_n519), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(G283), .B2(new_n802), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1124), .A2(new_n428), .A3(new_n1081), .A4(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(G125), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n286), .B1(new_n259), .B2(new_n739), .C1(new_n1128), .C2(new_n743), .ZN(new_n1129));
  XOR2_X1   g0929(.A(new_n1129), .B(KEYINPUT117), .Z(new_n1130));
  XNOR2_X1  g0930(.A(KEYINPUT54), .B(G143), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n802), .A2(G128), .B1(new_n729), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(G132), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n1133), .B1(new_n1134), .B2(new_n725), .C1(new_n947), .C2(new_n735), .ZN(new_n1135));
  OR3_X1    g0935(.A1(new_n737), .A2(KEYINPUT53), .A3(new_n273), .ZN(new_n1136));
  OAI21_X1  g0936(.A(KEYINPUT53), .B1(new_n737), .B2(new_n273), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1136), .B(new_n1137), .C1(new_n318), .C2(new_n746), .ZN(new_n1138));
  OR2_X1    g0938(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1127), .B1(new_n1130), .B2(new_n1139), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n1140), .A2(new_n719), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n708), .B1(new_n1025), .B2(new_n791), .ZN(new_n1142));
  NOR3_X1   g0942(.A1(new_n1122), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1143), .B1(new_n1144), .B2(new_n707), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1121), .A2(new_n1145), .ZN(G378));
  NAND2_X1  g0946(.A1(new_n276), .A2(new_n826), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n1147), .B(KEYINPUT55), .Z(new_n1148));
  XOR2_X1   g0948(.A(new_n315), .B(new_n1148), .Z(new_n1149));
  XOR2_X1   g0949(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n1150));
  XNOR2_X1  g0950(.A(new_n1149), .B(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n892), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1151), .B1(new_n902), .B2(G330), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n922), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n892), .A2(new_n1152), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n920), .B1(new_n911), .B2(new_n912), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n902), .A2(G330), .A3(new_n1151), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1155), .A2(new_n707), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n771), .B1(new_n259), .B2(new_n790), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n735), .A2(new_n1134), .B1(new_n728), .B2(new_n947), .ZN(new_n1162));
  XOR2_X1   g0962(.A(new_n1162), .B(KEYINPUT119), .Z(new_n1163));
  NOR2_X1   g0963(.A1(new_n746), .A2(new_n273), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n732), .A2(new_n1128), .B1(new_n737), .B2(new_n1131), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1164), .B(new_n1165), .C1(G128), .C2(new_n726), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1167), .A2(KEYINPUT59), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1167), .A2(KEYINPUT59), .ZN(new_n1169));
  AOI211_X1 g0969(.A(G33), .B(G41), .C1(new_n764), .C2(G124), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n318), .B2(new_n739), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n1168), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1030), .B1(new_n754), .B2(new_n743), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n735), .A2(new_n519), .B1(new_n739), .B2(new_n226), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n725), .A2(new_n228), .B1(new_n728), .B2(new_n437), .ZN(new_n1175));
  NOR3_X1   g0975(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n732), .A2(new_n218), .B1(new_n746), .B2(new_n334), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT118), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1176), .A2(new_n294), .A3(new_n377), .A4(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(KEYINPUT58), .ZN(new_n1181));
  AOI21_X1  g0981(.A(G50), .B1(new_n271), .B2(new_n294), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n342), .B2(G41), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1180), .A2(KEYINPUT58), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1172), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1161), .B1(new_n794), .B2(new_n1186), .C1(new_n1152), .C2(new_n717), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1160), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1088), .B1(new_n1144), .B2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1155), .A2(KEYINPUT57), .A3(new_n1159), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1057), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1157), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1120), .A2(new_n1089), .ZN(new_n1197));
  AOI21_X1  g0997(.A(KEYINPUT57), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1189), .B1(new_n1193), .B2(new_n1198), .ZN(G375));
  INV_X1    g0999(.A(new_n993), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1117), .A2(new_n1097), .A3(new_n1088), .A4(new_n1099), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1102), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n877), .A2(new_n717), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT121), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n708), .B1(G68), .B2(new_n791), .ZN(new_n1205));
  XOR2_X1   g1005(.A(new_n1205), .B(KEYINPUT122), .Z(new_n1206));
  AOI22_X1  g1006(.A1(G77), .A2(new_n740), .B1(new_n764), .B2(G303), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1207), .B1(new_n228), .B2(new_n728), .C1(new_n754), .C2(new_n725), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(G294), .A2(new_n802), .B1(new_n949), .B2(G116), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n519), .B2(new_n737), .ZN(new_n1210));
  NOR4_X1   g1010(.A1(new_n1208), .A2(new_n1210), .A3(new_n286), .A4(new_n1034), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1212), .A2(KEYINPUT123), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(KEYINPUT123), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n947), .A2(new_n725), .B1(new_n737), .B2(new_n318), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G150), .B2(new_n729), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n949), .A2(new_n1132), .B1(new_n740), .B2(G58), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n802), .A2(G132), .B1(new_n764), .B2(G128), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n377), .B1(G50), .B2(new_n747), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1213), .A2(new_n1214), .A3(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1206), .B1(new_n1221), .B2(new_n719), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1190), .A2(new_n707), .B1(new_n1204), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1202), .A2(new_n1223), .ZN(G381));
  INV_X1    g1024(.A(G378), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1225), .B(new_n1189), .C1(new_n1193), .C2(new_n1198), .ZN(new_n1226));
  OR4_X1    g1026(.A1(G396), .A2(G381), .A3(G393), .A4(G384), .ZN(new_n1227));
  OR4_X1    g1027(.A1(G387), .A2(new_n1226), .A3(new_n1227), .A4(G390), .ZN(G407));
  OAI211_X1 g1028(.A(G407), .B(G213), .C1(G343), .C2(new_n1226), .ZN(G409));
  INV_X1    g1029(.A(G390), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(G387), .A2(new_n1230), .ZN(new_n1231));
  OAI211_X1 g1031(.A(G390), .B(new_n959), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT124), .B1(G387), .B2(new_n1230), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(G393), .B(G396), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1233), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1235), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1231), .A2(KEYINPUT124), .A3(new_n1232), .A4(new_n1237), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1236), .A2(new_n1238), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1121), .A2(new_n1145), .A3(new_n1160), .A4(new_n1187), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1155), .A2(new_n1159), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(new_n1191), .A2(new_n1241), .A3(new_n993), .ZN(new_n1242));
  INV_X1    g1042(.A(G213), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n1240), .A2(new_n1242), .B1(new_n1243), .B2(G343), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G378), .B2(G375), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT60), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1201), .A2(new_n1246), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1113), .A2(new_n1117), .A3(KEYINPUT60), .A4(new_n1088), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1247), .A2(new_n1102), .A3(new_n1057), .A4(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n1223), .ZN(new_n1250));
  INV_X1    g1050(.A(G384), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(G384), .A2(new_n1249), .A3(new_n1223), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1245), .A2(KEYINPUT63), .A3(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT63), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1243), .A2(G343), .ZN(new_n1258));
  AND4_X1   g1058(.A1(new_n1121), .A2(new_n1145), .A3(new_n1160), .A4(new_n1187), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1196), .A2(new_n1200), .A3(new_n1197), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1258), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT57), .ZN(new_n1262));
  NOR3_X1   g1062(.A1(new_n1194), .A2(new_n1195), .A3(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1060), .B1(new_n1263), .B2(new_n1197), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1262), .B1(new_n1191), .B2(new_n1241), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1188), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1261), .B1(new_n1266), .B2(new_n1225), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1257), .B1(new_n1267), .B2(new_n1254), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1258), .A2(G2897), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(new_n1254), .B(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(KEYINPUT61), .B1(new_n1267), .B2(new_n1270), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1239), .A2(new_n1256), .A3(new_n1268), .A4(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT125), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT62), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1245), .A2(new_n1255), .A3(new_n1276), .A4(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G375), .A2(G378), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1279), .A2(new_n1255), .A3(new_n1261), .A4(new_n1277), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1275), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1278), .A2(new_n1281), .A3(new_n1271), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT126), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1278), .A2(new_n1281), .A3(new_n1271), .A4(KEYINPUT126), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1236), .A2(new_n1238), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1272), .B1(new_n1284), .B2(new_n1287), .ZN(G405));
  NAND2_X1  g1088(.A1(new_n1279), .A2(new_n1226), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT127), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1279), .A2(KEYINPUT127), .A3(new_n1226), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1254), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1291), .A2(new_n1254), .A3(new_n1292), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1294), .A2(new_n1239), .A3(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1295), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1286), .B1(new_n1297), .B2(new_n1293), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1296), .A2(new_n1298), .ZN(G402));
endmodule


