//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 1 1 0 1 0 1 0 1 0 1 1 1 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n732, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G210), .B1(G237), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G224), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G953), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n192), .B(KEYINPUT85), .ZN(new_n193));
  INV_X1    g007(.A(G128), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(KEYINPUT1), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G146), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G143), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n195), .A2(new_n197), .A3(new_n199), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n198), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n202), .B1(new_n196), .B2(G146), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n198), .A2(KEYINPUT64), .A3(G143), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n201), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n194), .B1(new_n199), .B2(KEYINPUT1), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n200), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  OR2_X1    g021(.A1(new_n207), .A2(G125), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  AND2_X1   g023(.A1(KEYINPUT0), .A2(G128), .ZN(new_n210));
  AND3_X1   g024(.A1(new_n197), .A2(new_n199), .A3(new_n210), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n198), .A2(KEYINPUT64), .A3(G143), .ZN(new_n212));
  AOI21_X1  g026(.A(KEYINPUT64), .B1(new_n198), .B2(G143), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n197), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(KEYINPUT0), .A2(G128), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n210), .A2(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n211), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G125), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT83), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n197), .A2(new_n199), .A3(new_n210), .ZN(new_n220));
  OR2_X1    g034(.A1(new_n210), .A2(new_n215), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n220), .B1(new_n205), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT83), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n223), .A3(G125), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n209), .B1(new_n225), .B2(KEYINPUT84), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT84), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n219), .A2(new_n227), .A3(new_n224), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n193), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n222), .A2(new_n223), .A3(G125), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n223), .B1(new_n222), .B2(G125), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT84), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  AND4_X1   g046(.A1(new_n193), .A2(new_n232), .A3(new_n228), .A4(new_n208), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(G110), .B(G122), .ZN(new_n235));
  AND2_X1   g049(.A1(KEYINPUT66), .A2(G119), .ZN(new_n236));
  NOR2_X1   g050(.A1(KEYINPUT66), .A2(G119), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT5), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(new_n239), .A3(G116), .ZN(new_n240));
  INV_X1    g054(.A(G116), .ZN(new_n241));
  OR2_X1    g055(.A1(KEYINPUT66), .A2(G119), .ZN(new_n242));
  NAND2_X1  g056(.A1(KEYINPUT66), .A2(G119), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(G116), .A2(G119), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OAI211_X1 g060(.A(G113), .B(new_n240), .C1(new_n246), .C2(new_n239), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT2), .B(G113), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n249), .B1(new_n244), .B2(new_n245), .ZN(new_n250));
  INV_X1    g064(.A(G107), .ZN(new_n251));
  AND2_X1   g065(.A1(KEYINPUT77), .A2(G104), .ZN(new_n252));
  NOR2_X1   g066(.A1(KEYINPUT77), .A2(G104), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G104), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G107), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G101), .ZN(new_n258));
  NOR3_X1   g072(.A1(new_n255), .A2(KEYINPUT3), .A3(G107), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n252), .A2(new_n253), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n259), .B1(new_n260), .B2(G107), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n262));
  INV_X1    g076(.A(G101), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n247), .A2(new_n250), .A3(new_n258), .A4(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n263), .B1(new_n261), .B2(new_n262), .ZN(new_n266));
  XOR2_X1   g080(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n267));
  AOI21_X1  g081(.A(KEYINPUT79), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT77), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n255), .ZN(new_n270));
  NAND2_X1  g084(.A1(KEYINPUT77), .A2(G104), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(G107), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT3), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(new_n251), .A3(G104), .ZN(new_n274));
  AOI21_X1  g088(.A(G107), .B1(new_n270), .B2(new_n271), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n272), .B(new_n274), .C1(new_n275), .C2(new_n273), .ZN(new_n276));
  AND4_X1   g090(.A1(KEYINPUT79), .A2(new_n276), .A3(G101), .A4(new_n267), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n268), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n246), .A2(KEYINPUT67), .A3(new_n248), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT67), .ZN(new_n280));
  OAI21_X1  g094(.A(G116), .B1(new_n236), .B2(new_n237), .ZN(new_n281));
  INV_X1    g095(.A(new_n245), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n248), .A3(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n250), .A2(new_n280), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n264), .A2(KEYINPUT4), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n279), .B(new_n284), .C1(new_n285), .C2(new_n266), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n235), .B(new_n265), .C1(new_n278), .C2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(KEYINPUT82), .A2(KEYINPUT6), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n284), .A2(new_n279), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n276), .A2(G101), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n292), .A2(KEYINPUT4), .A3(new_n264), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n291), .B(new_n293), .C1(new_n277), .C2(new_n268), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n265), .ZN(new_n295));
  INV_X1    g109(.A(new_n235), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n290), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n295), .A2(new_n296), .A3(new_n289), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n234), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G902), .ZN(new_n301));
  AND4_X1   g115(.A1(KEYINPUT7), .A2(new_n226), .A3(new_n193), .A4(new_n228), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n240), .A2(G113), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n239), .B1(new_n281), .B2(new_n282), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n250), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n264), .A2(new_n258), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n265), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT86), .B(KEYINPUT8), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n235), .B(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n219), .A2(new_n208), .A3(new_n224), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT87), .ZN(new_n312));
  OR2_X1    g126(.A1(new_n312), .A2(KEYINPUT7), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(KEYINPUT7), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n193), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  AOI22_X1  g129(.A1(new_n308), .A2(new_n310), .B1(new_n311), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n287), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n301), .B1(new_n302), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n190), .B1(new_n300), .B2(new_n318), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n287), .A2(new_n316), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n233), .A2(KEYINPUT7), .ZN(new_n321));
  AOI21_X1  g135(.A(G902), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  AOI211_X1 g136(.A(new_n235), .B(new_n288), .C1(new_n294), .C2(new_n265), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n323), .B1(new_n297), .B2(new_n290), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n322), .B(new_n189), .C1(new_n324), .C2(new_n234), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n188), .B1(new_n319), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G237), .ZN(new_n327));
  INV_X1    g141(.A(G953), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(new_n328), .A3(G214), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n196), .ZN(new_n330));
  NOR2_X1   g144(.A1(G237), .A2(G953), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(G143), .A3(G214), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G131), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT17), .ZN(new_n335));
  INV_X1    g149(.A(G131), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n330), .A2(new_n336), .A3(new_n332), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n334), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G140), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G125), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n218), .A2(G140), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT16), .ZN(new_n342));
  OR3_X1    g156(.A1(new_n218), .A2(KEYINPUT16), .A3(G140), .ZN(new_n343));
  AOI21_X1  g157(.A(G146), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n342), .A2(new_n343), .A3(G146), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n344), .B1(KEYINPUT74), .B2(new_n345), .ZN(new_n346));
  NOR3_X1   g160(.A1(new_n218), .A2(KEYINPUT16), .A3(G140), .ZN(new_n347));
  XNOR2_X1  g161(.A(G125), .B(G140), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n347), .B1(new_n348), .B2(KEYINPUT16), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT74), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n350), .A3(G146), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n333), .A2(KEYINPUT17), .A3(G131), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n338), .A2(new_n346), .A3(new_n351), .A4(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(G113), .B(G122), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n354), .B(KEYINPUT90), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(new_n255), .ZN(new_n356));
  NAND2_X1  g170(.A1(KEYINPUT18), .A2(G131), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n332), .ZN(new_n359));
  AOI21_X1  g173(.A(G143), .B1(new_n331), .B2(G214), .ZN(new_n360));
  NOR3_X1   g174(.A1(new_n359), .A2(new_n360), .A3(KEYINPUT88), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT88), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n362), .B1(new_n330), .B2(new_n332), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n358), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n330), .A2(new_n357), .A3(new_n332), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT89), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT89), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n330), .A2(new_n367), .A3(new_n357), .A4(new_n332), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n340), .A2(new_n341), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT75), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n348), .A2(KEYINPUT75), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n373), .A3(new_n198), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n370), .A2(G146), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n364), .A2(new_n369), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n353), .A2(new_n356), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n356), .B1(new_n353), .B2(new_n377), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n301), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G475), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT88), .B1(new_n359), .B2(new_n360), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n330), .A2(new_n362), .A3(new_n332), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n385), .A2(new_n358), .B1(new_n374), .B2(new_n375), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT19), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n372), .A2(new_n373), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n370), .A2(KEYINPUT19), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n198), .A3(new_n389), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n334), .A2(new_n337), .B1(G146), .B2(new_n349), .ZN(new_n391));
  AOI22_X1  g205(.A1(new_n386), .A2(new_n369), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n378), .B1(new_n392), .B2(new_n356), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT20), .ZN(new_n394));
  NOR2_X1   g208(.A1(G475), .A2(G902), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n394), .B1(new_n393), .B2(new_n395), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n382), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n196), .A2(KEYINPUT13), .A3(G128), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT91), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT91), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n402), .A2(new_n196), .A3(KEYINPUT13), .A4(G128), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n194), .A2(G143), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT13), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n405), .B1(new_n194), .B2(G143), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n401), .A2(new_n403), .A3(new_n404), .A4(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G134), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n241), .A2(G122), .ZN(new_n409));
  INV_X1    g223(.A(G122), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n410), .A2(G116), .ZN(new_n411));
  OAI21_X1  g225(.A(G107), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(G116), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n241), .A2(G122), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n414), .A3(new_n251), .ZN(new_n415));
  INV_X1    g229(.A(G134), .ZN(new_n416));
  XNOR2_X1  g230(.A(G128), .B(G143), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n412), .A2(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n408), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT92), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n408), .A2(new_n418), .A3(KEYINPUT92), .ZN(new_n422));
  XNOR2_X1  g236(.A(G116), .B(G122), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT14), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n251), .B1(new_n411), .B2(KEYINPUT14), .ZN(new_n426));
  AOI22_X1  g240(.A1(new_n425), .A2(new_n426), .B1(new_n251), .B2(new_n423), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n417), .B(new_n416), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n421), .A2(new_n422), .A3(new_n429), .ZN(new_n430));
  XOR2_X1   g244(.A(KEYINPUT70), .B(G217), .Z(new_n431));
  XOR2_X1   g245(.A(KEYINPUT9), .B(G234), .Z(new_n432));
  AND3_X1   g246(.A1(new_n431), .A2(new_n432), .A3(new_n328), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  AOI22_X1  g249(.A1(new_n419), .A2(new_n420), .B1(new_n428), .B2(new_n427), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(new_n422), .A3(new_n433), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n301), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT15), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(G478), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n439), .B(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n399), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n328), .A2(G952), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n444), .B1(G234), .B2(G237), .ZN(new_n445));
  AOI211_X1 g259(.A(new_n301), .B(new_n328), .C1(G234), .C2(G237), .ZN(new_n446));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(G898), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n443), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G221), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n450), .B1(new_n432), .B2(new_n301), .ZN(new_n451));
  INV_X1    g265(.A(G469), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(new_n301), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n217), .B(new_n293), .C1(new_n268), .C2(new_n277), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n263), .B1(new_n254), .B2(new_n256), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n270), .A2(new_n271), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n273), .B1(new_n456), .B2(new_n251), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n272), .A2(new_n274), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n455), .B1(new_n459), .B2(new_n263), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n207), .A2(KEYINPUT10), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n197), .A2(new_n199), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n200), .B1(new_n462), .B2(new_n206), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n258), .B(new_n463), .C1(new_n276), .C2(G101), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT10), .ZN(new_n465));
  AOI22_X1  g279(.A1(new_n460), .A2(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n454), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT11), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n468), .B1(new_n416), .B2(G137), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n416), .A2(G137), .ZN(new_n470));
  INV_X1    g284(.A(G137), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(KEYINPUT11), .A3(G134), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n469), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G131), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n469), .A2(new_n472), .A3(new_n336), .A4(new_n470), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n467), .A2(new_n476), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n474), .A2(new_n475), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n478), .B(KEYINPUT80), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n293), .A2(new_n217), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n466), .B(new_n479), .C1(new_n278), .C2(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(G110), .B(G140), .ZN(new_n482));
  INV_X1    g296(.A(G227), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n483), .A2(G953), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n482), .B(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(KEYINPUT12), .B1(new_n476), .B2(KEYINPUT81), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n264), .A2(new_n258), .A3(new_n463), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n207), .B1(new_n264), .B2(new_n258), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n489), .B(new_n476), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n464), .B1(new_n460), .B2(new_n207), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n489), .B1(new_n494), .B2(new_n476), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n481), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n477), .A2(new_n487), .B1(new_n496), .B2(new_n485), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n453), .B1(new_n497), .B2(G469), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n454), .A2(new_n466), .A3(new_n479), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n478), .B1(new_n454), .B2(new_n466), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n485), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n476), .B1(new_n490), .B2(new_n491), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n488), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n492), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n504), .A2(new_n481), .A3(new_n486), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(new_n452), .A3(new_n301), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n451), .B1(new_n498), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n326), .A2(new_n449), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT93), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n328), .A2(G221), .A3(G234), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(KEYINPUT22), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(G137), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(G110), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT66), .B(G119), .ZN(new_n517));
  OAI21_X1  g331(.A(KEYINPUT23), .B1(new_n517), .B2(new_n194), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT72), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g334(.A(KEYINPUT72), .B(KEYINPUT23), .C1(new_n517), .C2(new_n194), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT73), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n522), .B1(new_n238), .B2(G128), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n517), .A2(KEYINPUT73), .A3(new_n194), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n520), .A2(new_n521), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n194), .A2(G119), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT23), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n516), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n345), .A2(KEYINPUT74), .ZN(new_n529));
  INV_X1    g343(.A(new_n344), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n351), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n526), .B1(new_n238), .B2(G128), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT24), .B(G110), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n528), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n374), .A2(new_n345), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n521), .A2(new_n523), .A3(new_n524), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n238), .A2(G128), .ZN(new_n540));
  AOI21_X1  g354(.A(KEYINPUT72), .B1(new_n540), .B2(KEYINPUT23), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n516), .B(new_n527), .C1(new_n539), .C2(new_n541), .ZN(new_n542));
  OR2_X1    g356(.A1(new_n532), .A2(new_n534), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n538), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n515), .B1(new_n537), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n542), .A2(new_n543), .ZN(new_n546));
  INV_X1    g360(.A(new_n538), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n527), .B1(new_n539), .B2(new_n541), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(G110), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n346), .A2(new_n351), .B1(new_n532), .B2(new_n534), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n548), .A2(new_n552), .A3(new_n514), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n545), .A2(new_n553), .A3(new_n301), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT25), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT25), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n545), .A2(new_n553), .A3(new_n556), .A4(new_n301), .ZN(new_n557));
  INV_X1    g371(.A(G234), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n431), .B1(new_n558), .B2(G902), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(KEYINPUT71), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n555), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT76), .ZN(new_n562));
  INV_X1    g376(.A(new_n560), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n563), .B1(new_n554), .B2(KEYINPUT25), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT76), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(new_n565), .A3(new_n557), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n545), .A2(new_n553), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n560), .A2(G902), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n562), .A2(new_n566), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G472), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n217), .A2(new_n476), .ZN(new_n572));
  INV_X1    g386(.A(new_n470), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n416), .A2(G137), .ZN(new_n574));
  OAI21_X1  g388(.A(G131), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n207), .A2(new_n575), .A3(new_n475), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n572), .A2(new_n576), .A3(KEYINPUT30), .ZN(new_n577));
  INV_X1    g391(.A(new_n576), .ZN(new_n578));
  OAI21_X1  g392(.A(KEYINPUT65), .B1(new_n478), .B2(new_n222), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT65), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n217), .A2(new_n476), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n578), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n291), .B(new_n577), .C1(new_n582), .C2(KEYINPUT30), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n284), .A2(new_n279), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(new_n576), .A3(new_n572), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT27), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n331), .A2(new_n587), .A3(G210), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n587), .B1(new_n331), .B2(G210), .ZN(new_n590));
  OAI21_X1  g404(.A(KEYINPUT26), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n590), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT26), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n593), .A3(new_n588), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n591), .A2(new_n594), .A3(G101), .ZN(new_n595));
  AOI21_X1  g409(.A(G101), .B1(new_n591), .B2(new_n594), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n586), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT29), .ZN(new_n600));
  OR2_X1    g414(.A1(new_n582), .A2(new_n584), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT28), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n585), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n585), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(KEYINPUT28), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n601), .A2(new_n603), .A3(new_n605), .A4(new_n597), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n599), .A2(new_n600), .A3(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n598), .A2(new_n600), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n572), .A2(new_n576), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n291), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n605), .A2(new_n608), .A3(new_n603), .A4(new_n610), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n611), .A2(new_n301), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n571), .B1(new_n607), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(G472), .A2(G902), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT69), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT68), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n585), .B2(new_n597), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n585), .A2(new_n617), .A3(new_n597), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n583), .B(new_n616), .C1(new_n618), .C2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT31), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n618), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n619), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n625), .A2(new_n616), .A3(KEYINPUT31), .A4(new_n583), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n605), .A2(new_n603), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n601), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n598), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n615), .B1(new_n627), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n613), .B1(new_n631), .B2(KEYINPUT32), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT32), .ZN(new_n633));
  AOI22_X1  g447(.A1(new_n623), .A2(new_n626), .B1(new_n629), .B2(new_n598), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n633), .B1(new_n634), .B2(new_n615), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n570), .B1(new_n632), .B2(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n449), .A2(new_n326), .A3(new_n508), .A4(KEYINPUT93), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n511), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT94), .B(G101), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G3));
  NAND2_X1  g454(.A1(new_n301), .A2(G478), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT95), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n436), .A2(new_n422), .A3(new_n433), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n433), .B1(new_n436), .B2(new_n422), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n430), .A2(KEYINPUT33), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT33), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n646), .A2(new_n647), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n438), .A2(new_n650), .A3(new_n642), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n641), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(G478), .B1(new_n438), .B2(new_n301), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n399), .ZN(new_n655));
  INV_X1    g469(.A(new_n448), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n326), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n631), .ZN(new_n658));
  OAI21_X1  g472(.A(G472), .B1(new_n634), .B2(G902), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n451), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n477), .A2(new_n481), .A3(new_n486), .ZN(new_n663));
  AND2_X1   g477(.A1(new_n504), .A2(new_n481), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n663), .B(G469), .C1(new_n664), .C2(new_n486), .ZN(new_n665));
  INV_X1    g479(.A(new_n453), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI211_X1 g481(.A(G469), .B(G902), .C1(new_n501), .C2(new_n505), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n662), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n570), .A2(new_n669), .ZN(new_n670));
  AND4_X1   g484(.A1(new_n655), .A2(new_n657), .A3(new_n661), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT34), .B(G104), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT96), .B(KEYINPUT97), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G6));
  NOR2_X1   g489(.A1(new_n442), .A2(new_n398), .ZN(new_n676));
  AND3_X1   g490(.A1(new_n326), .A2(new_n656), .A3(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n677), .A2(new_n661), .A3(new_n670), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT35), .B(G107), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G9));
  AND3_X1   g494(.A1(new_n564), .A2(new_n565), .A3(new_n557), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n565), .B1(new_n564), .B2(new_n557), .ZN(new_n682));
  OAI22_X1  g496(.A1(new_n537), .A2(new_n544), .B1(KEYINPUT36), .B2(new_n515), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n515), .A2(KEYINPUT36), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n548), .A2(new_n552), .A3(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n683), .A2(new_n568), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT98), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n681), .A2(new_n682), .A3(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n660), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n511), .A2(new_n637), .A3(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT37), .B(G110), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G12));
  INV_X1    g507(.A(G900), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n445), .B1(new_n446), .B2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n676), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n697), .B1(new_n632), .B2(new_n635), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n686), .B(KEYINPUT98), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n562), .A2(new_n699), .A3(new_n566), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n326), .A2(new_n508), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G128), .ZN(G30));
  XOR2_X1   g517(.A(new_n695), .B(KEYINPUT39), .Z(new_n704));
  NAND2_X1  g518(.A1(new_n508), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT40), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n319), .A2(new_n325), .ZN(new_n707));
  XOR2_X1   g521(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT100), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n707), .B(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n399), .A2(new_n442), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n689), .A2(new_n187), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n631), .A2(KEYINPUT32), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n625), .A2(new_n583), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n597), .B1(new_n610), .B2(new_n585), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n301), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(G472), .ZN(new_n717));
  AND3_X1   g531(.A1(new_n713), .A2(new_n717), .A3(new_n635), .ZN(new_n718));
  NOR4_X1   g532(.A1(new_n706), .A2(new_n710), .A3(new_n712), .A4(new_n718), .ZN(new_n719));
  XOR2_X1   g533(.A(new_n719), .B(KEYINPUT101), .Z(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(new_n196), .ZN(G45));
  OAI211_X1 g535(.A(new_n398), .B(new_n696), .C1(new_n652), .C2(new_n653), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n632), .B2(new_n635), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n701), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(KEYINPUT102), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(new_n198), .ZN(G48));
  AOI21_X1  g540(.A(new_n452), .B1(new_n506), .B2(new_n301), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n727), .A2(new_n668), .A3(new_n451), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n636), .A2(new_n655), .A3(new_n657), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT41), .B(G113), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G15));
  NAND3_X1  g545(.A1(new_n636), .A2(new_n677), .A3(new_n728), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G116), .ZN(G18));
  AND3_X1   g547(.A1(new_n728), .A2(new_n326), .A3(new_n700), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n632), .A2(new_n635), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n734), .A2(new_n735), .A3(new_n449), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G119), .ZN(G21));
  AND3_X1   g551(.A1(new_n707), .A2(new_n187), .A3(new_n711), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n628), .A2(new_n610), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n598), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n627), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n614), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n659), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n570), .ZN(new_n744));
  NOR4_X1   g558(.A1(new_n727), .A2(new_n668), .A3(new_n448), .A4(new_n451), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n738), .A2(new_n743), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G122), .ZN(G24));
  AND2_X1   g561(.A1(new_n728), .A2(new_n326), .ZN(new_n748));
  INV_X1    g562(.A(new_n722), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n659), .A2(new_n742), .A3(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n748), .A2(new_n700), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G125), .ZN(G27));
  NOR3_X1   g566(.A1(new_n669), .A2(new_n707), .A3(new_n188), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n636), .A2(new_n749), .A3(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT42), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n635), .A2(KEYINPUT103), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n635), .A2(KEYINPUT103), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(new_n632), .A3(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n722), .A2(new_n755), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n759), .A2(new_n744), .A3(new_n753), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n756), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT104), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT104), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n756), .A2(new_n761), .A3(new_n764), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G131), .ZN(G33));
  NAND4_X1  g581(.A1(new_n636), .A2(new_n676), .A3(new_n696), .A4(new_n753), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G134), .ZN(G36));
  OAI21_X1  g583(.A(new_n663), .B1(new_n664), .B2(new_n486), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT45), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n497), .A2(KEYINPUT45), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n773), .A3(G469), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n666), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT46), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT105), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n774), .A2(KEYINPUT46), .A3(new_n666), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n779), .A2(new_n507), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT46), .B1(new_n774), .B2(new_n666), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT105), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n778), .A2(new_n780), .A3(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(new_n662), .A3(new_n704), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n707), .A2(new_n188), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n660), .A2(new_n700), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT106), .ZN(new_n788));
  OR3_X1    g602(.A1(new_n654), .A2(KEYINPUT43), .A3(new_n398), .ZN(new_n789));
  OAI21_X1  g603(.A(KEYINPUT43), .B1(new_n654), .B2(new_n398), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(KEYINPUT44), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n793), .A2(KEYINPUT107), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(KEYINPUT107), .ZN(new_n795));
  OAI221_X1 g609(.A(new_n786), .B1(KEYINPUT44), .B2(new_n792), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT108), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n785), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n798), .B1(new_n797), .B2(new_n796), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G137), .ZN(G39));
  OAI211_X1 g614(.A(new_n507), .B(new_n779), .C1(new_n781), .C2(new_n782), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n777), .A2(KEYINPUT105), .ZN(new_n802));
  OAI211_X1 g616(.A(KEYINPUT109), .B(new_n662), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT109), .B1(new_n784), .B2(new_n662), .ZN(new_n805));
  XOR2_X1   g619(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n806));
  NOR3_X1   g620(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n662), .B1(new_n801), .B2(new_n802), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT109), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n808), .B1(new_n811), .B2(new_n803), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n786), .A2(new_n570), .A3(new_n749), .ZN(new_n813));
  OR4_X1    g627(.A1(new_n735), .A2(new_n807), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G140), .ZN(G42));
  OR2_X1    g629(.A1(G952), .A2(G953), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n727), .A2(new_n668), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  OAI22_X1  g632(.A1(new_n807), .A2(new_n812), .B1(new_n662), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n743), .A2(new_n744), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n789), .A2(new_n445), .A3(new_n790), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(new_n786), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n819), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n710), .A2(new_n188), .A3(new_n728), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n822), .A2(new_n827), .ZN(new_n828));
  XOR2_X1   g642(.A(new_n828), .B(KEYINPUT50), .Z(new_n829));
  AND2_X1   g643(.A1(new_n786), .A2(new_n728), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n830), .A2(new_n821), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n831), .A2(new_n700), .A3(new_n743), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT118), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n830), .A2(new_n744), .A3(new_n445), .A4(new_n718), .ZN(new_n834));
  NOR4_X1   g648(.A1(new_n834), .A2(new_n398), .A3(new_n653), .A4(new_n652), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n829), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n836), .A2(KEYINPUT51), .ZN(new_n837));
  XOR2_X1   g651(.A(new_n444), .B(KEYINPUT120), .Z(new_n838));
  INV_X1    g652(.A(new_n655), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n834), .A2(new_n839), .ZN(new_n840));
  AOI211_X1 g654(.A(new_n838), .B(new_n840), .C1(new_n748), .C2(new_n823), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n759), .A2(new_n744), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n831), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT48), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n845), .A2(KEYINPUT121), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(KEYINPUT121), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n826), .A2(new_n837), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n819), .A2(new_n849), .A3(new_n825), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n818), .A2(new_n662), .ZN(new_n851));
  OAI22_X1  g665(.A1(new_n804), .A2(new_n805), .B1(KEYINPUT110), .B2(KEYINPUT47), .ZN(new_n852));
  INV_X1    g666(.A(new_n806), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n811), .A2(new_n803), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n851), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT117), .B1(new_n855), .B2(new_n824), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n850), .A2(new_n856), .A3(new_n836), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT51), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n857), .A2(KEYINPUT119), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT119), .B1(new_n857), .B2(new_n858), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n848), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT122), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n848), .B(KEYINPUT122), .C1(new_n859), .C2(new_n860), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n689), .A2(KEYINPUT112), .A3(new_n508), .A4(new_n696), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT112), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n662), .B(new_n696), .C1(new_n667), .C2(new_n668), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n868), .B1(new_n869), .B2(new_n700), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n713), .A2(new_n717), .A3(new_n635), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n867), .A2(new_n870), .A3(new_n871), .A4(new_n738), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n872), .A2(new_n702), .A3(new_n724), .A4(new_n751), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT52), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI22_X1  g689(.A1(new_n701), .A2(new_n698), .B1(new_n734), .B2(new_n750), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n876), .A2(KEYINPUT52), .A3(new_n724), .A4(new_n872), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  OR2_X1    g692(.A1(new_n655), .A2(new_n676), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n657), .A2(new_n661), .A3(new_n670), .A4(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n638), .A2(new_n691), .A3(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n729), .A2(new_n732), .A3(new_n736), .A4(new_n746), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n443), .A2(new_n695), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n750), .B1(new_n735), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n753), .A2(new_n700), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n768), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n881), .A2(new_n882), .A3(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n766), .A2(new_n866), .A3(new_n878), .A4(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n881), .A2(new_n882), .ZN(new_n889));
  INV_X1    g703(.A(new_n886), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n889), .A2(new_n763), .A3(new_n765), .A4(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n875), .A2(KEYINPUT113), .A3(new_n877), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT113), .B1(new_n875), .B2(new_n877), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n888), .B1(new_n894), .B2(new_n866), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT54), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n881), .A2(new_n886), .A3(new_n866), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n878), .ZN(new_n899));
  INV_X1    g713(.A(new_n882), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n762), .ZN(new_n901));
  OR2_X1    g715(.A1(new_n901), .A2(KEYINPUT115), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(KEYINPUT115), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n899), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT114), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n905), .B1(new_n894), .B2(KEYINPUT53), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT113), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n878), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n875), .A2(KEYINPUT113), .A3(new_n877), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n766), .A2(new_n908), .A3(new_n909), .A4(new_n887), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n910), .A2(KEYINPUT114), .A3(new_n866), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n904), .B1(new_n906), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n896), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n897), .B1(new_n913), .B2(KEYINPUT116), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n914), .B1(KEYINPUT116), .B2(new_n913), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n816), .B1(new_n865), .B2(new_n915), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n570), .A2(new_n188), .A3(new_n451), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT111), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT49), .ZN(new_n919));
  OAI221_X1 g733(.A(new_n399), .B1(new_n653), .B2(new_n652), .C1(new_n817), .C2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n920), .B1(new_n919), .B2(new_n817), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n918), .A2(new_n710), .A3(new_n718), .A4(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n916), .A2(new_n922), .ZN(G75));
  NOR2_X1   g737(.A1(new_n912), .A2(new_n301), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(G210), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n324), .B(new_n234), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT55), .Z(new_n927));
  INV_X1    g741(.A(KEYINPUT123), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n928), .A2(KEYINPUT56), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n925), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n927), .B1(new_n925), .B2(new_n929), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n328), .A2(G952), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(G51));
  NOR3_X1   g747(.A1(new_n912), .A2(new_n301), .A3(new_n774), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n453), .B(KEYINPUT124), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT57), .Z(new_n936));
  NAND2_X1  g750(.A1(new_n906), .A2(new_n911), .ZN(new_n937));
  INV_X1    g751(.A(new_n904), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n896), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AOI211_X1 g753(.A(KEYINPUT54), .B(new_n904), .C1(new_n906), .C2(new_n911), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n936), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n506), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT125), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n934), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n941), .A2(KEYINPUT125), .A3(new_n506), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n932), .B1(new_n944), .B2(new_n945), .ZN(G54));
  NAND3_X1  g760(.A1(new_n924), .A2(KEYINPUT58), .A3(G475), .ZN(new_n947));
  INV_X1    g761(.A(new_n393), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n947), .A2(new_n948), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n949), .A2(new_n950), .A3(new_n932), .ZN(G60));
  NAND2_X1  g765(.A1(new_n649), .A2(new_n651), .ZN(new_n952));
  NAND2_X1  g766(.A1(G478), .A2(G902), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT59), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n952), .B1(new_n915), .B2(new_n954), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n952), .B(new_n954), .C1(new_n939), .C2(new_n940), .ZN(new_n956));
  INV_X1    g770(.A(new_n932), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n955), .A2(new_n958), .ZN(G63));
  INV_X1    g773(.A(KEYINPUT126), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(KEYINPUT61), .ZN(new_n961));
  INV_X1    g775(.A(new_n912), .ZN(new_n962));
  NAND2_X1  g776(.A1(G217), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT60), .Z(new_n964));
  NAND4_X1  g778(.A1(new_n962), .A2(new_n685), .A3(new_n683), .A4(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n957), .B1(new_n960), .B2(KEYINPUT61), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n962), .A2(new_n964), .ZN(new_n969));
  INV_X1    g783(.A(new_n567), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n961), .B1(new_n968), .B2(new_n971), .ZN(new_n972));
  AND4_X1   g786(.A1(new_n961), .A2(new_n971), .A3(new_n965), .A4(new_n967), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n972), .A2(new_n973), .ZN(G66));
  NOR3_X1   g788(.A1(new_n447), .A2(new_n191), .A3(new_n328), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n975), .B1(new_n889), .B2(new_n328), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n324), .B1(G898), .B2(new_n328), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n976), .B(new_n977), .ZN(G69));
  OAI21_X1  g792(.A(new_n577), .B1(new_n582), .B2(KEYINPUT30), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT127), .Z(new_n980));
  NAND2_X1  g794(.A1(new_n388), .A2(new_n389), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n799), .A2(new_n814), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n842), .A2(new_n738), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n984), .A2(new_n785), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n876), .A2(new_n724), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n766), .A2(new_n768), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n988), .A2(G953), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n983), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n483), .A2(new_n328), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n982), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OR2_X1    g806(.A1(new_n982), .A2(G227), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n328), .B1(new_n993), .B2(G900), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT62), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n995), .B1(new_n720), .B2(new_n986), .ZN(new_n996));
  OR3_X1    g810(.A1(new_n720), .A2(new_n995), .A3(new_n986), .ZN(new_n997));
  AND4_X1   g811(.A1(new_n508), .A2(new_n879), .A3(new_n704), .A4(new_n786), .ZN(new_n998));
  AOI22_X1  g812(.A1(new_n996), .A2(new_n997), .B1(new_n636), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n983), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n982), .A2(G953), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n994), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n992), .A2(new_n1002), .ZN(G72));
  NOR3_X1   g817(.A1(new_n988), .A2(new_n882), .A3(new_n881), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n799), .A2(new_n814), .A3(new_n987), .A4(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(G472), .A2(G902), .ZN(new_n1006));
  XOR2_X1   g820(.A(new_n1006), .B(KEYINPUT63), .Z(new_n1007));
  AOI211_X1 g821(.A(new_n597), .B(new_n586), .C1(new_n1005), .C2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n586), .A2(new_n597), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n799), .A2(new_n814), .A3(new_n889), .A4(new_n999), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1009), .B1(new_n1010), .B2(new_n1007), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n597), .B1(new_n583), .B2(new_n585), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1007), .B1(new_n714), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n957), .B1(new_n895), .B2(new_n1013), .ZN(new_n1014));
  NOR3_X1   g828(.A1(new_n1008), .A2(new_n1011), .A3(new_n1014), .ZN(G57));
endmodule


