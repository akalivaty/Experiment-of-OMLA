//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 1 0 1 0 1 0 1 0 0 0 1 1 0 1 1 1 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n811, new_n812, new_n814, new_n815,
    new_n816, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928;
  INV_X1    g000(.A(KEYINPUT3), .ZN(new_n202));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT77), .B(KEYINPUT22), .Z(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  INV_X1    g004(.A(G218gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n203), .B1(new_n204), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n202), .B1(new_n210), .B2(KEYINPUT29), .ZN(new_n211));
  XNOR2_X1  g010(.A(G155gat), .B(G162gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(G141gat), .B(G148gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT81), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n213), .B(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n212), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G155gat), .ZN(new_n218));
  INV_X1    g017(.A(G162gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n216), .A2(new_n218), .A3(new_n219), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n213), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n217), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n211), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT82), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n227), .B1(new_n224), .B2(new_n202), .ZN(new_n228));
  NOR4_X1   g027(.A1(new_n217), .A2(KEYINPUT82), .A3(KEYINPUT3), .A4(new_n223), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n230), .A2(KEYINPUT29), .ZN(new_n231));
  INV_X1    g030(.A(new_n210), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n226), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G228gat), .A2(G233gat), .ZN(new_n234));
  OR2_X1    g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n234), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(G22gat), .B1(new_n237), .B2(KEYINPUT85), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT85), .ZN(new_n239));
  INV_X1    g038(.A(G22gat), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n235), .A2(new_n239), .A3(new_n240), .A4(new_n236), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n237), .A2(KEYINPUT85), .ZN(new_n243));
  XNOR2_X1  g042(.A(G50gat), .B(G78gat), .ZN(new_n244));
  INV_X1    g043(.A(G106gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(KEYINPUT84), .B(KEYINPUT31), .Z(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n243), .A2(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(new_n242), .B(new_n249), .Z(new_n250));
  INV_X1    g049(.A(KEYINPUT73), .ZN(new_n251));
  OAI21_X1  g050(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NOR3_X1   g052(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT23), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT65), .ZN(new_n256));
  NOR2_X1   g055(.A1(G169gat), .A2(G176gat), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n256), .B1(new_n257), .B2(KEYINPUT23), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT23), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n259), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G169gat), .A2(G176gat), .ZN(new_n262));
  AND4_X1   g061(.A1(KEYINPUT25), .A2(new_n255), .A3(new_n261), .A4(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT67), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(G183gat), .ZN(new_n270));
  INV_X1    g069(.A(G190gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g071(.A1(KEYINPUT68), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n269), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n275));
  AND3_X1   g074(.A1(new_n266), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n275), .B1(new_n266), .B2(new_n274), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n263), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT70), .ZN(new_n279));
  INV_X1    g078(.A(new_n264), .ZN(new_n280));
  AOI22_X1  g079(.A1(new_n280), .A2(KEYINPUT64), .B1(new_n270), .B2(new_n271), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n281), .B(new_n267), .C1(KEYINPUT64), .C2(new_n280), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n257), .A2(KEYINPUT23), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n282), .A2(new_n262), .A3(new_n283), .A4(new_n261), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT25), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n287), .B(new_n263), .C1(new_n276), .C2(new_n277), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n279), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G120gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G113gat), .ZN(new_n291));
  INV_X1    g090(.A(G113gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G120gat), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT1), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G127gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(KEYINPUT72), .A2(G127gat), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n296), .B1(new_n294), .B2(new_n297), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n298), .A2(G134gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n298), .A2(G134gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n253), .A2(new_n254), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n302), .B(new_n262), .C1(new_n303), .C2(KEYINPUT26), .ZN(new_n304));
  NAND2_X1  g103(.A1(G183gat), .A2(G190gat), .ZN(new_n305));
  XOR2_X1   g104(.A(KEYINPUT27), .B(G183gat), .Z(new_n306));
  OAI21_X1  g105(.A(KEYINPUT28), .B1(new_n306), .B2(G190gat), .ZN(new_n307));
  OR3_X1    g106(.A1(new_n270), .A2(KEYINPUT71), .A3(KEYINPUT27), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT28), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT27), .B1(new_n270), .B2(KEYINPUT71), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n308), .A2(new_n309), .A3(new_n271), .A4(new_n310), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n304), .A2(new_n305), .A3(new_n307), .A4(new_n311), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n289), .A2(new_n301), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n301), .B1(new_n289), .B2(new_n312), .ZN(new_n314));
  NAND2_X1  g113(.A1(G227gat), .A2(G233gat), .ZN(new_n315));
  NOR3_X1   g114(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n251), .B1(new_n316), .B2(KEYINPUT33), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n289), .A2(new_n312), .ZN(new_n318));
  OR2_X1    g117(.A1(new_n299), .A2(new_n300), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n289), .A2(new_n301), .A3(new_n312), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n320), .A2(G227gat), .A3(G233gat), .A4(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT33), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n322), .A2(KEYINPUT73), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(KEYINPUT32), .ZN(new_n325));
  XNOR2_X1  g124(.A(G15gat), .B(G43gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(G71gat), .ZN(new_n327));
  INV_X1    g126(.A(G99gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n327), .B(new_n328), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n317), .A2(new_n324), .A3(new_n325), .A4(new_n329), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n320), .A2(new_n321), .B1(G227gat), .B2(G233gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n331), .B(KEYINPUT34), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n329), .A2(KEYINPUT33), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n322), .A2(KEYINPUT32), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT74), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n322), .A2(new_n336), .A3(KEYINPUT32), .A4(new_n333), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n330), .A2(new_n332), .A3(new_n335), .A4(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT75), .ZN(new_n339));
  AND2_X1   g138(.A1(new_n335), .A2(new_n337), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n340), .A2(new_n341), .A3(new_n332), .A4(new_n330), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n340), .A2(new_n330), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n344), .A2(new_n332), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n250), .A2(new_n346), .ZN(new_n347));
  AND3_X1   g146(.A1(new_n318), .A2(G226gat), .A3(G233gat), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT29), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n318), .A2(new_n349), .B1(G226gat), .B2(G233gat), .ZN(new_n350));
  OR3_X1    g149(.A1(new_n348), .A2(new_n350), .A3(new_n210), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n210), .B1(new_n348), .B2(new_n350), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G8gat), .B(G36gat), .ZN(new_n354));
  INV_X1    g153(.A(G64gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n354), .B(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(G92gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT78), .B1(new_n353), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n360));
  INV_X1    g159(.A(new_n358), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n351), .A2(new_n360), .A3(new_n361), .A4(new_n352), .ZN(new_n362));
  XOR2_X1   g161(.A(KEYINPUT79), .B(KEYINPUT30), .Z(new_n363));
  NAND3_X1  g162(.A1(new_n359), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT80), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n361), .B1(new_n351), .B2(new_n352), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n353), .A2(new_n358), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n366), .B1(new_n367), .B2(KEYINPUT30), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n359), .A2(new_n369), .A3(new_n362), .A4(new_n363), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n365), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(KEYINPUT0), .B(G57gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n373), .B(G85gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(G1gat), .B(G29gat), .ZN(new_n375));
  XOR2_X1   g174(.A(new_n374), .B(new_n375), .Z(new_n376));
  NAND2_X1  g175(.A1(new_n319), .A2(new_n224), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT4), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT4), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n319), .A2(new_n379), .A3(new_n224), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  OAI221_X1 g180(.A(new_n301), .B1(new_n202), .B2(new_n224), .C1(new_n228), .C2(new_n229), .ZN(new_n382));
  NAND2_X1  g181(.A1(G225gat), .A2(G233gat), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n377), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n381), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  NOR3_X1   g185(.A1(new_n319), .A2(KEYINPUT83), .A3(new_n224), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT83), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n388), .B1(new_n225), .B2(new_n301), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n377), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n384), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n386), .A2(new_n391), .A3(KEYINPUT5), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n381), .A2(new_n382), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n384), .A2(KEYINPUT5), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n376), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT6), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n392), .A2(new_n395), .A3(new_n376), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n396), .A2(KEYINPUT6), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n372), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT35), .B1(new_n347), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT76), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n339), .A2(new_n405), .A3(new_n342), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n405), .B1(new_n339), .B2(new_n342), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n345), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n371), .A2(KEYINPUT35), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT88), .ZN(new_n412));
  AND3_X1   g211(.A1(new_n396), .A2(new_n412), .A3(KEYINPUT6), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n412), .B1(new_n396), .B2(KEYINPUT6), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT86), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT86), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n397), .A2(new_n417), .A3(new_n398), .A4(new_n399), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n415), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n410), .A2(new_n250), .A3(new_n411), .A4(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n421), .ZN(new_n422));
  OR2_X1    g221(.A1(new_n393), .A2(new_n383), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n423), .B(KEYINPUT39), .C1(new_n384), .C2(new_n390), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n424), .B(new_n376), .C1(KEYINPUT39), .C2(new_n423), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT40), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n396), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n371), .B(new_n427), .C1(new_n426), .C2(new_n425), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n359), .A2(new_n362), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n353), .A2(KEYINPUT37), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT37), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n351), .A2(new_n431), .A3(new_n352), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n430), .A2(new_n358), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n429), .B1(KEYINPUT38), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT87), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n435), .B1(new_n433), .B2(KEYINPUT38), .ZN(new_n436));
  OR3_X1    g235(.A1(new_n433), .A2(new_n435), .A3(KEYINPUT38), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n419), .A2(new_n434), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n428), .A2(new_n438), .A3(new_n250), .ZN(new_n439));
  INV_X1    g238(.A(new_n345), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT36), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n440), .B(new_n441), .C1(new_n406), .C2(new_n408), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT36), .B1(new_n343), .B2(new_n345), .ZN(new_n443));
  AND2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n250), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n403), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n439), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n422), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT17), .ZN(new_n449));
  INV_X1    g248(.A(G50gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(G43gat), .ZN(new_n451));
  INV_X1    g250(.A(G43gat), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(G50gat), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n451), .A2(new_n453), .A3(KEYINPUT15), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT15), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n452), .A2(G50gat), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n450), .A2(G43gat), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(G29gat), .A2(G36gat), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT14), .ZN(new_n460));
  INV_X1    g259(.A(G29gat), .ZN(new_n461));
  INV_X1    g260(.A(G36gat), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AND4_X1   g264(.A1(new_n454), .A2(new_n458), .A3(new_n459), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(KEYINPUT90), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT90), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n468), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n467), .A2(new_n469), .A3(new_n463), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n454), .B1(new_n470), .B2(new_n459), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT91), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n466), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n470), .A2(new_n459), .ZN(new_n474));
  INV_X1    g273(.A(new_n454), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n458), .A2(new_n454), .A3(new_n459), .A4(new_n465), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT91), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n449), .B1(new_n473), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(G15gat), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n480), .A2(new_n240), .ZN(new_n481));
  NOR2_X1   g280(.A1(G15gat), .A2(G22gat), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT92), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT16), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(new_n481), .B2(new_n482), .ZN(new_n485));
  INV_X1    g284(.A(G1gat), .ZN(new_n486));
  INV_X1    g285(.A(G8gat), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n487), .B1(new_n485), .B2(new_n486), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n483), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n490), .ZN(new_n492));
  INV_X1    g291(.A(new_n483), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n492), .A2(new_n493), .A3(new_n488), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n466), .A2(new_n471), .A3(new_n449), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n479), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(G229gat), .A2(G233gat), .ZN(new_n499));
  INV_X1    g298(.A(new_n495), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n472), .B1(new_n466), .B2(new_n471), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n476), .A2(KEYINPUT91), .A3(new_n477), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n498), .A2(KEYINPUT18), .A3(new_n499), .A4(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n499), .B(KEYINPUT13), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n500), .A2(new_n503), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n495), .B1(new_n501), .B2(new_n502), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(G113gat), .B(G141gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n512), .B(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G169gat), .B(G197gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(KEYINPUT12), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n498), .A2(new_n499), .A3(new_n504), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT18), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n511), .A2(new_n517), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT93), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n518), .A2(new_n523), .A3(new_n519), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n523), .B1(new_n518), .B2(new_n519), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n505), .A2(new_n510), .ZN(new_n526));
  NOR3_X1   g325(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT94), .B1(new_n527), .B2(new_n517), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n520), .A2(KEYINPUT93), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n518), .A2(new_n523), .A3(new_n519), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n529), .A2(new_n511), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT94), .ZN(new_n532));
  INV_X1    g331(.A(new_n517), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n522), .B1(new_n528), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT97), .ZN(new_n536));
  NAND2_X1  g335(.A1(G85gat), .A2(G92gat), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n536), .B1(new_n537), .B2(KEYINPUT98), .ZN(new_n538));
  NAND3_X1  g337(.A1(KEYINPUT97), .A2(G85gat), .A3(G92gat), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n538), .A2(KEYINPUT7), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(G85gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(new_n357), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT7), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n536), .B(new_n543), .C1(new_n537), .C2(KEYINPUT98), .ZN(new_n544));
  NAND2_X1  g343(.A1(G99gat), .A2(G106gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT8), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n540), .A2(new_n542), .A3(new_n544), .A4(new_n546), .ZN(new_n547));
  AND2_X1   g346(.A1(G99gat), .A2(G106gat), .ZN(new_n548));
  NOR2_X1   g347(.A1(G99gat), .A2(G106gat), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT99), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n328), .A2(new_n245), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT99), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(new_n552), .A3(new_n545), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n547), .A2(new_n554), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n550), .A2(new_n553), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n544), .A2(new_n546), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n556), .A2(new_n542), .A3(new_n557), .A4(new_n540), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(G57gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(G64gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n355), .A2(G57gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G71gat), .A2(G78gat), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT9), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(G71gat), .ZN(new_n567));
  INV_X1    g366(.A(G78gat), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n563), .A2(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n564), .B(KEYINPUT95), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT96), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n562), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n355), .A2(KEYINPUT96), .A3(G57gat), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n572), .A2(new_n561), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n567), .A2(new_n568), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n564), .B1(new_n575), .B2(new_n565), .ZN(new_n576));
  AOI22_X1  g375(.A1(new_n569), .A2(new_n570), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n559), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT10), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n555), .A2(new_n558), .A3(new_n577), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n559), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n583), .A2(KEYINPUT10), .A3(new_n577), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G230gat), .A2(G233gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n579), .A2(new_n581), .ZN(new_n588));
  INV_X1    g387(.A(new_n586), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(G120gat), .B(G148gat), .Z(new_n591));
  XNOR2_X1  g390(.A(G176gat), .B(G204gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n593), .B(new_n594), .Z(new_n595));
  NAND3_X1  g394(.A1(new_n587), .A2(new_n590), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT104), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n596), .A2(KEYINPUT104), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n589), .B1(new_n582), .B2(new_n584), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n600), .B1(new_n588), .B2(new_n589), .ZN(new_n601));
  OAI22_X1  g400(.A1(new_n598), .A2(new_n599), .B1(new_n601), .B2(new_n595), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n535), .A2(new_n602), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n448), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n479), .A2(new_n559), .A3(new_n497), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(KEYINPUT100), .ZN(new_n606));
  AND3_X1   g405(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n607), .B1(new_n503), .B2(new_n583), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n496), .B1(new_n503), .B2(new_n449), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT100), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n609), .A2(new_n610), .A3(new_n559), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n606), .A2(new_n608), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(G190gat), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n606), .A2(new_n611), .A3(new_n271), .A4(new_n608), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n613), .A2(G218gat), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(G218gat), .B1(new_n613), .B2(new_n614), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT101), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n610), .B1(new_n609), .B2(new_n559), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT17), .B1(new_n501), .B2(new_n502), .ZN(new_n619));
  NOR4_X1   g418(.A1(new_n619), .A2(new_n583), .A3(KEYINPUT100), .A4(new_n496), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n271), .B1(new_n621), .B2(new_n608), .ZN(new_n622));
  INV_X1    g421(.A(new_n614), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n206), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT101), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n613), .A2(G218gat), .A3(new_n614), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G134gat), .B(G162gat), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n617), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n630), .ZN(new_n632));
  OAI211_X1 g431(.A(KEYINPUT101), .B(new_n632), .C1(new_n615), .C2(new_n616), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n577), .A2(KEYINPUT21), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n495), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(G183gat), .ZN(new_n638));
  NAND2_X1  g437(.A1(G231gat), .A2(G233gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G127gat), .B(G155gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(G211gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n640), .B(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n577), .A2(KEYINPUT21), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n643), .B(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n635), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n604), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n650), .A2(new_n402), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(new_n486), .ZN(G1324gat));
  INV_X1    g451(.A(new_n650), .ZN(new_n653));
  NAND2_X1  g452(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n484), .A2(new_n487), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n653), .A2(new_n371), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n657));
  OR3_X1    g456(.A1(new_n656), .A2(KEYINPUT105), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n487), .B1(new_n653), .B2(new_n371), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n659), .B1(new_n657), .B2(new_n656), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT105), .B1(new_n656), .B2(new_n657), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n658), .A2(new_n660), .A3(new_n661), .ZN(G1325gat));
  NOR3_X1   g461(.A1(new_n650), .A2(new_n480), .A3(new_n444), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n653), .A2(new_n410), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n663), .B1(new_n480), .B2(new_n664), .ZN(G1326gat));
  NOR2_X1   g464(.A1(new_n650), .A2(new_n250), .ZN(new_n666));
  XOR2_X1   g465(.A(KEYINPUT43), .B(G22gat), .Z(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(G1327gat));
  AOI21_X1  g467(.A(new_n634), .B1(new_n422), .B2(new_n447), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n648), .A2(new_n603), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n672), .A2(G29gat), .A3(new_n402), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n673), .B(KEYINPUT45), .Z(new_n674));
  NAND2_X1  g473(.A1(new_n448), .A2(new_n635), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n669), .A2(KEYINPUT44), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(new_n671), .ZN(new_n680));
  OAI21_X1  g479(.A(G29gat), .B1(new_n680), .B2(new_n402), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n674), .A2(new_n681), .ZN(G1328gat));
  OAI21_X1  g481(.A(G36gat), .B1(new_n680), .B2(new_n372), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n672), .A2(G36gat), .A3(new_n372), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT46), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n685), .ZN(G1329gat));
  INV_X1    g485(.A(new_n410), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n452), .B1(new_n672), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n444), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(G43gat), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n688), .B1(new_n680), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g491(.A1(new_n677), .A2(new_n445), .A3(new_n671), .A4(new_n678), .ZN(new_n693));
  AOI21_X1  g492(.A(KEYINPUT106), .B1(new_n693), .B2(G50gat), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT48), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n672), .A2(G50gat), .A3(new_n250), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n697), .B1(new_n693), .B2(G50gat), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n696), .B(new_n698), .ZN(G1331gat));
  NOR2_X1   g498(.A1(new_n601), .A2(new_n595), .ZN(new_n700));
  OR2_X1    g499(.A1(new_n596), .A2(KEYINPUT104), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n700), .B1(new_n701), .B2(new_n597), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n702), .B1(new_n422), .B2(new_n447), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n532), .B1(new_n531), .B2(new_n533), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n521), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n635), .A2(new_n648), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n708), .A2(new_n402), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(new_n560), .ZN(G1332gat));
  AOI211_X1 g509(.A(new_n372), .B(new_n708), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n711));
  NOR2_X1   g510(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1333gat));
  NAND3_X1  g512(.A1(new_n703), .A2(new_n410), .A3(new_n707), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(KEYINPUT107), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n703), .A2(new_n716), .A3(new_n410), .A4(new_n707), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n715), .A2(new_n567), .A3(new_n717), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n703), .A2(G71gat), .A3(new_n689), .A4(new_n707), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT108), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT108), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n718), .A2(new_n722), .A3(new_n719), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n721), .A2(KEYINPUT50), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(KEYINPUT50), .B1(new_n721), .B2(new_n723), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(G1334gat));
  NOR2_X1   g525(.A1(new_n708), .A2(new_n250), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(new_n568), .ZN(G1335gat));
  NAND2_X1  g527(.A1(new_n648), .A2(new_n535), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT109), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n602), .ZN(new_n731));
  XOR2_X1   g530(.A(new_n731), .B(KEYINPUT110), .Z(new_n732));
  AND2_X1   g531(.A1(new_n679), .A2(new_n732), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n733), .A2(G85gat), .ZN(new_n734));
  INV_X1    g533(.A(new_n402), .ZN(new_n735));
  INV_X1    g534(.A(new_n730), .ZN(new_n736));
  OAI21_X1  g535(.A(KEYINPUT51), .B1(new_n675), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT51), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n669), .A2(new_n738), .A3(new_n730), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n740), .A2(new_n735), .A3(new_n602), .ZN(new_n741));
  AOI22_X1  g540(.A1(new_n734), .A2(new_n735), .B1(new_n541), .B2(new_n741), .ZN(G1336gat));
  NAND4_X1  g541(.A1(new_n679), .A2(G92gat), .A3(new_n371), .A4(new_n732), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n737), .A2(new_n602), .A3(new_n371), .A4(new_n739), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n357), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT52), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT111), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n743), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  OR2_X1    g547(.A1(new_n746), .A2(KEYINPUT111), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1337gat));
  AND2_X1   g549(.A1(new_n733), .A2(new_n689), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n740), .A2(new_n328), .A3(new_n602), .ZN(new_n752));
  OAI22_X1  g551(.A1(new_n751), .A2(new_n328), .B1(new_n687), .B2(new_n752), .ZN(G1338gat));
  NAND3_X1  g552(.A1(new_n740), .A2(new_n245), .A3(new_n602), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n754), .A2(new_n250), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n679), .A2(new_n445), .A3(new_n732), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n756), .A2(G106gat), .ZN(new_n757));
  OAI21_X1  g556(.A(KEYINPUT53), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(G106gat), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT53), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n759), .B(new_n760), .C1(new_n250), .C2(new_n754), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n758), .A2(new_n761), .ZN(G1339gat));
  INV_X1    g561(.A(new_n648), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n508), .A2(new_n509), .A3(new_n507), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n499), .B1(new_n498), .B2(new_n504), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n516), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n521), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n602), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n582), .A2(new_n584), .A3(new_n589), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n770), .A2(new_n600), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n595), .B1(new_n771), .B2(KEYINPUT54), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n773));
  XNOR2_X1  g572(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n600), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n772), .A2(new_n773), .A3(KEYINPUT55), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n701), .A2(new_n597), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n582), .A2(new_n584), .A3(new_n589), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n587), .A2(KEYINPUT54), .A3(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n595), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n779), .A2(new_n780), .A3(new_n775), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n779), .A2(KEYINPUT55), .A3(new_n780), .A4(new_n775), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT113), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n776), .A2(new_n777), .A3(new_n783), .A4(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n769), .B1(new_n535), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI211_X1 g588(.A(KEYINPUT115), .B(new_n769), .C1(new_n535), .C2(new_n786), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(new_n634), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n767), .A2(KEYINPUT114), .ZN(new_n792));
  AND4_X1   g591(.A1(new_n777), .A2(new_n776), .A3(new_n783), .A4(new_n785), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n631), .A2(new_n633), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n767), .A2(KEYINPUT114), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n763), .B1(new_n791), .B2(new_n797), .ZN(new_n798));
  NOR4_X1   g597(.A1(new_n635), .A2(new_n648), .A3(new_n602), .A4(new_n706), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n800), .A2(new_n445), .A3(new_n687), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n371), .A2(new_n402), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(G113gat), .B1(new_n803), .B2(new_n535), .ZN(new_n804));
  NOR4_X1   g603(.A1(new_n800), .A2(new_n402), .A3(new_n371), .A4(new_n347), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n805), .A2(new_n292), .A3(new_n706), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(G1340gat));
  OAI21_X1  g606(.A(G120gat), .B1(new_n803), .B2(new_n702), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n805), .A2(new_n290), .A3(new_n602), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(G1341gat));
  NOR3_X1   g609(.A1(new_n803), .A2(new_n295), .A3(new_n648), .ZN(new_n811));
  AOI21_X1  g610(.A(G127gat), .B1(new_n805), .B2(new_n763), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n811), .A2(new_n812), .ZN(G1342gat));
  XOR2_X1   g612(.A(KEYINPUT72), .B(G134gat), .Z(new_n814));
  NAND3_X1  g613(.A1(new_n805), .A2(new_n635), .A3(new_n814), .ZN(new_n815));
  XOR2_X1   g614(.A(new_n815), .B(KEYINPUT56), .Z(new_n816));
  OAI21_X1  g615(.A(G134gat), .B1(new_n803), .B2(new_n634), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(G1343gat));
  AND3_X1   g617(.A1(new_n776), .A2(new_n777), .A3(new_n785), .ZN(new_n819));
  XOR2_X1   g618(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n820));
  NAND2_X1  g619(.A1(new_n781), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n706), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n768), .A2(new_n602), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT116), .B1(new_n702), .B2(new_n767), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI22_X1  g625(.A1(new_n822), .A2(new_n826), .B1(new_n631), .B2(new_n633), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n648), .B1(new_n827), .B2(new_n796), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n649), .A2(new_n702), .A3(new_n535), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT57), .B1(new_n830), .B2(new_n250), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n832), .B(new_n445), .C1(new_n798), .C2(new_n799), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n442), .A2(new_n802), .A3(new_n443), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n831), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(G141gat), .B1(new_n835), .B2(new_n535), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT58), .ZN(new_n837));
  INV_X1    g636(.A(new_n834), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n838), .A2(new_n800), .A3(new_n250), .ZN(new_n839));
  INV_X1    g638(.A(G141gat), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n839), .A2(new_n840), .A3(new_n706), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n836), .A2(new_n837), .A3(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n843));
  INV_X1    g642(.A(new_n833), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n250), .B1(new_n828), .B2(new_n829), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n834), .B1(new_n845), .B2(new_n832), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n843), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n831), .A2(KEYINPUT118), .A3(new_n833), .A4(new_n834), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n535), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n841), .B1(new_n849), .B2(new_n840), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT119), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n850), .A2(new_n851), .A3(KEYINPUT58), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n851), .B1(new_n850), .B2(KEYINPUT58), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n842), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI211_X1 g655(.A(KEYINPUT120), .B(new_n842), .C1(new_n852), .C2(new_n853), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(G1344gat));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859));
  AOI211_X1 g658(.A(new_n859), .B(G148gat), .C1(new_n839), .C2(new_n602), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n847), .A2(new_n848), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n859), .B1(new_n862), .B2(new_n702), .ZN(new_n863));
  OAI211_X1 g662(.A(KEYINPUT57), .B(new_n445), .C1(new_n798), .C2(new_n799), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n864), .B1(KEYINPUT57), .B2(new_n845), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n602), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(KEYINPUT59), .A3(new_n834), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n860), .B1(new_n869), .B2(G148gat), .ZN(G1345gat));
  AOI21_X1  g669(.A(G155gat), .B1(new_n839), .B2(new_n763), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n862), .A2(new_n648), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n871), .B1(new_n872), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g672(.A(G162gat), .B1(new_n839), .B2(new_n635), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n862), .A2(new_n634), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n874), .B1(new_n875), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g675(.A1(new_n372), .A2(new_n735), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n801), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(G169gat), .B1(new_n878), .B2(new_n535), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT122), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n402), .B1(new_n798), .B2(new_n799), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT121), .ZN(new_n882));
  AND4_X1   g681(.A1(new_n371), .A2(new_n882), .A3(new_n346), .A4(new_n250), .ZN(new_n883));
  INV_X1    g682(.A(G169gat), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n883), .A2(new_n884), .A3(new_n706), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n880), .A2(new_n885), .ZN(G1348gat));
  AOI21_X1  g685(.A(G176gat), .B1(new_n883), .B2(new_n602), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n878), .A2(new_n702), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(G176gat), .B2(new_n888), .ZN(G1349gat));
  INV_X1    g688(.A(new_n306), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n883), .A2(new_n763), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(G183gat), .B1(new_n878), .B2(new_n648), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT60), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n894), .A2(KEYINPUT123), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n893), .B(new_n895), .ZN(G1350gat));
  OAI21_X1  g695(.A(G190gat), .B1(new_n878), .B2(new_n634), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT61), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n883), .A2(new_n271), .A3(new_n635), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1351gat));
  AND2_X1   g699(.A1(new_n444), .A2(new_n877), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n865), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(G197gat), .B1(new_n902), .B2(new_n535), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n444), .A2(new_n371), .A3(new_n445), .ZN(new_n904));
  XOR2_X1   g703(.A(new_n904), .B(KEYINPUT124), .Z(new_n905));
  AND2_X1   g704(.A1(new_n905), .A2(new_n882), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT125), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n535), .A2(G197gat), .ZN(new_n908));
  AND3_X1   g707(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n907), .B1(new_n906), .B2(new_n908), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n903), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(KEYINPUT126), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT126), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n903), .B(new_n913), .C1(new_n909), .C2(new_n910), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(G1352gat));
  INV_X1    g714(.A(G204gat), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n906), .A2(new_n916), .A3(new_n602), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT62), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n916), .B1(new_n867), .B2(new_n901), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n918), .A2(new_n919), .ZN(G1353gat));
  INV_X1    g719(.A(KEYINPUT127), .ZN(new_n921));
  OAI221_X1 g720(.A(G211gat), .B1(new_n921), .B2(KEYINPUT63), .C1(new_n902), .C2(new_n648), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(KEYINPUT63), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n922), .B(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n906), .A2(new_n205), .A3(new_n763), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1354gat));
  NAND3_X1  g725(.A1(new_n906), .A2(new_n206), .A3(new_n635), .ZN(new_n927));
  OAI21_X1  g726(.A(G218gat), .B1(new_n902), .B2(new_n634), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(G1355gat));
endmodule


