//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 1 0 1 0 1 0 1 0 0 1 1 1 0 1 1 1 0 1 1 1 0 1 1 1 1 1 1 1 1 1 1 1 1 0 0 0 0 0 1 0 1 1 1 0 0 0 0 0 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n577, new_n578, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n631, new_n632, new_n635, new_n636, new_n638, new_n639, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1214,
    new_n1215, new_n1216, new_n1217;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT66), .Z(new_n451));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  XOR2_X1   g029(.A(G325), .B(KEYINPUT67), .Z(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G567), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT68), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(KEYINPUT68), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n463), .A2(new_n468), .A3(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(KEYINPUT69), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n471), .A2(new_n474), .A3(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n461), .A2(new_n462), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n465), .A2(G2105), .ZN(new_n479));
  AOI22_X1  g054(.A1(new_n478), .A2(G137), .B1(G101), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n476), .A2(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n466), .A2(new_n467), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n478), .A2(G136), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n488), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n485), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  OAI211_X1 g066(.A(G126), .B(G2105), .C1(new_n461), .C2(new_n462), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT70), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n492), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n488), .A2(KEYINPUT4), .A3(G138), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n477), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n463), .A2(new_n468), .A3(G138), .A4(new_n488), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT71), .A2(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT71), .A2(G651), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT6), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n508), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G50), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n518), .B1(new_n511), .B2(new_n513), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G88), .ZN(new_n520));
  NAND2_X1  g095(.A1(G75), .A2(G543), .ZN(new_n521));
  INV_X1    g096(.A(G62), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n521), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n509), .A2(new_n510), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  AND3_X1   g101(.A1(new_n515), .A2(new_n520), .A3(new_n526), .ZN(G166));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT74), .ZN(new_n529));
  XOR2_X1   g104(.A(KEYINPUT73), .B(KEYINPUT7), .Z(new_n530));
  XNOR2_X1  g105(.A(new_n529), .B(new_n530), .ZN(new_n531));
  OR2_X1    g106(.A1(KEYINPUT5), .A2(G543), .ZN(new_n532));
  NAND2_X1  g107(.A1(KEYINPUT5), .A2(G543), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n534), .A2(G63), .A3(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(G89), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT6), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT71), .ZN(new_n539));
  INV_X1    g114(.A(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(KEYINPUT71), .A2(G651), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n538), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n534), .B1(new_n543), .B2(new_n512), .ZN(new_n544));
  OAI21_X1  g119(.A(G543), .B1(new_n543), .B2(new_n512), .ZN(new_n545));
  XNOR2_X1  g120(.A(KEYINPUT72), .B(G51), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n537), .A2(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n536), .A2(new_n547), .ZN(G168));
  INV_X1    g123(.A(G64), .ZN(new_n549));
  INV_X1    g124(.A(G77), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n518), .A2(new_n549), .B1(new_n550), .B2(new_n508), .ZN(new_n551));
  AOI22_X1  g126(.A1(G52), .A2(new_n514), .B1(new_n551), .B2(new_n525), .ZN(new_n552));
  OAI211_X1 g127(.A(G90), .B(new_n534), .C1(new_n543), .C2(new_n512), .ZN(new_n553));
  AOI21_X1  g128(.A(KEYINPUT75), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  OAI211_X1 g129(.A(G52), .B(G543), .C1(new_n543), .C2(new_n512), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n549), .B1(new_n532), .B2(new_n533), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n550), .A2(new_n508), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n525), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n553), .A2(new_n555), .A3(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n554), .A2(new_n561), .ZN(G301));
  INV_X1    g137(.A(G301), .ZN(G171));
  XOR2_X1   g138(.A(KEYINPUT76), .B(G81), .Z(new_n564));
  OAI211_X1 g139(.A(new_n534), .B(new_n564), .C1(new_n543), .C2(new_n512), .ZN(new_n565));
  OAI211_X1 g140(.A(G43), .B(G543), .C1(new_n543), .C2(new_n512), .ZN(new_n566));
  INV_X1    g141(.A(G56), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n567), .B1(new_n532), .B2(new_n533), .ZN(new_n568));
  INV_X1    g143(.A(G68), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n569), .A2(new_n508), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n525), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n565), .A2(new_n566), .A3(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G860), .ZN(G153));
  NAND4_X1  g149(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT77), .ZN(G176));
  NAND2_X1  g151(.A1(G1), .A2(G3), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT8), .ZN(new_n578));
  NAND4_X1  g153(.A1(G319), .A2(G483), .A3(G661), .A4(new_n578), .ZN(G188));
  AND2_X1   g154(.A1(G78), .A2(G543), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n580), .B1(new_n534), .B2(G65), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT78), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(G65), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(new_n532), .B2(new_n533), .ZN(new_n585));
  OAI21_X1  g160(.A(KEYINPUT78), .B1(new_n585), .B2(new_n580), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n583), .A2(G651), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n519), .A2(G91), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT9), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n514), .A2(new_n589), .A3(G53), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n589), .B1(new_n514), .B2(G53), .ZN(new_n592));
  OAI211_X1 g167(.A(new_n587), .B(new_n588), .C1(new_n591), .C2(new_n592), .ZN(G299));
  INV_X1    g168(.A(G168), .ZN(G286));
  NAND3_X1  g169(.A1(new_n515), .A2(new_n520), .A3(new_n526), .ZN(G303));
  NAND2_X1  g170(.A1(new_n514), .A2(G49), .ZN(new_n596));
  OAI211_X1 g171(.A(G87), .B(new_n534), .C1(new_n543), .C2(new_n512), .ZN(new_n597));
  OAI21_X1  g172(.A(G651), .B1(new_n534), .B2(G74), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(G288));
  NAND2_X1  g174(.A1(new_n519), .A2(G86), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n514), .A2(G48), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n534), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT79), .ZN(new_n603));
  NOR3_X1   g178(.A1(new_n602), .A2(new_n603), .A3(new_n524), .ZN(new_n604));
  NAND2_X1  g179(.A1(G73), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G61), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n518), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g182(.A(KEYINPUT79), .B1(new_n607), .B2(new_n525), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n600), .B(new_n601), .C1(new_n604), .C2(new_n608), .ZN(G305));
  OAI211_X1 g184(.A(G85), .B(new_n534), .C1(new_n543), .C2(new_n512), .ZN(new_n610));
  INV_X1    g185(.A(G60), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n611), .B1(new_n532), .B2(new_n533), .ZN(new_n612));
  INV_X1    g187(.A(G72), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n613), .A2(new_n508), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n525), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(G47), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n610), .B(new_n615), .C1(new_n545), .C2(new_n616), .ZN(G290));
  NAND2_X1  g192(.A1(G79), .A2(G543), .ZN(new_n618));
  INV_X1    g193(.A(G66), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n518), .B2(new_n619), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n514), .A2(G54), .B1(new_n620), .B2(G651), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT80), .B(KEYINPUT10), .ZN(new_n622));
  INV_X1    g197(.A(G92), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n544), .B2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(new_n622), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n519), .A2(G92), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n621), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n627), .A2(G868), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(G171), .B2(G868), .ZN(G284));
  AOI21_X1  g204(.A(new_n628), .B1(G171), .B2(G868), .ZN(G321));
  NAND2_X1  g205(.A1(G286), .A2(G868), .ZN(new_n631));
  INV_X1    g206(.A(G299), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(G868), .B2(new_n632), .ZN(G280));
  XNOR2_X1  g208(.A(G280), .B(KEYINPUT81), .ZN(G297));
  INV_X1    g209(.A(new_n627), .ZN(new_n635));
  INV_X1    g210(.A(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(G860), .ZN(G148));
  NAND2_X1  g212(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G868), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(G868), .B2(new_n573), .ZN(G323));
  XNOR2_X1  g215(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g216(.A1(new_n463), .A2(new_n468), .ZN(new_n642));
  NOR3_X1   g217(.A1(new_n642), .A2(new_n465), .A3(G2105), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT83), .B(KEYINPUT13), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n647), .A2(G2100), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(G2100), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n484), .A2(G123), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n478), .A2(G135), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n488), .A2(G111), .ZN(new_n652));
  OAI21_X1  g227(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n653));
  OAI211_X1 g228(.A(new_n650), .B(new_n651), .C1(new_n652), .C2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(KEYINPUT84), .B(G2096), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n648), .A2(new_n649), .A3(new_n656), .ZN(G156));
  XOR2_X1   g232(.A(G1341), .B(G1348), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT85), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2451), .B(G2454), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n659), .B(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT14), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2427), .B(G2438), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2430), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT15), .B(G2435), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n663), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n667), .B1(new_n666), .B2(new_n665), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n662), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2443), .B(G2446), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n671), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n672), .A2(G14), .A3(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT86), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G401));
  XNOR2_X1  g251(.A(G2072), .B(G2078), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT87), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT88), .B(KEYINPUT18), .Z(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G2084), .B(G2090), .Z(new_n681));
  XNOR2_X1  g256(.A(G2067), .B(G2678), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n678), .B1(new_n680), .B2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n683), .ZN(new_n685));
  OAI21_X1  g260(.A(KEYINPUT17), .B1(new_n681), .B2(new_n682), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n679), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n684), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G2096), .B(G2100), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(G227));
  XNOR2_X1  g265(.A(G1971), .B(G1976), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT19), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G1956), .B(G2474), .Z(new_n694));
  XOR2_X1   g269(.A(G1961), .B(G1966), .Z(new_n695));
  AND2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT20), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n694), .A2(new_n695), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  MUX2_X1   g276(.A(new_n701), .B(new_n700), .S(new_n693), .Z(new_n702));
  NOR2_X1   g277(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1991), .B(G1996), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(G1981), .B(G1986), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(G229));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G33), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n488), .A2(G103), .A3(G2104), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT25), .ZN(new_n714));
  INV_X1    g289(.A(new_n642), .ZN(new_n715));
  AOI22_X1  g290(.A1(new_n715), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n716), .A2(new_n488), .ZN(new_n717));
  AOI211_X1 g292(.A(new_n714), .B(new_n717), .C1(G139), .C2(new_n478), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n712), .B1(new_n718), .B2(new_n711), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(G2072), .Z(new_n720));
  NOR2_X1   g295(.A1(G5), .A2(G16), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G171), .B2(G16), .ZN(new_n722));
  INV_X1    g297(.A(G1961), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G16), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G21), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G168), .B2(new_n725), .ZN(new_n727));
  INV_X1    g302(.A(G1966), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n711), .A2(G26), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT28), .Z(new_n731));
  NAND2_X1  g306(.A1(new_n484), .A2(G128), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n478), .A2(G140), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n488), .A2(G116), .ZN(new_n734));
  OAI21_X1  g309(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n732), .B(new_n733), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n731), .B1(new_n736), .B2(G29), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(G2067), .Z(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT30), .B(G28), .ZN(new_n739));
  OR2_X1    g314(.A1(KEYINPUT31), .A2(G11), .ZN(new_n740));
  NAND2_X1  g315(.A1(KEYINPUT31), .A2(G11), .ZN(new_n741));
  AOI22_X1  g316(.A1(new_n739), .A2(new_n711), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n654), .B2(new_n711), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n711), .A2(G32), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n478), .A2(G141), .B1(G105), .B2(new_n479), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n484), .A2(G129), .ZN(new_n746));
  NAND3_X1  g321(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT26), .Z(new_n748));
  NAND3_X1  g323(.A1(new_n745), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n744), .B1(new_n749), .B2(G29), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT27), .B(G1996), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n743), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n750), .B2(new_n751), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n725), .A2(G19), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n573), .B2(new_n725), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G1341), .ZN(new_n756));
  NOR3_X1   g331(.A1(new_n738), .A2(new_n753), .A3(new_n756), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n720), .A2(new_n724), .A3(new_n729), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n711), .A2(G35), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G162), .B2(new_n711), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT29), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G2090), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT95), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n725), .A2(G20), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT23), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n632), .B2(new_n725), .ZN(new_n766));
  INV_X1    g341(.A(G1956), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n711), .A2(G27), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G164), .B2(new_n711), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G2078), .ZN(new_n771));
  INV_X1    g346(.A(new_n761), .ZN(new_n772));
  INV_X1    g347(.A(G2090), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT24), .ZN(new_n775));
  INV_X1    g350(.A(G34), .ZN(new_n776));
  AOI21_X1  g351(.A(G29), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n775), .B2(new_n776), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G160), .B2(new_n711), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n779), .A2(G2084), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n763), .A2(new_n768), .A3(new_n774), .A4(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(G4), .A2(G16), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n635), .B2(G16), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT93), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G1348), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n779), .A2(G2084), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT94), .Z(new_n787));
  NOR4_X1   g362(.A1(new_n758), .A2(new_n781), .A3(new_n785), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n725), .A2(G22), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G166), .B2(new_n725), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT90), .B(G1971), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n725), .A2(G6), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G305), .B2(G16), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT32), .B(G1981), .Z(new_n795));
  OR2_X1    g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n795), .B2(new_n794), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n725), .A2(G23), .ZN(new_n799));
  INV_X1    g374(.A(G288), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n725), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT33), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1976), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n798), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(KEYINPUT34), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT34), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n798), .A2(new_n803), .A3(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(G16), .A2(G24), .ZN(new_n808));
  XOR2_X1   g383(.A(G290), .B(KEYINPUT89), .Z(new_n809));
  AOI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(G16), .ZN(new_n810));
  INV_X1    g385(.A(G1986), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n711), .A2(G25), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n478), .A2(G131), .ZN(new_n814));
  OR2_X1    g389(.A1(G95), .A2(G2105), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n815), .B(G2104), .C1(G107), .C2(new_n488), .ZN(new_n816));
  INV_X1    g391(.A(G119), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n814), .B(new_n816), .C1(new_n817), .C2(new_n483), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n813), .B1(new_n819), .B2(new_n711), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT35), .B(G1991), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n805), .A2(new_n807), .A3(new_n812), .A4(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT91), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n824), .A2(KEYINPUT36), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(KEYINPUT36), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT92), .Z(new_n827));
  AND3_X1   g402(.A1(new_n823), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n827), .B1(new_n823), .B2(new_n825), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n788), .B1(new_n828), .B2(new_n829), .ZN(G150));
  INV_X1    g405(.A(KEYINPUT96), .ZN(new_n831));
  XNOR2_X1  g406(.A(G150), .B(new_n831), .ZN(G311));
  NOR2_X1   g407(.A1(new_n627), .A2(new_n636), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT38), .ZN(new_n834));
  OAI22_X1  g409(.A1(new_n518), .A2(new_n567), .B1(new_n569), .B2(new_n508), .ZN(new_n835));
  AOI22_X1  g410(.A1(G43), .A2(new_n514), .B1(new_n835), .B2(new_n525), .ZN(new_n836));
  NAND2_X1  g411(.A1(G80), .A2(G543), .ZN(new_n837));
  INV_X1    g412(.A(G67), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n837), .B1(new_n518), .B2(new_n838), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n514), .A2(G55), .B1(new_n839), .B2(new_n525), .ZN(new_n840));
  OAI211_X1 g415(.A(G93), .B(new_n534), .C1(new_n543), .C2(new_n512), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n836), .A2(new_n840), .A3(new_n565), .A4(new_n841), .ZN(new_n842));
  OAI211_X1 g417(.A(G55), .B(G543), .C1(new_n543), .C2(new_n512), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n838), .B1(new_n532), .B2(new_n533), .ZN(new_n844));
  INV_X1    g419(.A(new_n837), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n525), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n841), .A2(new_n843), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n572), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n842), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n834), .B(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n850), .A2(KEYINPUT39), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(KEYINPUT39), .ZN(new_n852));
  XOR2_X1   g427(.A(KEYINPUT97), .B(G860), .Z(new_n853));
  NAND3_X1  g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n847), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n855), .A2(new_n853), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT37), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n854), .A2(new_n857), .ZN(G145));
  INV_X1    g433(.A(G37), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n736), .B(new_n749), .Z(new_n860));
  NAND2_X1  g435(.A1(new_n503), .A2(new_n504), .ZN(new_n861));
  INV_X1    g436(.A(new_n502), .ZN(new_n862));
  INV_X1    g437(.A(new_n496), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n860), .B(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n718), .ZN(new_n866));
  AOI22_X1  g441(.A1(new_n484), .A2(G130), .B1(new_n478), .B2(G142), .ZN(new_n867));
  OAI21_X1  g442(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n868));
  INV_X1    g443(.A(G118), .ZN(new_n869));
  AOI22_X1  g444(.A1(new_n868), .A2(KEYINPUT98), .B1(new_n869), .B2(G2105), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n870), .B1(KEYINPUT98), .B2(new_n868), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n819), .B(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n645), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n866), .B(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(G160), .B(new_n654), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n490), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n859), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(KEYINPUT99), .B1(new_n866), .B2(new_n874), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n866), .A2(new_n874), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n866), .A2(KEYINPUT99), .A3(new_n874), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n877), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n879), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT40), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(G395));
  INV_X1    g462(.A(KEYINPUT104), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n849), .B(KEYINPUT100), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n638), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT41), .ZN(new_n891));
  NOR2_X1   g466(.A1(G299), .A2(new_n627), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n621), .A2(new_n624), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n540), .B1(new_n581), .B2(new_n582), .ZN(new_n894));
  AOI22_X1  g469(.A1(new_n894), .A2(new_n586), .B1(G91), .B2(new_n519), .ZN(new_n895));
  INV_X1    g470(.A(G53), .ZN(new_n896));
  OAI21_X1  g471(.A(KEYINPUT9), .B1(new_n545), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(new_n590), .ZN(new_n898));
  AOI22_X1  g473(.A1(new_n893), .A2(new_n626), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n891), .B1(new_n892), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n635), .A2(new_n898), .A3(new_n895), .ZN(new_n901));
  NAND2_X1  g476(.A1(G299), .A2(new_n627), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(KEYINPUT41), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n890), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT101), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(new_n892), .B2(new_n899), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n901), .A2(KEYINPUT101), .A3(new_n902), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n890), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n905), .A2(KEYINPUT103), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(KEYINPUT103), .B1(new_n905), .B2(new_n910), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT102), .ZN(new_n913));
  AND2_X1   g488(.A1(G288), .A2(G290), .ZN(new_n914));
  NOR2_X1   g489(.A1(G288), .A2(G290), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n597), .A2(new_n598), .ZN(new_n917));
  OAI22_X1  g492(.A1(new_n518), .A2(new_n611), .B1(new_n613), .B2(new_n508), .ZN(new_n918));
  AOI22_X1  g493(.A1(G47), .A2(new_n514), .B1(new_n918), .B2(new_n525), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n917), .A2(new_n919), .A3(new_n596), .A4(new_n610), .ZN(new_n920));
  NAND2_X1  g495(.A1(G288), .A2(G290), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(new_n921), .A3(KEYINPUT102), .ZN(new_n922));
  NAND2_X1  g497(.A1(G305), .A2(G303), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n603), .B1(new_n602), .B2(new_n524), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n607), .A2(KEYINPUT79), .A3(new_n525), .ZN(new_n925));
  AOI22_X1  g500(.A1(new_n924), .A2(new_n925), .B1(G48), .B2(new_n514), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n926), .A2(G166), .A3(new_n600), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n916), .A2(new_n922), .A3(new_n923), .A4(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n923), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n914), .A2(new_n915), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(KEYINPUT102), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(KEYINPUT42), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n911), .B1(new_n912), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n933), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n905), .A2(new_n935), .A3(KEYINPUT103), .A4(new_n910), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(G868), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n855), .A2(G868), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n888), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  AOI211_X1 g516(.A(KEYINPUT104), .B(new_n939), .C1(new_n937), .C2(G868), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(G295));
  NAND2_X1  g518(.A1(new_n938), .A2(new_n940), .ZN(G331));
  NAND3_X1  g519(.A1(new_n552), .A2(KEYINPUT75), .A3(new_n553), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n559), .A2(new_n560), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n572), .A2(new_n847), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n572), .A2(new_n847), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n945), .B(new_n946), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n842), .B(new_n848), .C1(new_n554), .C2(new_n561), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n949), .A2(G168), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(G168), .B1(new_n949), .B2(new_n950), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n900), .B(new_n903), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n932), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n949), .A2(new_n950), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(G286), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n892), .A2(new_n899), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n949), .A2(new_n950), .A3(G168), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n953), .A2(new_n954), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n859), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT105), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n932), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n928), .A2(new_n931), .A3(KEYINPUT105), .ZN(new_n964));
  AOI22_X1  g539(.A1(new_n953), .A2(new_n959), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT43), .B1(new_n961), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n909), .A2(new_n958), .A3(new_n956), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n953), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n963), .A2(new_n964), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT43), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n970), .A2(new_n971), .A3(new_n859), .A4(new_n960), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n966), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n953), .A2(new_n967), .B1(new_n963), .B2(new_n964), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT106), .B1(new_n961), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT106), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n970), .A2(new_n978), .A3(new_n859), .A4(new_n960), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n977), .A2(new_n979), .A3(KEYINPUT43), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n961), .A2(new_n965), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n974), .B1(new_n981), .B2(new_n971), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n980), .A2(new_n982), .A3(KEYINPUT107), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT107), .B1(new_n980), .B2(new_n982), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n975), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT108), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI211_X1 g562(.A(KEYINPUT108), .B(new_n975), .C1(new_n983), .C2(new_n984), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(G397));
  INV_X1    g564(.A(G1384), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n864), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n480), .A2(G40), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n474), .B1(new_n471), .B2(G2105), .ZN(new_n995));
  AOI211_X1 g570(.A(KEYINPUT69), .B(new_n488), .C1(new_n469), .C2(new_n470), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n994), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n993), .A2(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n736), .B(G2067), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n999), .B(KEYINPUT110), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n749), .B(G1996), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OR2_X1    g578(.A1(new_n819), .A2(new_n821), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n819), .A2(new_n821), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G290), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n811), .ZN(new_n1008));
  XOR2_X1   g583(.A(new_n1008), .B(KEYINPUT109), .Z(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1010), .B1(new_n811), .B2(new_n1007), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n998), .B1(new_n1006), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT45), .B1(new_n506), .B2(new_n990), .ZN(new_n1013));
  AOI211_X1 g588(.A(new_n992), .B(G1384), .C1(new_n505), .C2(new_n863), .ZN(new_n1014));
  NOR3_X1   g589(.A1(new_n1013), .A2(new_n1014), .A3(new_n997), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1015), .A2(G1971), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n991), .A2(KEYINPUT50), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n480), .A2(G40), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1018), .B1(new_n473), .B2(new_n475), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n506), .A2(new_n990), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1017), .B(new_n1019), .C1(KEYINPUT50), .C2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1021), .A2(G2090), .ZN(new_n1022));
  OAI21_X1  g597(.A(KEYINPUT114), .B1(new_n1016), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1020), .A2(new_n992), .ZN(new_n1024));
  AOI21_X1  g599(.A(G1384), .B1(new_n505), .B2(new_n863), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT45), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1024), .A2(new_n1019), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G1971), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1029), .B(new_n1030), .C1(G2090), .C2(new_n1021), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1023), .A2(G8), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(G303), .A2(G8), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1033), .B(KEYINPUT55), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT112), .B(G86), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n519), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n926), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(G1981), .ZN(new_n1039));
  INV_X1    g614(.A(G1981), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n926), .A2(new_n1040), .A3(new_n600), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1039), .A2(new_n1041), .A3(KEYINPUT49), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT49), .ZN(new_n1043));
  NOR2_X1   g618(.A1(G305), .A2(G1981), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1040), .B1(new_n926), .B2(new_n1037), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G8), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1047), .B1(new_n1019), .B2(new_n1025), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1042), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n800), .A2(G1976), .ZN(new_n1050));
  OAI211_X1 g625(.A(G8), .B(new_n1050), .C1(new_n997), .C2(new_n991), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT52), .ZN(new_n1052));
  INV_X1    g627(.A(G1976), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT52), .B1(G288), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1048), .A2(new_n1050), .A3(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1049), .A2(new_n1052), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT115), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT115), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1049), .A2(new_n1052), .A3(new_n1058), .A4(new_n1055), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1034), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1020), .A2(KEYINPUT50), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT50), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1025), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1062), .A2(new_n1019), .A3(new_n1064), .ZN(new_n1065));
  OAI22_X1  g640(.A1(new_n1016), .A2(KEYINPUT111), .B1(G2090), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT111), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1029), .A2(new_n1067), .ZN(new_n1068));
  OAI211_X1 g643(.A(G8), .B(new_n1061), .C1(new_n1066), .C2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n506), .A2(KEYINPUT45), .A3(new_n990), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n993), .A2(new_n1019), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n728), .ZN(new_n1072));
  INV_X1    g647(.A(G2084), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1062), .A2(new_n1073), .A3(new_n1019), .A4(new_n1064), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(G168), .A2(G8), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT116), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT116), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1078), .A2(new_n1079), .A3(G8), .A4(G168), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1035), .A2(new_n1060), .A3(new_n1069), .A4(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT63), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1065), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1029), .A2(new_n1067), .B1(new_n1085), .B2(new_n773), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1016), .A2(KEYINPUT111), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1047), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n1061), .A2(KEYINPUT117), .ZN(new_n1089));
  OR2_X1    g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1056), .A2(new_n1083), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1090), .A2(new_n1081), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1049), .A2(new_n1053), .A3(new_n800), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1048), .B1(new_n1094), .B2(new_n1044), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n1069), .B2(new_n1056), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT113), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1095), .B(KEYINPUT113), .C1(new_n1069), .C2(new_n1056), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1084), .A2(new_n1093), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT124), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1072), .A2(G168), .A3(new_n1074), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(G8), .ZN(new_n1103));
  AOI21_X1  g678(.A(G168), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT51), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT62), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT51), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1102), .A2(new_n1107), .A3(G8), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1105), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1106), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT53), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1112), .B1(new_n1027), .B2(G2078), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1065), .A2(new_n723), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1112), .A2(G2078), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1113), .B(new_n1114), .C1(new_n1071), .C2(new_n1116), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1117), .A2(G171), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1035), .A2(new_n1060), .A3(new_n1069), .A4(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1101), .B1(new_n1111), .B2(new_n1120), .ZN(new_n1121));
  NOR4_X1   g696(.A1(new_n1119), .A2(new_n1109), .A3(new_n1110), .A4(KEYINPUT124), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1100), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  OR2_X1    g698(.A1(G301), .A2(KEYINPUT54), .ZN(new_n1124));
  NAND2_X1  g699(.A1(G301), .A2(KEYINPUT54), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1117), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1026), .A2(new_n472), .A3(new_n994), .A4(new_n1115), .ZN(new_n1128));
  INV_X1    g703(.A(new_n993), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1124), .B(new_n1125), .C1(new_n1128), .C2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT123), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1114), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1065), .A2(KEYINPUT123), .A3(new_n723), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1131), .A2(new_n1113), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1127), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1136), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1137), .A2(new_n1060), .A3(new_n1069), .A4(new_n1035), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n1139));
  OAI21_X1  g714(.A(KEYINPUT118), .B1(new_n997), .B2(new_n991), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT118), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n476), .A2(new_n1141), .A3(new_n994), .A4(new_n1025), .ZN(new_n1142));
  XOR2_X1   g717(.A(KEYINPUT58), .B(G1341), .Z(new_n1143));
  NAND3_X1  g718(.A1(new_n1140), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT121), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(G1996), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1015), .A2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1140), .A2(new_n1142), .A3(KEYINPUT121), .A4(new_n1143), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1146), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT59), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1150), .A2(new_n1151), .A3(new_n573), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1151), .B1(new_n1150), .B2(new_n573), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g730(.A(KEYINPUT56), .B(G2072), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1024), .A2(new_n1019), .A3(new_n1026), .A4(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT57), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n895), .A2(new_n898), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1158), .B1(new_n895), .B2(new_n898), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AOI211_X1 g737(.A(KEYINPUT50), .B(G1384), .C1(new_n500), .C2(new_n505), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1063), .B1(new_n864), .B2(new_n990), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1163), .A2(new_n997), .A3(new_n1164), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1157), .B(new_n1162), .C1(new_n1165), .C2(G1956), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1166), .A2(KEYINPUT61), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1157), .B1(new_n1165), .B2(G1956), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT120), .ZN(new_n1169));
  OAI21_X1  g744(.A(KEYINPUT119), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1161), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT119), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1171), .A2(new_n1172), .A3(new_n1159), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1170), .A2(new_n1173), .ZN(new_n1174));
  AND3_X1   g749(.A1(new_n1168), .A2(new_n1169), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1169), .B1(new_n1168), .B2(new_n1174), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1167), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1162), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1168), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(new_n1166), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1177), .A2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1139), .B1(new_n1155), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1150), .A2(new_n573), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(KEYINPUT59), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(new_n1152), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1187), .A2(KEYINPUT122), .A3(new_n1177), .A4(new_n1182), .ZN(new_n1188));
  AOI21_X1  g763(.A(G2067), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1189));
  INV_X1    g764(.A(G1348), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1189), .B1(new_n1190), .B2(new_n1065), .ZN(new_n1191));
  AND3_X1   g766(.A1(new_n1191), .A2(KEYINPUT60), .A3(new_n627), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n627), .B1(new_n1191), .B2(KEYINPUT60), .ZN(new_n1193));
  OAI22_X1  g768(.A1(new_n1192), .A2(new_n1193), .B1(KEYINPUT60), .B2(new_n1191), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1184), .A2(new_n1188), .A3(new_n1194), .ZN(new_n1195));
  OAI22_X1  g770(.A1(new_n1175), .A2(new_n1176), .B1(new_n627), .B2(new_n1191), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1196), .A2(new_n1166), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1138), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1012), .B1(new_n1123), .B2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g774(.A(KEYINPUT48), .B1(new_n1009), .B2(new_n998), .ZN(new_n1200));
  AND3_X1   g775(.A1(new_n1009), .A2(KEYINPUT48), .A3(new_n998), .ZN(new_n1201));
  AOI211_X1 g776(.A(new_n1200), .B(new_n1201), .C1(new_n1006), .C2(new_n998), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n998), .B1(new_n1001), .B2(new_n749), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n998), .A2(new_n1147), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n1204), .B(KEYINPUT46), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1206));
  XOR2_X1   g781(.A(new_n1206), .B(KEYINPUT47), .Z(new_n1207));
  XOR2_X1   g782(.A(new_n1005), .B(KEYINPUT125), .Z(new_n1208));
  NAND2_X1  g783(.A1(new_n1003), .A2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1209), .B1(G2067), .B2(new_n736), .ZN(new_n1210));
  AOI211_X1 g785(.A(new_n1202), .B(new_n1207), .C1(new_n998), .C2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1199), .A2(new_n1211), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g787(.A1(G401), .A2(new_n458), .A3(G227), .ZN(new_n1214));
  INV_X1    g788(.A(KEYINPUT126), .ZN(new_n1215));
  AND3_X1   g789(.A1(new_n1214), .A2(new_n1215), .A3(new_n709), .ZN(new_n1216));
  AOI21_X1  g790(.A(new_n1215), .B1(new_n1214), .B2(new_n709), .ZN(new_n1217));
  OAI221_X1 g791(.A(new_n973), .B1(new_n879), .B2(new_n884), .C1(new_n1216), .C2(new_n1217), .ZN(G225));
  INV_X1    g792(.A(G225), .ZN(G308));
endmodule


