//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 0 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 0 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1225, new_n1226, new_n1227, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1290, new_n1291, new_n1292, new_n1293;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n209), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT65), .Z(new_n225));
  INV_X1    g0025(.A(KEYINPUT1), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n225), .A2(new_n226), .ZN(new_n228));
  AND3_X1   g0028(.A1(new_n217), .A2(new_n227), .A3(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G58), .B(G77), .Z(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n240), .B(KEYINPUT66), .Z(new_n241));
  XNOR2_X1  g0041(.A(G87), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G97), .B(G107), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(G179), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n206), .A2(G45), .ZN(new_n247));
  OR2_X1    g0047(.A1(KEYINPUT5), .A2(G41), .ZN(new_n248));
  NAND2_X1  g0048(.A1(KEYINPUT5), .A2(G41), .ZN(new_n249));
  AOI21_X1  g0049(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G274), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  AND2_X1   g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(new_n213), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n252), .B1(G257), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT3), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G33), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n258), .A2(new_n260), .A3(G250), .A4(G1698), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G33), .A2(G283), .ZN(new_n262));
  AND2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n258), .A2(new_n260), .A3(G244), .A4(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT4), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n258), .A2(new_n260), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n264), .A2(KEYINPUT4), .A3(G244), .ZN(new_n269));
  OAI21_X1  g0069(.A(KEYINPUT81), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT81), .ZN(new_n272));
  AND3_X1   g0072(.A1(new_n264), .A2(KEYINPUT4), .A3(G244), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n263), .A2(new_n267), .A3(new_n270), .A4(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT82), .ZN(new_n276));
  AND3_X1   g0076(.A1(new_n275), .A2(new_n276), .A3(new_n254), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n276), .B1(new_n275), .B2(new_n254), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n246), .B(new_n256), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n270), .A2(new_n262), .A3(new_n274), .A4(new_n261), .ZN(new_n280));
  INV_X1    g0080(.A(new_n267), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n254), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n256), .ZN(new_n283));
  INV_X1    g0083(.A(G169), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AND2_X1   g0085(.A1(new_n279), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT70), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT70), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n289), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n288), .A2(new_n213), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT6), .ZN(new_n292));
  INV_X1    g0092(.A(G97), .ZN(new_n293));
  NOR3_X1   g0093(.A1(new_n292), .A2(new_n293), .A3(G107), .ZN(new_n294));
  XNOR2_X1  g0094(.A(G97), .B(G107), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n294), .B1(new_n292), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G20), .A2(G33), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  OAI22_X1  g0098(.A1(new_n296), .A2(new_n207), .B1(new_n202), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G107), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n257), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT7), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(G20), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n301), .B(new_n303), .C1(new_n268), .C2(KEYINPUT79), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n302), .B1(new_n271), .B2(G20), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n300), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n291), .B1(new_n299), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n291), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n206), .A2(G33), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n310), .A2(G97), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n309), .A2(new_n293), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n307), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n256), .B1(new_n277), .B2(new_n278), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G200), .ZN(new_n316));
  INV_X1    g0116(.A(G190), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n283), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n318), .A2(new_n314), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n286), .A2(new_n314), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  AND3_X1   g0120(.A1(new_n288), .A2(new_n213), .A3(new_n290), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n308), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n206), .A2(G20), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G50), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n322), .A2(new_n324), .B1(G50), .B2(new_n308), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT73), .ZN(new_n326));
  XNOR2_X1  g0126(.A(new_n325), .B(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G58), .ZN(new_n328));
  OAI21_X1  g0128(.A(KEYINPUT71), .B1(new_n328), .B2(KEYINPUT72), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT8), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI211_X1 g0131(.A(KEYINPUT71), .B(KEYINPUT8), .C1(new_n328), .C2(KEYINPUT72), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT71), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n333), .A2(KEYINPUT8), .A3(G58), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n331), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n335), .A2(new_n207), .A3(G33), .ZN(new_n336));
  INV_X1    g0136(.A(G150), .ZN(new_n337));
  OAI22_X1  g0137(.A1(new_n337), .A2(new_n298), .B1(new_n201), .B2(new_n207), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n291), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n327), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n340), .B(KEYINPUT9), .ZN(new_n341));
  NAND2_X1  g0141(.A1(G33), .A2(G41), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(G1), .A3(G13), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT69), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n271), .A2(new_n264), .ZN(new_n345));
  INV_X1    g0145(.A(G222), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n271), .A2(KEYINPUT69), .A3(G222), .A4(new_n264), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n268), .A2(new_n264), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n350), .A2(G223), .B1(G77), .B2(new_n268), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n343), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(G41), .A2(G45), .ZN(new_n353));
  OAI22_X1  g0153(.A1(new_n253), .A2(new_n213), .B1(new_n353), .B2(G1), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT68), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT68), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n343), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G226), .ZN(new_n360));
  XNOR2_X1  g0160(.A(KEYINPUT67), .B(G45), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n206), .B(G274), .C1(new_n361), .C2(G41), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n352), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G200), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(G190), .B2(new_n364), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n341), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT74), .ZN(new_n369));
  AOI21_X1  g0169(.A(KEYINPUT10), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n341), .B(new_n367), .C1(new_n369), .C2(KEYINPUT10), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n284), .B1(new_n352), .B2(new_n363), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n364), .A2(new_n246), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n340), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n371), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n335), .A2(new_n321), .A3(new_n308), .A4(new_n323), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n331), .A2(new_n309), .A3(new_n332), .A4(new_n334), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT80), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT80), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n377), .A2(new_n381), .A3(new_n378), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G68), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n328), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(G58), .A2(G68), .ZN(new_n386));
  OAI21_X1  g0186(.A(G20), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n297), .A2(G159), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(G20), .B1(new_n258), .B2(new_n260), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT78), .B1(new_n390), .B2(KEYINPUT7), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT78), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n392), .B(new_n302), .C1(new_n271), .C2(G20), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n268), .A2(new_n303), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n391), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n389), .B1(new_n395), .B2(G68), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n321), .B1(new_n396), .B2(KEYINPUT16), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT16), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n384), .B1(new_n304), .B2(new_n305), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n398), .B1(new_n399), .B2(new_n389), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n383), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  OR2_X1    g0201(.A1(new_n264), .A2(G226), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n271), .B(new_n402), .C1(G223), .C2(G1698), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G33), .A2(G87), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n343), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(G232), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n362), .B1(new_n406), .B2(new_n354), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(G179), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n284), .B2(new_n408), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT18), .B1(new_n401), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n395), .A2(G68), .ZN(new_n413));
  INV_X1    g0213(.A(new_n389), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(KEYINPUT16), .A3(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n415), .A2(new_n291), .A3(new_n400), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n380), .A2(new_n382), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n206), .A2(G274), .ZN(new_n418));
  AND2_X1   g0218(.A1(KEYINPUT67), .A2(G45), .ZN(new_n419));
  NOR2_X1   g0219(.A1(KEYINPUT67), .A2(G45), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(G41), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n418), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n354), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n423), .B1(G232), .B2(new_n424), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n403), .A2(new_n404), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n425), .B(G190), .C1(new_n426), .C2(new_n343), .ZN(new_n427));
  OAI21_X1  g0227(.A(G200), .B1(new_n405), .B2(new_n407), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n416), .A2(new_n417), .A3(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT17), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n416), .A2(new_n417), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT18), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n433), .A2(new_n434), .A3(new_n410), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n416), .A2(new_n417), .A3(KEYINPUT17), .A4(new_n429), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n412), .A2(new_n432), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT14), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n257), .A2(new_n293), .ZN(new_n439));
  NOR2_X1   g0239(.A1(G226), .A2(G1698), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n440), .B1(new_n406), .B2(G1698), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n439), .B1(new_n441), .B2(new_n271), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n362), .B1(new_n442), .B2(new_n343), .ZN(new_n443));
  INV_X1    g0243(.A(G238), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n444), .B1(new_n355), .B2(new_n358), .ZN(new_n445));
  NOR3_X1   g0245(.A1(new_n443), .A2(new_n445), .A3(KEYINPUT13), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT13), .ZN(new_n447));
  INV_X1    g0247(.A(new_n439), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n406), .A2(G1698), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(G226), .B2(G1698), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n448), .B1(new_n450), .B2(new_n268), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n423), .B1(new_n451), .B2(new_n254), .ZN(new_n452));
  INV_X1    g0252(.A(new_n358), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n356), .B1(new_n343), .B2(new_n357), .ZN(new_n454));
  OAI21_X1  g0254(.A(G238), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n447), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n438), .B(G169), .C1(new_n446), .C2(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT13), .B1(new_n443), .B2(new_n445), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n452), .A2(new_n447), .A3(new_n455), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n458), .A2(G179), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n458), .A2(new_n459), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n438), .B1(new_n462), .B2(G169), .ZN(new_n463));
  OAI21_X1  g0263(.A(KEYINPUT77), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(G169), .B1(new_n446), .B2(new_n456), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT14), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT77), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n466), .A2(new_n467), .A3(new_n460), .A4(new_n457), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n207), .A2(G33), .ZN(new_n470));
  OAI22_X1  g0270(.A1(new_n470), .A2(new_n202), .B1(new_n207), .B2(G68), .ZN(new_n471));
  INV_X1    g0271(.A(G50), .ZN(new_n472));
  OAI22_X1  g0272(.A1(new_n471), .A2(KEYINPUT75), .B1(new_n472), .B2(new_n298), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n471), .A2(KEYINPUT75), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n291), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT76), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT11), .ZN(new_n478));
  OAI211_X1 g0278(.A(KEYINPUT76), .B(new_n291), .C1(new_n473), .C2(new_n474), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n478), .B1(new_n477), .B2(new_n479), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n310), .A2(G68), .A3(new_n323), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT12), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n483), .B1(new_n309), .B2(new_n384), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n308), .A2(KEYINPUT12), .A3(G68), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR3_X1   g0286(.A1(new_n480), .A2(new_n481), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n469), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n462), .A2(G200), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n487), .B(new_n490), .C1(new_n317), .C2(new_n462), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n423), .B1(new_n359), .B2(G244), .ZN(new_n492));
  OAI22_X1  g0292(.A1(new_n345), .A2(new_n406), .B1(new_n300), .B2(new_n271), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n493), .B1(G238), .B2(new_n350), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n492), .B1(new_n494), .B2(new_n343), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n284), .ZN(new_n496));
  XOR2_X1   g0296(.A(KEYINPUT8), .B(G58), .Z(new_n497));
  AOI22_X1  g0297(.A1(new_n497), .A2(new_n297), .B1(G20), .B2(G77), .ZN(new_n498));
  XNOR2_X1  g0298(.A(KEYINPUT15), .B(G87), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n498), .B1(new_n470), .B2(new_n499), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n500), .A2(new_n291), .B1(new_n202), .B2(new_n309), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n310), .A2(G77), .A3(new_n323), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n496), .B(new_n503), .C1(G179), .C2(new_n495), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n503), .B1(new_n495), .B2(G200), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(new_n317), .B2(new_n495), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n489), .A2(new_n491), .A3(new_n504), .A4(new_n506), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n376), .A2(new_n437), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n310), .A2(G116), .A3(new_n311), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n308), .A2(G116), .ZN(new_n510));
  XNOR2_X1  g0310(.A(new_n510), .B(KEYINPUT85), .ZN(new_n511));
  AOI21_X1  g0311(.A(G20), .B1(G33), .B2(G283), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n257), .A2(G97), .ZN(new_n513));
  INV_X1    g0313(.A(G116), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n512), .A2(new_n513), .B1(G20), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(KEYINPUT20), .B1(new_n291), .B2(new_n515), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n291), .A2(KEYINPUT20), .A3(new_n515), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n509), .B(new_n511), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n255), .A2(G270), .B1(G274), .B2(new_n250), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n258), .A2(new_n260), .A3(G257), .A4(new_n264), .ZN(new_n520));
  INV_X1    g0320(.A(G303), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n520), .B1(new_n521), .B2(new_n271), .ZN(new_n522));
  INV_X1    g0322(.A(G264), .ZN(new_n523));
  NOR3_X1   g0323(.A1(new_n268), .A2(new_n523), .A3(new_n264), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n254), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n518), .A2(new_n526), .A3(G169), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT21), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n526), .A2(G200), .ZN(new_n530));
  INV_X1    g0330(.A(new_n518), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n530), .B(new_n531), .C1(new_n317), .C2(new_n526), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n518), .A2(G179), .A3(new_n525), .A4(new_n519), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n518), .A2(new_n526), .A3(KEYINPUT21), .A4(G169), .ZN(new_n534));
  AND4_X1   g0334(.A1(new_n529), .A2(new_n532), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n206), .A2(G45), .A3(G274), .ZN(new_n536));
  INV_X1    g0336(.A(G45), .ZN(new_n537));
  OAI21_X1  g0337(.A(G250), .B1(new_n537), .B2(G1), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n536), .B1(new_n254), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT83), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n343), .A2(G250), .A3(new_n247), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT83), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n541), .A2(new_n542), .A3(new_n536), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n258), .A2(new_n260), .A3(G244), .A4(G1698), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n258), .A2(new_n260), .A3(G238), .A4(new_n264), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G33), .A2(G116), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n540), .A2(new_n543), .B1(new_n547), .B2(new_n254), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G190), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n258), .A2(new_n260), .A3(new_n207), .A4(G68), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT19), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n470), .B2(new_n293), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g0353(.A(KEYINPUT84), .B(G87), .ZN(new_n554));
  NOR2_X1   g0354(.A1(G97), .A2(G107), .ZN(new_n555));
  NAND3_X1  g0355(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n554), .A2(new_n555), .B1(new_n207), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n291), .B1(new_n553), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n499), .A2(new_n309), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n321), .A2(G87), .A3(new_n308), .A4(new_n311), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n549), .B(new_n561), .C1(new_n365), .C2(new_n548), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n310), .A2(new_n311), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n558), .B(new_n559), .C1(new_n563), .C2(new_n499), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n540), .A2(new_n543), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n547), .A2(new_n254), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(new_n246), .A3(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n564), .B(new_n567), .C1(G169), .C2(new_n548), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n562), .A2(new_n568), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n250), .A2(new_n523), .A3(new_n254), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n258), .A2(new_n260), .A3(G250), .A4(new_n264), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT86), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT86), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n271), .A2(new_n573), .A3(G250), .A4(new_n264), .ZN(new_n574));
  NAND2_X1  g0374(.A1(G33), .A2(G294), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n271), .A2(G257), .A3(G1698), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n572), .A2(new_n574), .A3(new_n575), .A4(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n570), .B1(new_n577), .B2(new_n254), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n251), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n284), .ZN(new_n580));
  AOI211_X1 g0380(.A(new_n570), .B(new_n252), .C1(new_n577), .C2(new_n254), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n246), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT24), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n258), .A2(new_n260), .A3(new_n207), .A4(G87), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT22), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT22), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n271), .A2(new_n586), .A3(new_n207), .A4(G87), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n546), .A2(G20), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT23), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(new_n207), .B2(G107), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n300), .A2(KEYINPUT23), .A3(G20), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n589), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n583), .B1(new_n588), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n588), .A2(new_n583), .A3(new_n593), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n321), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n563), .A2(new_n300), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n309), .A2(new_n300), .ZN(new_n599));
  XNOR2_X1  g0399(.A(new_n599), .B(KEYINPUT25), .ZN(new_n600));
  OR2_X1    g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n580), .B(new_n582), .C1(new_n597), .C2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n579), .A2(G200), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n581), .A2(G190), .ZN(new_n604));
  INV_X1    g0404(.A(new_n596), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n291), .B1(new_n605), .B2(new_n594), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n598), .A2(new_n600), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n603), .A2(new_n604), .A3(new_n606), .A4(new_n607), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n569), .A2(new_n602), .A3(new_n608), .ZN(new_n609));
  AND4_X1   g0409(.A1(new_n320), .A2(new_n508), .A3(new_n535), .A4(new_n609), .ZN(G372));
  INV_X1    g0410(.A(new_n375), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT88), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n504), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n504), .A2(new_n612), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n613), .A2(new_n491), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n487), .B1(new_n464), .B2(new_n468), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n432), .B(new_n436), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n412), .A2(new_n435), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n371), .A2(new_n372), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n611), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n529), .A2(new_n533), .A3(new_n534), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n602), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n569), .A2(new_n608), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n320), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n568), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n286), .A2(new_n314), .A3(new_n569), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n629), .B1(new_n630), .B2(KEYINPUT26), .ZN(new_n631));
  INV_X1    g0431(.A(new_n314), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n279), .A2(new_n285), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n632), .B1(new_n633), .B2(KEYINPUT87), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT26), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT87), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n279), .A2(new_n636), .A3(new_n285), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n634), .A2(new_n635), .A3(new_n569), .A4(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n628), .A2(new_n631), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n508), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n622), .A2(new_n640), .ZN(G369));
  NAND3_X1  g0441(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT27), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n644), .A2(new_n206), .A3(new_n207), .A4(G13), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n643), .A2(G213), .A3(new_n645), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n646), .A2(KEYINPUT89), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(KEYINPUT89), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(G343), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n651), .A2(KEYINPUT90), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(KEYINPUT90), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n597), .B2(new_n601), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n655), .A2(new_n608), .A3(new_n602), .ZN(new_n656));
  INV_X1    g0456(.A(new_n654), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n623), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n602), .B2(new_n654), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n661), .A2(KEYINPUT91), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(KEYINPUT91), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n535), .B1(new_n657), .B2(new_n531), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n654), .A2(new_n623), .A3(new_n518), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(G330), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n602), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n654), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n656), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n664), .A2(new_n677), .ZN(G399));
  NAND3_X1  g0478(.A1(new_n554), .A2(new_n514), .A3(new_n555), .ZN(new_n679));
  XOR2_X1   g0479(.A(new_n679), .B(KEYINPUT92), .Z(new_n680));
  INV_X1    g0480(.A(new_n210), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(G41), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n680), .A2(G1), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n215), .B2(new_n683), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT28), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n319), .A2(new_n316), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n279), .A2(new_n285), .A3(new_n314), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n687), .A2(KEYINPUT98), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT98), .B1(new_n687), .B2(new_n688), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n626), .B1(new_n624), .B2(new_n602), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n629), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n279), .A2(new_n636), .A3(new_n285), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n636), .B1(new_n279), .B2(new_n285), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n694), .A2(new_n695), .A3(new_n632), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n696), .A2(KEYINPUT97), .A3(KEYINPUT26), .A4(new_n569), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n634), .A2(KEYINPUT26), .A3(new_n569), .A4(new_n637), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n562), .A2(new_n568), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n635), .B1(new_n688), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(KEYINPUT97), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n654), .B1(new_n693), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT29), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n639), .A2(new_n657), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT96), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n706), .B(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n705), .B1(new_n708), .B2(KEYINPUT29), .ZN(new_n709));
  INV_X1    g0509(.A(new_n256), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n282), .A2(KEYINPUT82), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n275), .A2(new_n276), .A3(new_n254), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n548), .ZN(new_n714));
  AOI21_X1  g0514(.A(G179), .B1(new_n519), .B2(new_n525), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n579), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(KEYINPUT95), .B1(new_n713), .B2(new_n716), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n715), .A2(new_n714), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT95), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n315), .A2(new_n718), .A3(new_n719), .A4(new_n579), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n578), .A2(new_n282), .A3(new_n256), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n548), .A2(G179), .A3(new_n525), .A4(new_n519), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n723), .A2(new_n724), .A3(new_n722), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT94), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI211_X1 g0528(.A(KEYINPUT94), .B(new_n722), .C1(new_n723), .C2(new_n724), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n721), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(new_n654), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT31), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n320), .A2(new_n609), .A3(new_n535), .A4(new_n657), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n725), .B1(new_n713), .B2(new_n716), .ZN(new_n735));
  OAI211_X1 g0535(.A(KEYINPUT31), .B(new_n654), .C1(new_n735), .C2(new_n726), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT93), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n736), .A2(new_n737), .ZN(new_n739));
  OAI211_X1 g0539(.A(new_n733), .B(new_n734), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G330), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n709), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n686), .B1(new_n742), .B2(G1), .ZN(G364));
  XOR2_X1   g0543(.A(new_n670), .B(KEYINPUT99), .Z(new_n744));
  INV_X1    g0544(.A(G13), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n745), .A2(new_n537), .A3(G20), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n746), .A2(KEYINPUT100), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(KEYINPUT100), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n747), .A2(G1), .A3(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n682), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n750), .B1(new_n668), .B2(new_n669), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n744), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT101), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n213), .B1(G20), .B2(new_n284), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XOR2_X1   g0558(.A(new_n758), .B(KEYINPUT102), .Z(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT103), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n210), .A2(new_n271), .ZN(new_n761));
  INV_X1    g0561(.A(G355), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n761), .A2(new_n762), .B1(G116), .B2(new_n210), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n681), .A2(new_n271), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n765), .B1(new_n216), .B2(new_n421), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n240), .A2(new_n537), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n763), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n750), .B1(new_n760), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n317), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n207), .A2(G190), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n246), .A2(G200), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n772), .A2(new_n472), .B1(new_n775), .B2(new_n202), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n207), .A2(new_n317), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(new_n774), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT104), .Z(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n776), .B1(new_n780), .B2(G58), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT105), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n773), .A2(new_n246), .A3(G200), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT106), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G107), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n777), .A2(new_n246), .A3(G200), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n271), .B1(new_n786), .B2(new_n554), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G179), .A2(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n773), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G159), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n789), .A2(KEYINPUT32), .A3(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(KEYINPUT32), .B1(new_n789), .B2(new_n790), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n207), .B1(new_n788), .B2(G190), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n293), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n770), .A2(G190), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n795), .B1(new_n796), .B2(G68), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n785), .A2(new_n792), .A3(new_n793), .A4(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G322), .ZN(new_n799));
  INV_X1    g0599(.A(G329), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n778), .A2(new_n799), .B1(new_n789), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G311), .ZN(new_n802));
  INV_X1    g0602(.A(new_n796), .ZN(new_n803));
  XOR2_X1   g0603(.A(KEYINPUT33), .B(G317), .Z(new_n804));
  OAI221_X1 g0604(.A(new_n268), .B1(new_n775), .B2(new_n802), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n786), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n801), .B(new_n805), .C1(G303), .C2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G283), .ZN(new_n808));
  INV_X1    g0608(.A(new_n784), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n794), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n811), .A2(G294), .B1(G326), .B2(new_n771), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n812), .B(KEYINPUT107), .Z(new_n813));
  OAI22_X1  g0613(.A1(new_n782), .A2(new_n798), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n769), .B1(new_n814), .B2(new_n757), .ZN(new_n815));
  INV_X1    g0615(.A(new_n756), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n815), .B1(new_n667), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n753), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT108), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G396));
  NAND4_X1  g0620(.A1(new_n613), .A2(new_n503), .A3(new_n614), .A4(new_n654), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n654), .A2(new_n503), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n822), .A2(new_n506), .A3(new_n504), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n639), .A2(new_n824), .A3(new_n657), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n708), .B2(new_n824), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n750), .B1(new_n826), .B2(new_n741), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n741), .B2(new_n826), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n757), .A2(new_n754), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n750), .B1(G77), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n775), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n271), .B(new_n795), .C1(G116), .C2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(G294), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n786), .A2(new_n300), .B1(new_n778), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n789), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n835), .B1(G311), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n784), .A2(G87), .ZN(new_n838));
  AOI22_X1  g0638(.A1(G283), .A2(new_n796), .B1(new_n771), .B2(G303), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n833), .A2(new_n837), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n832), .A2(G159), .B1(G137), .B2(new_n771), .ZN(new_n841));
  INV_X1    g0641(.A(G143), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n841), .B1(new_n337), .B2(new_n803), .C1(new_n779), .C2(new_n842), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT34), .Z(new_n844));
  OAI21_X1  g0644(.A(new_n271), .B1(new_n786), .B2(new_n472), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(G132), .B2(new_n836), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n846), .B1(new_n328), .B2(new_n794), .C1(new_n809), .C2(new_n384), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n840), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n831), .B1(new_n848), .B2(new_n757), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n824), .B2(new_n755), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n828), .A2(new_n850), .ZN(G384));
  INV_X1    g0651(.A(new_n296), .ZN(new_n852));
  OR2_X1    g0652(.A1(new_n852), .A2(KEYINPUT35), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(KEYINPUT35), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n853), .A2(G116), .A3(new_n214), .A4(new_n854), .ZN(new_n855));
  XOR2_X1   g0655(.A(new_n855), .B(KEYINPUT36), .Z(new_n856));
  NOR3_X1   g0656(.A1(new_n385), .A2(new_n215), .A3(new_n202), .ZN(new_n857));
  OR2_X1    g0657(.A1(new_n857), .A2(KEYINPUT109), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n857), .A2(KEYINPUT109), .B1(new_n472), .B2(G68), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n206), .B(G13), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(G1), .B1(new_n745), .B2(G20), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n508), .B(new_n705), .C1(new_n708), .C2(KEYINPUT29), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n622), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n413), .A2(new_n414), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n398), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n383), .B1(new_n866), .B2(new_n397), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n430), .B1(new_n867), .B2(new_n411), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n867), .A2(new_n649), .ZN(new_n869));
  OAI21_X1  g0669(.A(KEYINPUT37), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n433), .A2(new_n410), .ZN(new_n871));
  XOR2_X1   g0671(.A(new_n649), .B(KEYINPUT111), .Z(new_n872));
  NAND2_X1  g0672(.A1(new_n433), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT37), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n871), .A2(new_n873), .A3(new_n874), .A4(new_n430), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n437), .A2(new_n869), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(new_n877), .A3(KEYINPUT38), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n871), .A2(new_n873), .A3(new_n430), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT37), .ZN(new_n880));
  INV_X1    g0680(.A(new_n873), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n880), .A2(new_n875), .B1(new_n437), .B2(new_n881), .ZN(new_n882));
  XNOR2_X1  g0682(.A(KEYINPUT112), .B(KEYINPUT38), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n878), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT39), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT110), .B1(new_n469), .B2(new_n488), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT110), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n888), .B(new_n487), .C1(new_n464), .C2(new_n468), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n876), .A2(new_n877), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT38), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(KEYINPUT39), .A3(new_n878), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n886), .A2(new_n657), .A3(new_n891), .A4(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n504), .A2(new_n654), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n825), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n894), .A2(new_n878), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n489), .A2(new_n888), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n616), .A2(KEYINPUT110), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n488), .A2(new_n654), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n903), .A2(new_n491), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n489), .A2(new_n657), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n899), .A2(new_n900), .A3(new_n908), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n619), .A2(new_n872), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n896), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n864), .B(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n729), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(new_n717), .B2(new_n720), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n657), .B1(new_n914), .B2(new_n728), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(KEYINPUT31), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n733), .A2(new_n916), .A3(new_n734), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n884), .A2(new_n908), .A3(new_n824), .A4(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n734), .B1(new_n915), .B2(KEYINPUT31), .ZN(new_n919));
  AOI211_X1 g0719(.A(new_n732), .B(new_n657), .C1(new_n914), .C2(new_n728), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n824), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n906), .B1(new_n890), .B2(new_n904), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT40), .B1(new_n894), .B2(new_n878), .ZN(new_n924));
  AOI22_X1  g0724(.A1(KEYINPUT40), .A2(new_n918), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n508), .A2(new_n917), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n669), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n927), .B2(new_n926), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n862), .B1(new_n912), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT113), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n912), .A2(new_n929), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n930), .B2(new_n931), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n861), .B1(new_n932), .B2(new_n934), .ZN(G367));
  OAI21_X1  g0735(.A(new_n691), .B1(new_n632), .B2(new_n657), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n696), .A2(new_n654), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n659), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n939), .B(KEYINPUT42), .Z(new_n940));
  INV_X1    g0740(.A(new_n938), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n688), .B1(new_n941), .B2(new_n602), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n657), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n657), .A2(new_n561), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT114), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(new_n699), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n940), .A2(new_n943), .B1(KEYINPUT43), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n946), .A2(KEYINPUT43), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n947), .B(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n676), .A2(new_n938), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n949), .B(new_n950), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n682), .B(KEYINPUT41), .Z(new_n952));
  NOR2_X1   g0752(.A1(new_n664), .A2(new_n938), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT44), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n941), .B1(new_n662), .B2(new_n663), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT45), .ZN(new_n956));
  AND3_X1   g0756(.A1(new_n954), .A2(new_n956), .A3(new_n677), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n677), .B1(new_n954), .B2(new_n956), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n675), .A2(new_n658), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n660), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n671), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(new_n744), .B2(new_n960), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n742), .A2(new_n962), .ZN(new_n963));
  OR3_X1    g0763(.A1(new_n957), .A2(new_n958), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n952), .B1(new_n964), .B2(new_n742), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n951), .B1(new_n965), .B2(new_n749), .ZN(new_n966));
  INV_X1    g0766(.A(new_n759), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n210), .B2(new_n499), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n765), .A2(new_n236), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n750), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n202), .A2(new_n783), .B1(new_n778), .B2(new_n337), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n271), .B1(new_n786), .B2(new_n328), .C1(new_n790), .C2(new_n803), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n811), .A2(G68), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n772), .B2(new_n842), .ZN(new_n974));
  INV_X1    g0774(.A(G137), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n775), .A2(new_n472), .B1(new_n789), .B2(new_n975), .ZN(new_n976));
  OR4_X1    g0776(.A1(new_n971), .A2(new_n972), .A3(new_n974), .A4(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(G317), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n783), .A2(new_n293), .B1(new_n789), .B2(new_n978), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n271), .B(new_n979), .C1(G283), .C2(new_n832), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n786), .A2(new_n514), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n981), .A2(KEYINPUT46), .B1(new_n796), .B2(G294), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n980), .B(new_n982), .C1(new_n521), .C2(new_n779), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n771), .A2(G311), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n984), .B1(new_n300), .B2(new_n794), .C1(new_n981), .C2(KEYINPUT46), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n977), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT47), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n970), .B1(new_n987), .B2(new_n757), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT115), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n946), .B2(new_n816), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n966), .A2(new_n990), .ZN(G387));
  OAI21_X1  g0791(.A(new_n764), .B1(new_n233), .B2(new_n421), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n680), .B2(new_n761), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n497), .A2(new_n472), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT50), .Z(new_n995));
  AOI21_X1  g0795(.A(G45), .B1(G68), .B2(G77), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n995), .A2(new_n680), .A3(new_n996), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n993), .A2(new_n997), .B1(new_n300), .B2(new_n681), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n750), .B1(new_n998), .B2(new_n760), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n832), .A2(G303), .B1(G311), .B2(new_n796), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(new_n799), .B2(new_n772), .C1(new_n779), .C2(new_n978), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT48), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n806), .A2(G294), .B1(new_n811), .B2(G283), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT49), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n783), .A2(new_n514), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n271), .B(new_n1010), .C1(G326), .C2(new_n836), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n806), .A2(G77), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1013), .B(new_n271), .C1(new_n790), .C2(new_n772), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n794), .A2(new_n499), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n335), .A2(new_n796), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n784), .A2(G97), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n778), .A2(new_n472), .B1(new_n775), .B2(new_n384), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(G150), .B2(new_n836), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .A4(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1012), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n999), .B1(new_n1022), .B2(new_n757), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n674), .B2(new_n816), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT116), .Z(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n962), .B2(new_n749), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n963), .A2(new_n682), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n742), .A2(new_n962), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(G393));
  OAI21_X1  g0829(.A(new_n963), .B1(new_n957), .B2(new_n958), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n964), .A2(new_n682), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n749), .ZN(new_n1032));
  NOR3_X1   g0832(.A1(new_n957), .A2(new_n958), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n941), .A2(new_n756), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n967), .B1(new_n293), .B2(new_n210), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n764), .A2(new_n244), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n750), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n794), .A2(new_n202), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n497), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n271), .B1(new_n1039), .B2(new_n775), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1038), .B(new_n1040), .C1(G50), .C2(new_n796), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n786), .A2(new_n384), .B1(new_n789), .B2(new_n842), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT117), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1041), .A2(new_n838), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n778), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n1047), .A2(G159), .B1(G150), .B2(new_n771), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT51), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n1047), .A2(G311), .B1(G317), .B2(new_n771), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT52), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n271), .B1(new_n806), .B2(G283), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G294), .A2(new_n832), .B1(new_n836), .B2(G322), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n811), .A2(G116), .B1(G303), .B2(new_n796), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n785), .A2(new_n1052), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n1046), .A2(new_n1049), .B1(new_n1051), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1037), .B1(new_n1056), .B2(new_n757), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1033), .B1(new_n1034), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1031), .A2(new_n1058), .ZN(G390));
  AND2_X1   g0859(.A1(new_n697), .A2(new_n702), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n687), .A2(new_n688), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT98), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n687), .A2(KEYINPUT98), .A3(new_n688), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n692), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n568), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n657), .B(new_n824), .C1(new_n1060), .C2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n922), .B1(new_n1067), .B2(new_n898), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n891), .A2(new_n657), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n884), .ZN(new_n1070));
  OAI21_X1  g0870(.A(KEYINPUT118), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT118), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1070), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n897), .B1(new_n704), .B2(new_n824), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1072), .B(new_n1073), .C1(new_n1074), .C2(new_n922), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1071), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n899), .A2(new_n908), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1077), .A2(new_n1069), .B1(new_n886), .B2(new_n895), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n908), .A2(new_n740), .A3(G330), .A4(new_n824), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1076), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1078), .B1(new_n1071), .B2(new_n1075), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n917), .A2(G330), .A3(new_n824), .ZN(new_n1083));
  OR3_X1    g0883(.A1(new_n1083), .A2(KEYINPUT119), .A3(new_n922), .ZN(new_n1084));
  OAI21_X1  g0884(.A(KEYINPUT119), .B1(new_n1083), .B2(new_n922), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1081), .B1(new_n1082), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n824), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n922), .B1(new_n741), .B2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1084), .A2(new_n1085), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n899), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1083), .A2(new_n922), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1092), .A2(new_n1080), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n1074), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1091), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n508), .A2(G330), .A3(new_n917), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n863), .A2(new_n622), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n683), .B1(new_n1087), .B2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1082), .A2(new_n1086), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1080), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1102), .B(new_n1078), .C1(new_n1071), .C2(new_n1075), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1090), .A2(new_n899), .B1(new_n1074), .B2(new_n1093), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1105), .A2(new_n1097), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1100), .A2(new_n1107), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n772), .A2(new_n808), .B1(new_n202), .B2(new_n794), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(G116), .A2(new_n1047), .B1(new_n832), .B2(G97), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n1110), .B1(new_n834), .B2(new_n789), .C1(new_n809), .C2(new_n384), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1109), .B(new_n1111), .C1(G107), .C2(new_n796), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n271), .B1(new_n806), .B2(G87), .ZN(new_n1113));
  XOR2_X1   g0913(.A(new_n1113), .B(KEYINPUT120), .Z(new_n1114));
  NOR2_X1   g0914(.A1(new_n794), .A2(new_n790), .ZN(new_n1115));
  INV_X1    g0915(.A(G132), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n271), .B1(new_n778), .B2(new_n1116), .C1(new_n975), .C2(new_n803), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1115), .B(new_n1117), .C1(G128), .C2(new_n771), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n836), .A2(G125), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(KEYINPUT54), .B(G143), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1119), .B1(new_n472), .B2(new_n783), .C1(new_n775), .C2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT53), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n786), .B2(new_n337), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n806), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1121), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n1112), .A2(new_n1114), .B1(new_n1118), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n757), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n750), .B1(new_n335), .B2(new_n830), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n886), .A2(new_n895), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1128), .B1(new_n1129), .B2(new_n754), .ZN(new_n1130));
  OR2_X1    g0930(.A1(new_n1130), .A2(KEYINPUT121), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(KEYINPUT121), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1104), .A2(new_n749), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1108), .A2(new_n1133), .ZN(G378));
  OAI21_X1  g0934(.A(new_n750), .B1(G50), .B2(new_n830), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n649), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n340), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n376), .A2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n371), .A2(new_n372), .A3(new_n375), .A4(new_n1137), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1139), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1146), .A2(new_n755), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n803), .A2(new_n1116), .B1(new_n794), .B2(new_n337), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1120), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n806), .A2(new_n1149), .B1(new_n1047), .B2(G128), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n975), .B2(new_n775), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1148), .B(new_n1151), .C1(G125), .C2(new_n771), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  OR2_X1    g0953(.A1(new_n1153), .A2(KEYINPUT59), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(KEYINPUT59), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n257), .B(new_n422), .C1(new_n783), .C2(new_n790), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(G124), .B2(new_n836), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1154), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n271), .A2(G41), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(G97), .A2(new_n796), .B1(new_n771), .B2(G116), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1013), .A2(new_n973), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n783), .A2(new_n328), .B1(new_n775), .B2(new_n499), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n778), .A2(new_n300), .B1(new_n789), .B2(new_n808), .ZN(new_n1163));
  NOR3_X1   g0963(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(KEYINPUT58), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1159), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1166), .B(new_n472), .C1(G33), .C2(G41), .ZN(new_n1167));
  OR2_X1    g0967(.A1(new_n1164), .A2(KEYINPUT58), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1158), .A2(new_n1165), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1135), .B(new_n1147), .C1(new_n757), .C2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(KEYINPUT122), .B1(new_n925), .B2(new_n669), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1146), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT122), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT40), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n923), .B2(new_n884), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n900), .A2(new_n1174), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n908), .A2(new_n824), .A3(new_n917), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1173), .B(G330), .C1(new_n1175), .C2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1171), .A2(new_n1172), .A3(new_n1179), .ZN(new_n1180));
  OAI211_X1 g0980(.A(G330), .B(new_n1146), .C1(new_n1175), .C2(new_n1178), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n911), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n918), .A2(KEYINPUT40), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n923), .A2(new_n924), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n669), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n911), .B1(new_n1186), .B2(new_n1146), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT123), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n1180), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1188), .B1(new_n1180), .B2(new_n1187), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1183), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1170), .B1(new_n1191), .B2(new_n749), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1098), .B1(new_n1087), .B2(new_n1099), .ZN(new_n1193));
  AOI21_X1  g0993(.A(KEYINPUT57), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1097), .B1(new_n1104), .B2(new_n1095), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n896), .A2(new_n909), .A3(new_n910), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1181), .A2(new_n1196), .ZN(new_n1198));
  OAI21_X1  g0998(.A(G330), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1146), .B1(new_n1199), .B2(KEYINPUT122), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1198), .B1(new_n1200), .B2(new_n1179), .ZN(new_n1201));
  OAI21_X1  g1001(.A(KEYINPUT57), .B1(new_n1197), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n682), .B1(new_n1195), .B2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1192), .B1(new_n1194), .B2(new_n1203), .ZN(G375));
  AOI211_X1 g1004(.A(new_n749), .B(new_n682), .C1(new_n384), .C2(new_n829), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n803), .A2(new_n514), .B1(new_n772), .B2(new_n834), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n268), .B1(new_n789), .B2(new_n521), .ZN(new_n1207));
  NOR3_X1   g1007(.A1(new_n1206), .A2(new_n1015), .A3(new_n1207), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(G283), .A2(new_n1047), .B1(new_n832), .B2(G107), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n293), .B2(new_n786), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G77), .B2(new_n784), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(G150), .A2(new_n832), .B1(new_n836), .B2(G128), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n790), .B2(new_n786), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G137), .B2(new_n780), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n271), .B1(new_n783), .B2(new_n328), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n772), .A2(new_n1116), .B1(new_n794), .B2(new_n472), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(new_n796), .C2(new_n1149), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n1208), .A2(new_n1211), .B1(new_n1214), .B2(new_n1217), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1205), .B1(new_n1127), .B2(new_n1218), .C1(new_n908), .C2(new_n755), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(new_n1105), .B2(new_n1032), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1106), .A2(new_n952), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1105), .A2(new_n1097), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1220), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(G381));
  INV_X1    g1024(.A(G387), .ZN(new_n1225));
  NOR4_X1   g1025(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1225), .A2(new_n1226), .A3(new_n1223), .ZN(new_n1227));
  OR3_X1    g1027(.A1(new_n1227), .A2(G378), .A3(G375), .ZN(G407));
  AND2_X1   g1028(.A1(new_n1108), .A2(new_n1133), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n650), .A2(G213), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1232));
  OAI211_X1 g1032(.A(G407), .B(G213), .C1(G375), .C2(new_n1232), .ZN(G409));
  XNOR2_X1  g1033(.A(new_n819), .B(G393), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n1234), .A2(G390), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(G390), .A2(new_n1234), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(G387), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1225), .A2(new_n1236), .A3(new_n1235), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1240), .A2(KEYINPUT61), .ZN(new_n1241));
  OAI211_X1 g1041(.A(G378), .B(new_n1192), .C1(new_n1194), .C2(new_n1203), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n952), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1191), .A2(new_n1243), .A3(new_n1193), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1180), .A2(new_n1187), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1183), .A2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1170), .B1(new_n1246), .B2(new_n749), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1244), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1229), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1242), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT124), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1242), .A2(new_n1249), .A3(KEYINPUT124), .ZN(new_n1253));
  INV_X1    g1053(.A(G384), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1091), .A2(new_n1097), .A3(KEYINPUT60), .A4(new_n1094), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n682), .ZN(new_n1256));
  OAI21_X1  g1056(.A(KEYINPUT60), .B1(new_n1105), .B2(new_n1097), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1256), .B1(new_n1222), .B2(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1254), .B1(new_n1258), .B2(new_n1220), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1220), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1257), .A2(new_n1222), .ZN(new_n1261));
  OAI211_X1 g1061(.A(G384), .B(new_n1260), .C1(new_n1261), .C2(new_n1256), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1259), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1252), .A2(new_n1230), .A3(new_n1253), .A4(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT63), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1252), .A2(new_n1230), .A3(new_n1253), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1231), .A2(G2897), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n1263), .B2(KEYINPUT125), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT125), .ZN(new_n1271));
  AND3_X1   g1071(.A1(new_n1259), .A2(new_n1271), .A3(new_n1262), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1271), .B1(new_n1259), .B2(new_n1262), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1268), .B(new_n1270), .C1(new_n1269), .C2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1231), .B1(new_n1242), .B2(new_n1249), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(KEYINPUT63), .A3(new_n1264), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1241), .A2(new_n1267), .A3(new_n1275), .A4(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT61), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1270), .B1(new_n1274), .B2(new_n1269), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1279), .B1(new_n1280), .B2(new_n1276), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT62), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1265), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1276), .A2(KEYINPUT62), .A3(new_n1264), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1281), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT126), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1240), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  AOI211_X1 g1087(.A(KEYINPUT126), .B(new_n1281), .C1(new_n1283), .C2(new_n1284), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1278), .B1(new_n1287), .B2(new_n1288), .ZN(G405));
  NAND2_X1  g1089(.A1(G375), .A2(new_n1229), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1290), .B(new_n1264), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1242), .A2(KEYINPUT127), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1291), .B(new_n1292), .ZN(new_n1293));
  XNOR2_X1  g1093(.A(new_n1293), .B(new_n1240), .ZN(G402));
endmodule


