//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 1 1 1 1 0 1 0 0 0 1 0 0 0 0 1 0 0 1 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1209, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT0), .Z(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G107), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n217), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G50), .ZN(new_n219));
  INV_X1    g0019(.A(G226), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G58), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n208), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT65), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT1), .Z(new_n229));
  AND3_X1   g0029(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n230));
  AOI21_X1  g0030(.A(KEYINPUT64), .B1(G1), .B2(G13), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n232), .A2(new_n206), .ZN(new_n233));
  NOR2_X1   g0033(.A1(G58), .A2(G68), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n235), .A2(G50), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(new_n237));
  AOI211_X1 g0037(.A(new_n211), .B(new_n229), .C1(new_n233), .C2(new_n237), .ZN(G361));
  XOR2_X1   g0038(.A(G238), .B(G244), .Z(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G226), .B(G232), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n216), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G270), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G358));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G87), .B(G116), .Z(new_n251));
  XNOR2_X1  g0051(.A(G97), .B(G107), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  NAND2_X1  g0054(.A1(new_n225), .A2(G1698), .ZN(new_n255));
  AND2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  OAI221_X1 g0057(.A(new_n255), .B1(G226), .B2(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT72), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G97), .ZN(new_n260));
  AND3_X1   g0060(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n259), .B1(new_n258), .B2(new_n260), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  OAI22_X1  g0064(.A1(new_n230), .A2(new_n231), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NOR3_X1   g0065(.A1(new_n261), .A2(new_n262), .A3(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G274), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  AOI211_X1 g0068(.A(G1), .B(new_n267), .C1(new_n264), .C2(new_n268), .ZN(new_n269));
  AND2_X1   g0069(.A1(KEYINPUT67), .A2(G1), .ZN(new_n270));
  NOR2_X1   g0070(.A1(KEYINPUT67), .A2(G1), .ZN(new_n271));
  OAI22_X1  g0071(.A1(new_n270), .A2(new_n271), .B1(G41), .B2(G45), .ZN(new_n272));
  OAI211_X1 g0072(.A(G1), .B(G13), .C1(new_n263), .C2(new_n264), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n269), .B1(new_n274), .B2(G238), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(KEYINPUT13), .B1(new_n266), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n262), .ZN(new_n278));
  INV_X1    g0078(.A(new_n265), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT13), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(new_n282), .A3(new_n275), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT73), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n277), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  OAI211_X1 g0085(.A(KEYINPUT73), .B(KEYINPUT13), .C1(new_n266), .C2(new_n276), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(G200), .A3(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n263), .A2(G20), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n288), .A2(G77), .B1(G20), .B2(new_n213), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n289), .B1(new_n219), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n232), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT11), .ZN(new_n296));
  OR2_X1    g0096(.A1(KEYINPUT67), .A2(G1), .ZN(new_n297));
  NAND2_X1  g0097(.A1(KEYINPUT67), .A2(G1), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n294), .B1(G20), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n296), .B1(new_n213), .B2(new_n301), .ZN(new_n302));
  OAI211_X1 g0102(.A(G13), .B(G20), .C1(new_n270), .C2(new_n271), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT74), .B1(new_n303), .B2(G68), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n304), .B(KEYINPUT12), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n277), .A2(new_n283), .A3(G190), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n287), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n285), .A2(G169), .A3(new_n286), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT14), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT14), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n285), .A2(new_n312), .A3(G169), .A4(new_n286), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n277), .A2(new_n283), .A3(G179), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n311), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n306), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n309), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n300), .A2(G50), .ZN(new_n318));
  INV_X1    g0118(.A(G150), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n291), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n206), .B1(new_n234), .B2(new_n219), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n224), .A2(KEYINPUT8), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT69), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT69), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n324), .B(KEYINPUT8), .C1(new_n224), .C2(KEYINPUT70), .ZN(new_n325));
  OR2_X1    g0125(.A1(new_n224), .A2(KEYINPUT8), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n323), .B(new_n325), .C1(new_n326), .C2(KEYINPUT70), .ZN(new_n327));
  AOI211_X1 g0127(.A(new_n320), .B(new_n321), .C1(new_n327), .C2(new_n288), .ZN(new_n328));
  INV_X1    g0128(.A(new_n231), .ZN(new_n329));
  NAND3_X1  g0129(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n330));
  AND3_X1   g0130(.A1(new_n329), .A2(new_n330), .A3(new_n293), .ZN(new_n331));
  OAI221_X1 g0131(.A(new_n318), .B1(G50), .B2(new_n303), .C1(new_n328), .C2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT9), .ZN(new_n333));
  OR2_X1    g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT3), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n263), .ZN(new_n336));
  NAND2_X1  g0136(.A1(KEYINPUT3), .A2(G33), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G1698), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G222), .ZN(new_n340));
  INV_X1    g0140(.A(G223), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n338), .B(new_n340), .C1(new_n341), .C2(new_n339), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(G77), .B2(new_n338), .ZN(new_n343));
  OR2_X1    g0143(.A1(new_n343), .A2(KEYINPUT68), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(KEYINPUT68), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n344), .A2(new_n279), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n269), .B1(new_n274), .B2(G226), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G200), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n332), .A2(new_n333), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n346), .A2(G190), .A3(new_n347), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n334), .A2(new_n349), .A3(new_n350), .A4(new_n351), .ZN(new_n352));
  OR2_X1    g0152(.A1(new_n352), .A2(KEYINPUT10), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(KEYINPUT10), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n256), .A2(new_n257), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n356), .B1(G238), .B2(G1698), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n225), .B2(G1698), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n358), .B(new_n279), .C1(G107), .C2(new_n338), .ZN(new_n359));
  INV_X1    g0159(.A(new_n269), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n272), .A2(new_n273), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n359), .B(new_n360), .C1(new_n222), .C2(new_n361), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n362), .A2(G200), .ZN(new_n363));
  INV_X1    g0163(.A(G190), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n300), .A2(G77), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n326), .A2(new_n322), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n367), .A2(new_n291), .B1(new_n206), .B2(new_n221), .ZN(new_n368));
  XOR2_X1   g0168(.A(KEYINPUT15), .B(G87), .Z(new_n369));
  AOI21_X1  g0169(.A(new_n368), .B1(new_n369), .B2(new_n288), .ZN(new_n370));
  OAI221_X1 g0170(.A(new_n366), .B1(G77), .B2(new_n303), .C1(new_n370), .C2(new_n331), .ZN(new_n371));
  OR3_X1    g0171(.A1(new_n363), .A2(new_n365), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n317), .A2(new_n355), .A3(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G169), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n348), .A2(new_n374), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n375), .B(new_n332), .C1(G179), .C2(new_n348), .ZN(new_n376));
  XNOR2_X1  g0176(.A(new_n376), .B(KEYINPUT71), .ZN(new_n377));
  OR2_X1    g0177(.A1(new_n362), .A2(G179), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n362), .A2(new_n374), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(new_n371), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(G250), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n382), .B1(new_n336), .B2(new_n337), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT78), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n384), .A2(KEYINPUT4), .ZN(new_n385));
  OAI21_X1  g0185(.A(G1698), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G283), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n263), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(G244), .B1(new_n256), .B2(new_n257), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n388), .B1(new_n389), .B2(new_n385), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT4), .ZN(new_n392));
  OAI211_X1 g0192(.A(G244), .B(new_n339), .C1(new_n256), .C2(new_n257), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n392), .B1(new_n393), .B2(KEYINPUT78), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n279), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  XOR2_X1   g0195(.A(KEYINPUT5), .B(G41), .Z(new_n396));
  OAI21_X1  g0196(.A(G45), .B1(new_n270), .B2(new_n271), .ZN(new_n397));
  OAI211_X1 g0197(.A(G257), .B(new_n273), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n268), .B1(new_n297), .B2(new_n298), .ZN(new_n399));
  XNOR2_X1  g0199(.A(KEYINPUT5), .B(G41), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n399), .A2(G274), .A3(new_n273), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n395), .A2(G179), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n222), .B1(new_n336), .B2(new_n337), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n384), .B1(new_n405), .B2(new_n339), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n386), .B(new_n390), .C1(new_n406), .C2(new_n392), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n402), .B1(new_n407), .B2(new_n279), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n404), .B1(new_n374), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT7), .B1(new_n356), .B2(new_n206), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT7), .ZN(new_n411));
  NOR4_X1   g0211(.A1(new_n256), .A2(new_n257), .A3(new_n411), .A4(G20), .ZN(new_n412));
  OAI21_X1  g0212(.A(G107), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT6), .ZN(new_n414));
  INV_X1    g0214(.A(G97), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n415), .A2(new_n215), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n414), .B1(new_n416), .B2(new_n202), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n215), .A2(KEYINPUT6), .A3(G97), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G20), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n290), .A2(G77), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n413), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n294), .ZN(new_n423));
  OAI21_X1  g0223(.A(G33), .B1(new_n270), .B2(new_n271), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n303), .A2(new_n232), .A3(new_n424), .A4(new_n293), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT77), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n331), .A2(KEYINPUT77), .A3(new_n303), .A4(new_n424), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(new_n428), .A3(G97), .ZN(new_n429));
  INV_X1    g0229(.A(new_n303), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n415), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n423), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n409), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n385), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n405), .A2(new_n434), .B1(new_n263), .B2(new_n387), .ZN(new_n435));
  OAI21_X1  g0235(.A(G250), .B1(new_n256), .B2(new_n257), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n339), .B1(new_n436), .B2(new_n434), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n394), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n265), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(G200), .B1(new_n440), .B2(new_n402), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n408), .A2(G190), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n422), .A2(new_n294), .B1(new_n415), .B2(new_n430), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n441), .A2(new_n442), .A3(new_n429), .A4(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n382), .A2(new_n339), .ZN(new_n445));
  OAI221_X1 g0245(.A(new_n445), .B1(G257), .B2(new_n339), .C1(new_n256), .C2(new_n257), .ZN(new_n446));
  INV_X1    g0246(.A(G294), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n446), .B1(new_n263), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n279), .ZN(new_n449));
  OAI211_X1 g0249(.A(G264), .B(new_n273), .C1(new_n396), .C2(new_n397), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n449), .A2(KEYINPUT86), .A3(new_n401), .A4(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(G257), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n336), .A2(new_n337), .B1(new_n452), .B2(G1698), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n453), .A2(new_n445), .B1(G33), .B2(G294), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n401), .B(new_n450), .C1(new_n454), .C2(new_n265), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT86), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n451), .A2(new_n457), .A3(new_n364), .ZN(new_n458));
  INV_X1    g0258(.A(G200), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n206), .A2(G33), .A3(G116), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n206), .A2(G107), .ZN(new_n463));
  XNOR2_X1  g0263(.A(new_n463), .B(KEYINPUT23), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n206), .B(G87), .C1(new_n256), .C2(new_n257), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n465), .A2(KEYINPUT22), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n465), .A2(KEYINPUT22), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n462), .B(new_n464), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT24), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g0270(.A(new_n465), .B(KEYINPUT22), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n471), .A2(KEYINPUT24), .A3(new_n462), .A4(new_n464), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n470), .A2(new_n294), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT25), .ZN(new_n474));
  OR2_X1    g0274(.A1(new_n474), .A2(KEYINPUT84), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(KEYINPUT84), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n430), .A2(new_n215), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT85), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n475), .B(new_n476), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(new_n478), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n477), .A2(new_n478), .A3(new_n475), .A4(new_n476), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n427), .A2(new_n428), .A3(G107), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n473), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n433), .B(new_n444), .C1(new_n461), .C2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n303), .A2(new_n369), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n338), .A2(new_n206), .A3(G68), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n288), .A2(G97), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT19), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g0291(.A(KEYINPUT79), .B(G87), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n492), .A2(new_n203), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n260), .A2(new_n490), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n494), .A2(G20), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n488), .B(new_n491), .C1(new_n493), .C2(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n487), .B1(new_n496), .B2(new_n294), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n427), .A2(new_n428), .A3(G87), .ZN(new_n498));
  AND2_X1   g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n214), .A2(new_n339), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n222), .A2(G1698), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n500), .B(new_n501), .C1(new_n256), .C2(new_n257), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G33), .A2(G116), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n279), .ZN(new_n505));
  OAI211_X1 g0305(.A(G45), .B(new_n267), .C1(new_n270), .C2(new_n271), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n506), .B(new_n273), .C1(new_n399), .C2(G250), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n505), .A2(new_n364), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n505), .A2(new_n507), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n508), .B1(new_n510), .B2(G200), .ZN(new_n511));
  INV_X1    g0311(.A(G179), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n505), .A2(new_n512), .A3(new_n507), .ZN(new_n513));
  AOI21_X1  g0313(.A(G169), .B1(new_n505), .B2(new_n507), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n427), .A2(new_n428), .A3(new_n369), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n497), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n499), .A2(new_n511), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n486), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n339), .A2(G257), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n338), .B(new_n521), .C1(new_n216), .C2(new_n339), .ZN(new_n522));
  XOR2_X1   g0322(.A(KEYINPUT81), .B(G303), .Z(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n356), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n279), .A3(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(G270), .B(new_n273), .C1(new_n396), .C2(new_n397), .ZN(new_n526));
  AND3_X1   g0326(.A1(new_n526), .A2(KEYINPUT80), .A3(new_n401), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT80), .B1(new_n526), .B2(new_n401), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(KEYINPUT82), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT82), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n531), .B(new_n525), .C1(new_n527), .C2(new_n528), .ZN(new_n532));
  AND2_X1   g0332(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(G200), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n303), .A2(G116), .ZN(new_n535));
  INV_X1    g0335(.A(G116), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G20), .ZN(new_n537));
  AOI21_X1  g0337(.A(G20), .B1(G33), .B2(G283), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n263), .A2(G97), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT83), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n540), .B1(new_n538), .B2(new_n539), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n294), .B(new_n537), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT20), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n543), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n541), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n548), .A2(KEYINPUT20), .A3(new_n294), .A4(new_n537), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n535), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  OR2_X1    g0350(.A1(new_n425), .A2(new_n536), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n534), .B(new_n553), .C1(new_n364), .C2(new_n533), .ZN(new_n554));
  NOR3_X1   g0354(.A1(new_n553), .A2(new_n512), .A3(new_n529), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n374), .B1(new_n550), .B2(new_n551), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n556), .A2(new_n530), .A3(new_n532), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT21), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT21), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n556), .A2(new_n559), .A3(new_n530), .A4(new_n532), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n555), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n374), .B1(new_n451), .B2(new_n457), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n455), .A2(new_n512), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n485), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n520), .A2(new_n554), .A3(new_n561), .A4(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT16), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n411), .B1(new_n338), .B2(G20), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n356), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n213), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G58), .A2(G68), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT75), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(KEYINPUT75), .A2(G58), .A3(G68), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n235), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(G20), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n290), .A2(G159), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n566), .B1(new_n569), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(G68), .B1(new_n410), .B2(new_n412), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n574), .A2(G20), .B1(G159), .B2(new_n290), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n579), .A2(new_n580), .A3(KEYINPUT16), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n578), .A2(new_n294), .A3(new_n581), .ZN(new_n582));
  OR2_X1    g0382(.A1(new_n327), .A2(new_n303), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n300), .A2(new_n327), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n269), .B1(new_n274), .B2(G232), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n220), .A2(G1698), .ZN(new_n587));
  OAI221_X1 g0387(.A(new_n587), .B1(G223), .B2(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n588));
  NAND2_X1  g0388(.A1(G33), .A2(G87), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n279), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT76), .B1(new_n586), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n360), .B1(new_n361), .B2(new_n225), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n265), .B1(new_n588), .B2(new_n589), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT76), .ZN(new_n595));
  NOR3_X1   g0395(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n459), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n593), .A2(new_n594), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n364), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n585), .A2(new_n600), .A3(KEYINPUT17), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT17), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n586), .A2(KEYINPUT76), .A3(new_n591), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n595), .B1(new_n593), .B2(new_n594), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n605), .A2(new_n459), .B1(new_n364), .B2(new_n598), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n602), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n601), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n605), .A2(new_n374), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n598), .A2(new_n512), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n607), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT18), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n607), .A2(KEYINPUT18), .A3(new_n610), .A4(new_n611), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n609), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NOR4_X1   g0417(.A1(new_n373), .A2(new_n381), .A3(new_n565), .A4(new_n617), .ZN(G372));
  INV_X1    g0418(.A(new_n377), .ZN(new_n619));
  INV_X1    g0419(.A(new_n380), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n315), .A2(new_n316), .B1(new_n620), .B2(new_n308), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n621), .A2(new_n609), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n614), .A2(new_n615), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT88), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT88), .B1(new_n614), .B2(new_n615), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n622), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT89), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n353), .A2(new_n354), .A3(KEYINPUT90), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT90), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n355), .A2(new_n631), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n628), .A2(new_n629), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT89), .B1(new_n622), .B2(new_n627), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n619), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n373), .A2(new_n381), .A3(new_n617), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n458), .A2(new_n460), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n637), .A2(new_n484), .A3(new_n473), .A4(new_n483), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n638), .A2(new_n518), .A3(new_n433), .A4(new_n444), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n639), .B1(new_n561), .B2(new_n564), .ZN(new_n640));
  OAI21_X1  g0440(.A(G169), .B1(new_n440), .B2(new_n402), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n641), .A2(new_n404), .B1(new_n443), .B2(new_n429), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n642), .A2(new_n518), .A3(KEYINPUT26), .ZN(new_n643));
  AOI211_X1 g0443(.A(KEYINPUT87), .B(KEYINPUT26), .C1(new_n642), .C2(new_n518), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT87), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n515), .A2(new_n517), .ZN(new_n646));
  INV_X1    g0446(.A(new_n508), .ZN(new_n647));
  AOI21_X1  g0447(.A(G200), .B1(new_n505), .B2(new_n507), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n497), .B(new_n498), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n409), .A2(new_n646), .A3(new_n649), .A4(new_n432), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT26), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n645), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n643), .B1(new_n644), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n646), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n636), .B1(new_n640), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n635), .A2(new_n655), .ZN(G369));
  NAND2_X1  g0456(.A1(new_n558), .A2(new_n560), .ZN(new_n657));
  INV_X1    g0457(.A(new_n555), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(G13), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n660), .A2(G20), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n299), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT27), .ZN(new_n663));
  OR3_X1    g0463(.A1(new_n662), .A2(KEYINPUT91), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(G213), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n665), .B1(new_n662), .B2(new_n663), .ZN(new_n666));
  OAI21_X1  g0466(.A(KEYINPUT91), .B1(new_n662), .B2(new_n663), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n664), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n668), .A2(G343), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n659), .B1(new_n553), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n561), .A2(new_n552), .A3(new_n669), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n671), .A2(new_n554), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(G330), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n564), .A2(new_n669), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n485), .A2(new_n669), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n638), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n675), .B1(new_n677), .B2(new_n564), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT92), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n561), .B2(new_n669), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n659), .A2(KEYINPUT92), .A3(new_n670), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n679), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(new_n675), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n681), .A2(new_n686), .ZN(G399));
  INV_X1    g0487(.A(new_n209), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G41), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n493), .A2(new_n536), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n690), .A2(G1), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n236), .B2(new_n690), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT28), .ZN(new_n695));
  INV_X1    g0495(.A(G330), .ZN(new_n696));
  OAI21_X1  g0496(.A(KEYINPUT31), .B1(new_n565), .B2(new_n669), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n449), .A2(new_n450), .ZN(new_n698));
  NOR3_X1   g0498(.A1(new_n529), .A2(new_n698), .A3(new_n509), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n699), .A2(KEYINPUT30), .A3(G179), .A4(new_n408), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT94), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n699), .A2(G179), .A3(new_n408), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT30), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n408), .A2(G179), .A3(new_n510), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n533), .A2(new_n455), .A3(new_n706), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n670), .B1(new_n702), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n697), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n708), .A2(KEYINPUT93), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n702), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n708), .A2(KEYINPUT93), .ZN(new_n714));
  OAI211_X1 g0514(.A(KEYINPUT31), .B(new_n669), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n696), .B1(new_n711), .B2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT29), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n561), .A2(new_n564), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT95), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n486), .B1(new_n499), .B2(new_n511), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n561), .A2(KEYINPUT95), .A3(new_n564), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n650), .A2(new_n651), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n643), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n723), .A2(new_n646), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n717), .B1(new_n726), .B2(new_n670), .ZN(new_n727));
  INV_X1    g0527(.A(new_n654), .ZN(new_n728));
  INV_X1    g0528(.A(new_n640), .ZN(new_n729));
  AOI211_X1 g0529(.A(KEYINPUT29), .B(new_n669), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n716), .A2(new_n727), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n695), .B1(new_n731), .B2(G1), .ZN(G364));
  NAND2_X1  g0532(.A1(new_n661), .A2(G45), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n690), .A2(G1), .A3(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n674), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n673), .A2(G330), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(G13), .A2(G33), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n673), .A2(G20), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n232), .B1(G20), .B2(new_n374), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n206), .A2(new_n364), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n512), .A2(G200), .ZN(new_n744));
  AND3_X1   g0544(.A1(new_n743), .A2(KEYINPUT96), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(KEYINPUT96), .B1(new_n743), .B2(new_n744), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(G322), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n206), .A2(G190), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G179), .A2(G200), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G329), .ZN(new_n754));
  NAND3_X1  g0554(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n364), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n756), .B(KEYINPUT97), .Z(new_n757));
  AOI21_X1  g0557(.A(new_n206), .B1(new_n751), .B2(G190), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n757), .A2(G326), .B1(G294), .B2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT98), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n754), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n459), .A2(G179), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n743), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n749), .B(new_n762), .C1(G303), .C2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n755), .A2(G190), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G317), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n769), .A2(KEYINPUT33), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(KEYINPUT33), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n768), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n338), .B(new_n772), .C1(new_n760), .C2(new_n761), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n766), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n750), .A2(new_n763), .ZN(new_n775));
  INV_X1    g0575(.A(G311), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n750), .A2(new_n744), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n774), .B1(new_n387), .B2(new_n775), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n756), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n779), .A2(new_n219), .B1(new_n758), .B2(new_n415), .ZN(new_n780));
  INV_X1    g0580(.A(new_n747), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n356), .B1(new_n781), .B2(G58), .ZN(new_n782));
  INV_X1    g0582(.A(G159), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n752), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT32), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n782), .B(new_n785), .C1(new_n215), .C2(new_n775), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n780), .B(new_n786), .C1(new_n492), .C2(new_n765), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n787), .B1(new_n213), .B2(new_n768), .C1(new_n221), .C2(new_n777), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n742), .B1(new_n778), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n739), .A2(G20), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n741), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n688), .A2(new_n338), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n793), .B1(new_n268), .B2(new_n237), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(new_n250), .B2(new_n268), .ZN(new_n795));
  INV_X1    g0595(.A(G355), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n209), .A2(new_n338), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n795), .B1(G116), .B2(new_n209), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n740), .B(new_n789), .C1(new_n791), .C2(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n737), .B1(new_n799), .B2(new_n734), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT99), .Z(G396));
  OAI21_X1  g0601(.A(new_n670), .B1(new_n654), .B2(new_n640), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n380), .A2(new_n669), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n669), .A2(new_n371), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n372), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n803), .B1(new_n805), .B2(new_n380), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n802), .B(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n716), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n808), .B1(new_n809), .B2(KEYINPUT100), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(KEYINPUT100), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n809), .A2(KEYINPUT100), .A3(new_n808), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n812), .A2(new_n734), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n807), .A2(new_n738), .ZN(new_n815));
  INV_X1    g0615(.A(new_n734), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n741), .A2(new_n738), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n221), .ZN(new_n818));
  INV_X1    g0618(.A(G132), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n338), .B1(new_n752), .B2(new_n819), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n767), .A2(G150), .B1(new_n756), .B2(G137), .ZN(new_n821));
  INV_X1    g0621(.A(G143), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n821), .B1(new_n783), .B2(new_n777), .C1(new_n747), .C2(new_n822), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT34), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n824), .B1(new_n219), .B2(new_n764), .C1(new_n213), .C2(new_n775), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n820), .B(new_n825), .C1(G58), .C2(new_n759), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n758), .A2(new_n415), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n338), .B(new_n827), .C1(G283), .C2(new_n767), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n781), .A2(G294), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n765), .A2(G107), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n777), .A2(new_n536), .B1(new_n752), .B2(new_n776), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(G303), .B2(new_n756), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n828), .A2(new_n829), .A3(new_n830), .A4(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n775), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n833), .B1(G87), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n741), .B1(new_n826), .B2(new_n835), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n815), .A2(new_n816), .A3(new_n818), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n814), .A2(new_n837), .ZN(G384));
  NAND2_X1  g0638(.A1(new_n585), .A2(new_n600), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n607), .A2(new_n668), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n839), .A2(new_n612), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(KEYINPUT37), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT37), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n839), .A2(new_n843), .A3(new_n612), .A4(new_n840), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n845), .B(KEYINPUT38), .C1(new_n616), .C2(new_n840), .ZN(new_n846));
  INV_X1    g0646(.A(new_n845), .ZN(new_n847));
  OR2_X1    g0647(.A1(new_n609), .A2(KEYINPUT103), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n609), .A2(KEYINPUT103), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n848), .B(new_n849), .C1(new_n625), .C2(new_n626), .ZN(new_n850));
  INV_X1    g0650(.A(new_n840), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n847), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n846), .B1(new_n852), .B2(KEYINPUT38), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT39), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n315), .A2(new_n316), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n670), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT102), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n845), .B1(new_n616), .B2(new_n840), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT38), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n846), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n855), .A2(new_n858), .A3(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n627), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n866), .A2(new_n668), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n316), .A2(new_n669), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n856), .A2(new_n669), .B1(new_n317), .B2(new_n868), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n670), .B(new_n806), .C1(new_n654), .C2(new_n640), .ZN(new_n870));
  INV_X1    g0670(.A(new_n803), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI211_X1 g0672(.A(KEYINPUT101), .B(new_n867), .C1(new_n872), .C2(new_n862), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT101), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n870), .A2(new_n871), .ZN(new_n875));
  INV_X1    g0675(.A(new_n869), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n875), .A2(new_n876), .A3(new_n862), .ZN(new_n877));
  INV_X1    g0677(.A(new_n867), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n874), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n865), .B1(new_n873), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n636), .B1(new_n727), .B2(new_n730), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n635), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n880), .B(new_n882), .Z(new_n883));
  INV_X1    g0683(.A(KEYINPUT31), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n884), .B(new_n670), .C1(new_n702), .C2(new_n708), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(new_n697), .B2(new_n710), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n886), .A2(new_n807), .A3(new_n869), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n853), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n863), .A2(KEYINPUT40), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n888), .A2(KEYINPUT40), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n886), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n636), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n696), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n890), .B2(new_n892), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n883), .B(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(new_n299), .B2(new_n661), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n536), .B1(new_n419), .B2(KEYINPUT35), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n897), .B(new_n233), .C1(KEYINPUT35), .C2(new_n419), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n898), .B(KEYINPUT36), .ZN(new_n899));
  AND4_X1   g0699(.A1(G77), .A2(new_n237), .A3(new_n572), .A4(new_n573), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n213), .A2(G50), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n660), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n896), .B(new_n899), .C1(new_n299), .C2(new_n902), .ZN(G367));
  NAND2_X1  g0703(.A1(new_n669), .A2(new_n432), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n904), .A2(new_n433), .A3(new_n444), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n642), .A2(new_n669), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n685), .B2(new_n675), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n909), .B(KEYINPUT44), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT45), .B1(new_n686), .B2(new_n907), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT45), .ZN(new_n913));
  NOR4_X1   g0713(.A1(new_n685), .A2(new_n913), .A3(new_n675), .A4(new_n908), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n911), .A2(new_n916), .A3(new_n681), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n680), .B1(new_n910), .B2(new_n915), .ZN(new_n918));
  INV_X1    g0718(.A(new_n685), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n679), .A2(new_n684), .A3(new_n683), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(new_n735), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n917), .A2(new_n918), .A3(new_n731), .A4(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n731), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n689), .B(KEYINPUT41), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT105), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT105), .ZN(new_n928));
  INV_X1    g0728(.A(new_n925), .ZN(new_n929));
  AOI211_X1 g0729(.A(new_n928), .B(new_n929), .C1(new_n923), .C2(new_n731), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n733), .A2(G1), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n927), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  OR3_X1    g0734(.A1(new_n670), .A2(new_n646), .A3(new_n499), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n518), .B1(new_n670), .B2(new_n499), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n685), .A2(new_n907), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n940), .B(KEYINPUT42), .Z(new_n941));
  OAI21_X1  g0741(.A(new_n433), .B1(new_n905), .B2(new_n564), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n670), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n939), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n681), .A2(new_n908), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT104), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n944), .A2(new_n939), .A3(new_n945), .ZN(new_n950));
  AND3_X1   g0750(.A1(new_n947), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n949), .B1(new_n947), .B2(new_n950), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n934), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n768), .A2(new_n783), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n764), .A2(new_n224), .B1(new_n758), .B2(new_n213), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n338), .B1(new_n775), .B2(new_n221), .ZN(new_n957));
  INV_X1    g0757(.A(G137), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n777), .A2(new_n219), .B1(new_n752), .B2(new_n958), .ZN(new_n959));
  NOR4_X1   g0759(.A1(new_n955), .A2(new_n956), .A3(new_n957), .A4(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n757), .ZN(new_n961));
  OAI221_X1 g0761(.A(new_n960), .B1(new_n822), .B2(new_n961), .C1(new_n319), .C2(new_n747), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n356), .B1(new_n961), .B2(new_n776), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n764), .A2(new_n536), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT46), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n758), .A2(new_n215), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n775), .A2(new_n415), .B1(new_n752), .B2(new_n769), .ZN(new_n967));
  NOR4_X1   g0767(.A1(new_n963), .A2(new_n965), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n968), .B1(new_n387), .B2(new_n777), .C1(new_n523), .C2(new_n747), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n768), .A2(new_n447), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n962), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT47), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n741), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n935), .A2(new_n790), .A3(new_n936), .ZN(new_n974));
  INV_X1    g0774(.A(new_n369), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n791), .B1(new_n209), .B2(new_n975), .C1(new_n246), .C2(new_n793), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT106), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n973), .A2(new_n816), .A3(new_n974), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n954), .A2(new_n978), .ZN(G387));
  NAND2_X1  g0779(.A1(new_n243), .A2(G45), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n691), .B(KEYINPUT107), .Z(new_n981));
  NOR2_X1   g0781(.A1(new_n367), .A2(G50), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(G45), .B1(new_n983), .B2(KEYINPUT50), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT50), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n982), .A2(new_n985), .B1(G68), .B2(G77), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n981), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n980), .A2(new_n987), .A3(new_n792), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(G107), .B2(new_n209), .C1(new_n692), .C2(new_n797), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n989), .A2(new_n791), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n781), .A2(G50), .B1(new_n369), .B2(new_n759), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n991), .B1(new_n213), .B2(new_n777), .C1(new_n415), .C2(new_n775), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(new_n327), .B2(new_n767), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n756), .A2(G159), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n764), .A2(new_n221), .B1(new_n752), .B2(new_n319), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT108), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n993), .A2(new_n338), .A3(new_n994), .A4(new_n996), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n747), .A2(new_n769), .B1(new_n523), .B2(new_n777), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT109), .Z(new_n999));
  OAI221_X1 g0799(.A(new_n999), .B1(new_n776), .B2(new_n768), .C1(new_n748), .C2(new_n961), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT48), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1001), .B1(new_n387), .B2(new_n758), .C1(new_n447), .C2(new_n764), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT49), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n834), .A2(G116), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n753), .A2(G326), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1004), .A2(new_n356), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  AND2_X1   g0807(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n997), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n734), .B(new_n990), .C1(new_n1009), .C2(new_n741), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n679), .A2(new_n790), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n1010), .A2(new_n1011), .B1(new_n932), .B2(new_n922), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n922), .A2(new_n731), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n922), .A2(new_n731), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1013), .A2(new_n689), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1012), .A2(new_n1015), .ZN(G393));
  NAND3_X1  g0816(.A1(new_n917), .A2(new_n932), .A3(new_n918), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n747), .A2(new_n776), .B1(new_n769), .B2(new_n779), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT52), .Z(new_n1019));
  INV_X1    g0819(.A(new_n777), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n338), .B(new_n1019), .C1(G294), .C2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n536), .B2(new_n758), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n764), .A2(new_n387), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n768), .A2(new_n523), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n775), .A2(new_n215), .B1(new_n752), .B2(new_n748), .ZN(new_n1025));
  NOR4_X1   g0825(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(G87), .A2(new_n834), .B1(new_n753), .B2(G143), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n367), .A2(new_n777), .B1(new_n219), .B2(new_n768), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1027), .B1(new_n1028), .B2(KEYINPUT111), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n747), .A2(new_n783), .B1(new_n319), .B2(new_n779), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT51), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n758), .A2(new_n221), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(new_n1028), .B2(KEYINPUT111), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1031), .A2(new_n338), .A3(new_n1033), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n1029), .B(new_n1034), .C1(G68), .C2(new_n765), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n741), .B1(new_n1026), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n908), .A2(new_n790), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n791), .B1(new_n415), .B2(new_n209), .C1(new_n793), .C2(new_n253), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n816), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT110), .Z(new_n1040));
  NAND3_X1  g0840(.A1(new_n1036), .A2(new_n1037), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1017), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(KEYINPUT112), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT112), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1017), .A2(new_n1044), .A3(new_n1041), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n917), .A2(new_n918), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n1014), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1048), .A2(new_n689), .A3(new_n923), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1046), .A2(new_n1049), .ZN(G390));
  NAND3_X1  g0850(.A1(new_n891), .A2(G330), .A3(new_n636), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n881), .A2(new_n635), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n876), .B1(new_n716), .B2(new_n806), .ZN(new_n1054));
  NOR4_X1   g0854(.A1(new_n886), .A2(new_n696), .A3(new_n807), .A4(new_n869), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n875), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n805), .A2(new_n380), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n726), .A2(new_n670), .A3(new_n1057), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n1058), .A2(new_n871), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n716), .A2(new_n806), .A3(new_n876), .ZN(new_n1060));
  AND3_X1   g0860(.A1(new_n657), .A2(new_n564), .A3(new_n658), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1061), .A2(new_n554), .A3(new_n520), .A4(new_n670), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n709), .B1(new_n1062), .B2(KEYINPUT31), .ZN(new_n1063));
  OAI211_X1 g0863(.A(G330), .B(new_n806), .C1(new_n1063), .C2(new_n885), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n869), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1059), .A2(new_n1060), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1056), .A2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n862), .A2(new_n854), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n853), .B2(new_n854), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n872), .A2(new_n858), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n869), .B1(new_n1058), .B2(new_n871), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n857), .B(KEYINPUT102), .Z(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n853), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n1069), .A2(new_n1070), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1055), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1074), .A2(new_n1060), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1053), .B(new_n1067), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1067), .A2(new_n1053), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT113), .ZN(new_n1080));
  OR2_X1    g0880(.A1(new_n1074), .A2(new_n1060), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n689), .B(new_n1078), .C1(new_n1080), .C2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n932), .ZN(new_n1085));
  XOR2_X1   g0885(.A(KEYINPUT54), .B(G143), .Z(new_n1086));
  AOI22_X1  g0886(.A1(new_n1020), .A2(new_n1086), .B1(new_n759), .B2(G159), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n958), .B2(new_n768), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT114), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n356), .B(new_n1089), .C1(G132), .C2(new_n781), .ZN(new_n1090));
  INV_X1    g0890(.A(G128), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1090), .B1(new_n1091), .B2(new_n779), .ZN(new_n1092));
  NOR3_X1   g0892(.A1(new_n764), .A2(KEYINPUT53), .A3(new_n319), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n775), .A2(new_n219), .ZN(new_n1094));
  OAI21_X1  g0894(.A(KEYINPUT53), .B1(new_n764), .B2(new_n319), .ZN(new_n1095));
  INV_X1    g0895(.A(G125), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1095), .B1(new_n1096), .B2(new_n752), .ZN(new_n1097));
  NOR4_X1   g0897(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .A4(new_n1097), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n338), .B(new_n1032), .C1(G283), .C2(new_n756), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n781), .A2(G116), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n765), .A2(G87), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n775), .A2(new_n213), .B1(new_n752), .B2(new_n447), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G107), .B2(new_n767), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .A4(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(G97), .B2(new_n1020), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n741), .B1(new_n1098), .B2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n816), .B(new_n1106), .C1(new_n1069), .C2(new_n739), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n817), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1108), .B1(new_n327), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1084), .A2(new_n1085), .A3(new_n1110), .ZN(G378));
  AOI21_X1  g0911(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1112));
  OAI21_X1  g0912(.A(KEYINPUT118), .B1(new_n1112), .B2(new_n1052), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n632), .A2(new_n630), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n332), .A2(new_n668), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1115), .B(new_n1116), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n1114), .A2(new_n376), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1117), .B1(new_n1114), .B2(new_n376), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT116), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n890), .A2(new_n696), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1122), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n877), .A2(new_n878), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(KEYINPUT101), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n877), .A2(new_n874), .A3(new_n878), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1124), .B1(new_n1128), .B2(new_n865), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n865), .B(new_n1124), .C1(new_n873), .C2(new_n879), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1123), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n880), .A2(new_n1122), .A3(new_n1121), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n1118), .A2(new_n1119), .A3(new_n1122), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n853), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n876), .B(new_n806), .C1(new_n1063), .C2(new_n885), .ZN(new_n1136));
  OAI21_X1  g0936(.A(KEYINPUT40), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n889), .A2(new_n887), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1134), .B1(new_n1139), .B2(G330), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1133), .A2(new_n1140), .A3(new_n1130), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n1132), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT118), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1078), .A2(new_n1143), .A3(new_n1053), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1113), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT57), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1113), .A2(new_n1144), .A3(KEYINPUT57), .A4(new_n1142), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1147), .A2(new_n689), .A3(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1132), .A2(new_n932), .A3(new_n1141), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n219), .B1(new_n256), .B2(G41), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n356), .B1(new_n752), .B2(new_n387), .C1(new_n224), .C2(new_n775), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n975), .A2(new_n777), .B1(new_n221), .B2(new_n764), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n768), .A2(new_n415), .B1(new_n758), .B2(new_n213), .ZN(new_n1154));
  NOR4_X1   g0954(.A1(new_n1152), .A2(new_n1153), .A3(G41), .A4(new_n1154), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n1155), .B1(new_n215), .B2(new_n747), .C1(new_n536), .C2(new_n779), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT58), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n768), .A2(new_n819), .B1(new_n779), .B2(new_n1096), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1086), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n747), .A2(new_n1091), .B1(new_n764), .B2(new_n1159), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1158), .B(new_n1160), .C1(G137), .C2(new_n1020), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n319), .B2(new_n758), .ZN(new_n1162));
  OR2_X1    g0962(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n834), .A2(G159), .ZN(new_n1164));
  AOI21_X1  g0964(.A(G41), .B1(new_n753), .B2(G124), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1163), .A2(new_n263), .A3(new_n1164), .A4(new_n1165), .ZN(new_n1166));
  AND2_X1   g0966(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1151), .B(new_n1157), .C1(new_n1166), .C2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n741), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n734), .B1(new_n817), .B2(new_n219), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT115), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1169), .B(new_n1171), .C1(new_n1120), .C2(new_n739), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1150), .A2(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT117), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1149), .A2(new_n1174), .ZN(G375));
  OAI22_X1  g0975(.A1(new_n975), .A2(new_n758), .B1(new_n536), .B2(new_n768), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n779), .A2(new_n447), .B1(new_n775), .B2(new_n221), .ZN(new_n1177));
  NOR3_X1   g0977(.A1(new_n1176), .A2(new_n1177), .A3(new_n338), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n781), .A2(G283), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n753), .A2(G303), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(G97), .A2(new_n765), .B1(new_n1020), .B2(G107), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n775), .A2(new_n224), .B1(new_n752), .B2(new_n1091), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n356), .B(new_n1183), .C1(G50), .C2(new_n759), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1184), .B1(new_n319), .B2(new_n777), .C1(new_n783), .C2(new_n764), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n1185), .A2(KEYINPUT119), .B1(G132), .B2(new_n756), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1186), .B1(KEYINPUT119), .B2(new_n1185), .C1(new_n768), .C2(new_n1159), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n747), .A2(new_n958), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1182), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n1189), .B(KEYINPUT120), .Z(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n741), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n869), .A2(new_n738), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n817), .A2(new_n213), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n816), .A4(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n1067), .B2(new_n932), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1052), .A2(new_n1056), .A3(new_n1066), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1080), .A2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1196), .B1(new_n1199), .B2(new_n929), .ZN(G381));
  INV_X1    g1000(.A(G375), .ZN(new_n1201));
  INV_X1    g1001(.A(G390), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n954), .A2(new_n978), .A3(new_n1202), .ZN(new_n1203));
  OR2_X1    g1003(.A1(G393), .A2(G396), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(G378), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(G381), .A2(G384), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1201), .A2(new_n1205), .A3(new_n1206), .A4(new_n1207), .ZN(G407));
  NAND2_X1  g1008(.A1(new_n1201), .A2(new_n1206), .ZN(new_n1209));
  OAI211_X1 g1009(.A(G407), .B(G213), .C1(G343), .C2(new_n1209), .ZN(G409));
  INV_X1    g1010(.A(new_n953), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n926), .A2(new_n930), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1211), .B1(new_n1212), .B2(new_n933), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n978), .ZN(new_n1214));
  OAI21_X1  g1014(.A(G390), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(G393), .A2(G396), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1204), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT125), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1204), .A2(KEYINPUT125), .A3(new_n1216), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1215), .A2(new_n1221), .A3(new_n1203), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1220), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n1215), .B2(new_n1203), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n665), .A2(G343), .ZN(new_n1227));
  INV_X1    g1027(.A(G384), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT60), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1197), .A2(new_n1229), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1230), .A2(KEYINPUT123), .A3(new_n1079), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT123), .B1(new_n1230), .B2(new_n1079), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n689), .B1(new_n1197), .B2(new_n1229), .ZN(new_n1233));
  NOR3_X1   g1033(.A1(new_n1231), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1196), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1228), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1232), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1233), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1230), .A2(KEYINPUT123), .A3(new_n1079), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1240), .A2(G384), .A3(new_n1196), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1236), .A2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1132), .A2(KEYINPUT121), .A3(new_n1141), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n932), .ZN(new_n1244));
  AOI21_X1  g1044(.A(KEYINPUT121), .B1(new_n1132), .B2(new_n1141), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1172), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(KEYINPUT122), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1113), .A2(new_n1144), .A3(new_n925), .A4(new_n1142), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT122), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1249), .B(new_n1172), .C1(new_n1244), .C2(new_n1245), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1247), .A2(new_n1248), .A3(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n1206), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1149), .A2(new_n1174), .A3(G378), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n1227), .B(new_n1242), .C1(new_n1252), .C2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT62), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1227), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1227), .A2(G2897), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT124), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1257), .B1(new_n1242), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1257), .ZN(new_n1260));
  AOI211_X1 g1060(.A(KEYINPUT124), .B(new_n1260), .C1(new_n1236), .C2(new_n1241), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n1259), .A2(new_n1261), .B1(new_n1258), .B2(new_n1242), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n1254), .A2(new_n1255), .B1(new_n1256), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1227), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1242), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1264), .A2(new_n1255), .A3(new_n1265), .A4(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT61), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1226), .B1(new_n1263), .B2(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(KEYINPUT63), .B1(new_n1256), .B2(new_n1262), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1256), .A2(new_n1266), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1226), .A2(KEYINPUT61), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1254), .A2(KEYINPUT63), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1273), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1270), .A2(new_n1276), .ZN(G405));
  NAND2_X1  g1077(.A1(G375), .A2(new_n1206), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT126), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1278), .B(new_n1279), .ZN(new_n1280));
  OR2_X1    g1080(.A1(new_n1242), .A2(KEYINPUT127), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1280), .A2(new_n1253), .A3(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1202), .B1(new_n954), .B2(new_n978), .ZN(new_n1283));
  AOI211_X1 g1083(.A(new_n1214), .B(G390), .C1(new_n934), .C2(new_n953), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1220), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1242), .A2(KEYINPUT127), .ZN(new_n1286));
  AND3_X1   g1086(.A1(new_n1285), .A2(new_n1222), .A3(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1286), .B1(new_n1285), .B2(new_n1222), .ZN(new_n1288));
  OR2_X1    g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1282), .A2(new_n1289), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1291), .A2(new_n1253), .A3(new_n1281), .A4(new_n1280), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(G402));
endmodule


