

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U548 ( .A1(G651), .A2(n644), .ZN(n646) );
  NOR2_X1 U549 ( .A1(G2084), .A2(n723), .ZN(n725) );
  AND2_X1 U550 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X4 U551 ( .A1(n535), .A2(n534), .ZN(G160) );
  BUF_X2 U552 ( .A(n575), .Z(n650) );
  XNOR2_X1 U553 ( .A(n747), .B(KEYINPUT32), .ZN(n757) );
  NAND2_X1 U554 ( .A1(n585), .A2(n584), .ZN(n955) );
  INV_X1 U555 ( .A(KEYINPUT29), .ZN(n716) );
  OR2_X1 U556 ( .A1(n684), .A2(G1384), .ZN(n685) );
  INV_X1 U557 ( .A(KEYINPUT17), .ZN(n529) );
  NOR2_X1 U558 ( .A1(G2104), .A2(G2105), .ZN(n530) );
  XOR2_X1 U559 ( .A(KEYINPUT31), .B(n733), .Z(n510) );
  NOR2_X1 U560 ( .A1(n512), .A2(n709), .ZN(n511) );
  AND2_X1 U561 ( .A1(n711), .A2(n944), .ZN(n512) );
  AND2_X1 U562 ( .A1(n941), .A2(n825), .ZN(n513) );
  AND2_X1 U563 ( .A1(n718), .A2(G1996), .ZN(n694) );
  NOR2_X1 U564 ( .A1(n750), .A2(n726), .ZN(n727) );
  INV_X1 U565 ( .A(G168), .ZN(n728) );
  AND2_X1 U566 ( .A1(n729), .A2(n728), .ZN(n732) );
  BUF_X1 U567 ( .A(n723), .Z(n738) );
  XNOR2_X1 U568 ( .A(n717), .B(n716), .ZN(n722) );
  NOR2_X1 U569 ( .A1(n773), .A2(G1966), .ZN(n750) );
  NOR2_X1 U570 ( .A1(KEYINPUT33), .A2(n761), .ZN(n762) );
  NOR2_X1 U571 ( .A1(n780), .A2(n781), .ZN(n693) );
  INV_X1 U572 ( .A(G2105), .ZN(n531) );
  OR2_X1 U573 ( .A1(n813), .A2(n513), .ZN(n814) );
  AND2_X2 U574 ( .A1(G2104), .A2(G2105), .ZN(n881) );
  OR2_X1 U575 ( .A1(n815), .A2(n814), .ZN(n828) );
  NAND2_X1 U576 ( .A1(n878), .A2(G137), .ZN(n533) );
  NOR2_X2 U577 ( .A1(G651), .A2(G543), .ZN(n635) );
  NAND2_X1 U578 ( .A1(n635), .A2(G89), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n514), .B(KEYINPUT4), .ZN(n516) );
  XOR2_X1 U580 ( .A(G543), .B(KEYINPUT0), .Z(n644) );
  INV_X1 U581 ( .A(G651), .ZN(n518) );
  NOR2_X1 U582 ( .A1(n644), .A2(n518), .ZN(n589) );
  BUF_X1 U583 ( .A(n589), .Z(n638) );
  NAND2_X1 U584 ( .A1(G76), .A2(n638), .ZN(n515) );
  NAND2_X1 U585 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U586 ( .A(n517), .B(KEYINPUT5), .ZN(n524) );
  NOR2_X1 U587 ( .A1(G543), .A2(n518), .ZN(n519) );
  XOR2_X1 U588 ( .A(KEYINPUT1), .B(n519), .Z(n575) );
  NAND2_X1 U589 ( .A1(G63), .A2(n650), .ZN(n521) );
  NAND2_X1 U590 ( .A1(G51), .A2(n646), .ZN(n520) );
  NAND2_X1 U591 ( .A1(n521), .A2(n520), .ZN(n522) );
  XOR2_X1 U592 ( .A(KEYINPUT6), .B(n522), .Z(n523) );
  NAND2_X1 U593 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U594 ( .A(n525), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U595 ( .A1(n881), .A2(G113), .ZN(n528) );
  AND2_X4 U596 ( .A1(n531), .A2(G2104), .ZN(n877) );
  NAND2_X1 U597 ( .A1(G101), .A2(n877), .ZN(n526) );
  XOR2_X1 U598 ( .A(KEYINPUT23), .B(n526), .Z(n527) );
  NAND2_X1 U599 ( .A1(n528), .A2(n527), .ZN(n535) );
  XNOR2_X2 U600 ( .A(n530), .B(n529), .ZN(n878) );
  NOR2_X1 U601 ( .A1(G2104), .A2(n531), .ZN(n567) );
  BUF_X1 U602 ( .A(n567), .Z(n882) );
  NAND2_X1 U603 ( .A1(G125), .A2(n882), .ZN(n532) );
  NAND2_X1 U604 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U605 ( .A1(G85), .A2(n635), .ZN(n537) );
  NAND2_X1 U606 ( .A1(G72), .A2(n638), .ZN(n536) );
  NAND2_X1 U607 ( .A1(n537), .A2(n536), .ZN(n541) );
  NAND2_X1 U608 ( .A1(G60), .A2(n650), .ZN(n539) );
  NAND2_X1 U609 ( .A1(G47), .A2(n646), .ZN(n538) );
  NAND2_X1 U610 ( .A1(n539), .A2(n538), .ZN(n540) );
  OR2_X1 U611 ( .A1(n541), .A2(n540), .ZN(G290) );
  XOR2_X1 U612 ( .A(G2427), .B(G2435), .Z(n543) );
  XNOR2_X1 U613 ( .A(G2454), .B(G2443), .ZN(n542) );
  XNOR2_X1 U614 ( .A(n543), .B(n542), .ZN(n550) );
  XOR2_X1 U615 ( .A(G2451), .B(KEYINPUT99), .Z(n545) );
  XNOR2_X1 U616 ( .A(G2430), .B(G2438), .ZN(n544) );
  XNOR2_X1 U617 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U618 ( .A(n546), .B(G2446), .Z(n548) );
  XNOR2_X1 U619 ( .A(G1348), .B(G1341), .ZN(n547) );
  XNOR2_X1 U620 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U621 ( .A(n550), .B(n549), .ZN(n551) );
  AND2_X1 U622 ( .A1(n551), .A2(G14), .ZN(G401) );
  NAND2_X1 U623 ( .A1(G64), .A2(n650), .ZN(n553) );
  NAND2_X1 U624 ( .A1(G52), .A2(n646), .ZN(n552) );
  NAND2_X1 U625 ( .A1(n553), .A2(n552), .ZN(n558) );
  NAND2_X1 U626 ( .A1(G90), .A2(n635), .ZN(n555) );
  NAND2_X1 U627 ( .A1(G77), .A2(n638), .ZN(n554) );
  NAND2_X1 U628 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U629 ( .A(KEYINPUT9), .B(n556), .Z(n557) );
  NOR2_X1 U630 ( .A1(n558), .A2(n557), .ZN(G171) );
  AND2_X1 U631 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U632 ( .A1(G111), .A2(n881), .ZN(n560) );
  NAND2_X1 U633 ( .A1(G135), .A2(n878), .ZN(n559) );
  NAND2_X1 U634 ( .A1(n560), .A2(n559), .ZN(n563) );
  NAND2_X1 U635 ( .A1(n882), .A2(G123), .ZN(n561) );
  XOR2_X1 U636 ( .A(KEYINPUT18), .B(n561), .Z(n562) );
  NOR2_X1 U637 ( .A1(n563), .A2(n562), .ZN(n565) );
  NAND2_X1 U638 ( .A1(n877), .A2(G99), .ZN(n564) );
  NAND2_X1 U639 ( .A1(n565), .A2(n564), .ZN(n995) );
  XNOR2_X1 U640 ( .A(G2096), .B(n995), .ZN(n566) );
  OR2_X1 U641 ( .A1(G2100), .A2(n566), .ZN(G156) );
  NAND2_X1 U642 ( .A1(n878), .A2(G138), .ZN(n572) );
  NAND2_X1 U643 ( .A1(G126), .A2(n567), .ZN(n569) );
  NAND2_X1 U644 ( .A1(G114), .A2(n881), .ZN(n568) );
  NAND2_X1 U645 ( .A1(n569), .A2(n568), .ZN(n571) );
  AND2_X1 U646 ( .A1(G102), .A2(n877), .ZN(n570) );
  NOR2_X1 U647 ( .A1(n571), .A2(n570), .ZN(n684) );
  AND2_X1 U648 ( .A1(n572), .A2(n684), .ZN(G164) );
  INV_X1 U649 ( .A(G132), .ZN(G219) );
  INV_X1 U650 ( .A(G82), .ZN(G220) );
  XOR2_X1 U651 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U652 ( .A1(G7), .A2(G661), .ZN(n573) );
  XNOR2_X1 U653 ( .A(n573), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U654 ( .A(G223), .ZN(n831) );
  NAND2_X1 U655 ( .A1(n831), .A2(G567), .ZN(n574) );
  XOR2_X1 U656 ( .A(KEYINPUT11), .B(n574), .Z(G234) );
  NAND2_X1 U657 ( .A1(n650), .A2(G56), .ZN(n576) );
  XOR2_X1 U658 ( .A(KEYINPUT14), .B(n576), .Z(n582) );
  NAND2_X1 U659 ( .A1(n635), .A2(G81), .ZN(n577) );
  XNOR2_X1 U660 ( .A(n577), .B(KEYINPUT12), .ZN(n579) );
  NAND2_X1 U661 ( .A1(G68), .A2(n589), .ZN(n578) );
  NAND2_X1 U662 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U663 ( .A(KEYINPUT13), .B(n580), .Z(n581) );
  NOR2_X1 U664 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U665 ( .A(n583), .B(KEYINPUT68), .ZN(n585) );
  NAND2_X1 U666 ( .A1(G43), .A2(n646), .ZN(n584) );
  INV_X1 U667 ( .A(n955), .ZN(n586) );
  XOR2_X1 U668 ( .A(G860), .B(KEYINPUT69), .Z(n612) );
  NAND2_X1 U669 ( .A1(n586), .A2(n612), .ZN(G153) );
  XOR2_X1 U670 ( .A(G171), .B(KEYINPUT70), .Z(G301) );
  NAND2_X1 U671 ( .A1(G54), .A2(n646), .ZN(n594) );
  NAND2_X1 U672 ( .A1(G92), .A2(n635), .ZN(n588) );
  NAND2_X1 U673 ( .A1(G66), .A2(n650), .ZN(n587) );
  NAND2_X1 U674 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U675 ( .A1(G79), .A2(n589), .ZN(n590) );
  XNOR2_X1 U676 ( .A(KEYINPUT71), .B(n590), .ZN(n591) );
  NOR2_X1 U677 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U678 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U679 ( .A(n595), .B(KEYINPUT15), .ZN(n596) );
  XNOR2_X1 U680 ( .A(KEYINPUT72), .B(n596), .ZN(n619) );
  NOR2_X1 U681 ( .A1(G868), .A2(n619), .ZN(n597) );
  XNOR2_X1 U682 ( .A(n597), .B(KEYINPUT73), .ZN(n599) );
  NAND2_X1 U683 ( .A1(G301), .A2(G868), .ZN(n598) );
  NAND2_X1 U684 ( .A1(n599), .A2(n598), .ZN(G284) );
  NAND2_X1 U685 ( .A1(G91), .A2(n635), .ZN(n601) );
  NAND2_X1 U686 ( .A1(G78), .A2(n638), .ZN(n600) );
  NAND2_X1 U687 ( .A1(n601), .A2(n600), .ZN(n604) );
  NAND2_X1 U688 ( .A1(n650), .A2(G65), .ZN(n602) );
  XOR2_X1 U689 ( .A(KEYINPUT66), .B(n602), .Z(n603) );
  NOR2_X1 U690 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U691 ( .A1(n646), .A2(G53), .ZN(n605) );
  NAND2_X1 U692 ( .A1(n606), .A2(n605), .ZN(G299) );
  INV_X1 U693 ( .A(G868), .ZN(n607) );
  NOR2_X1 U694 ( .A1(G286), .A2(n607), .ZN(n609) );
  NOR2_X1 U695 ( .A1(G868), .A2(G299), .ZN(n608) );
  NOR2_X1 U696 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U697 ( .A(KEYINPUT74), .B(n610), .ZN(G297) );
  INV_X1 U698 ( .A(n619), .ZN(n937) );
  INV_X1 U699 ( .A(G559), .ZN(n611) );
  NOR2_X1 U700 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U701 ( .A1(n937), .A2(n613), .ZN(n614) );
  XNOR2_X1 U702 ( .A(n614), .B(KEYINPUT75), .ZN(n615) );
  XNOR2_X1 U703 ( .A(n615), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U704 ( .A1(G868), .A2(n955), .ZN(n618) );
  NAND2_X1 U705 ( .A1(n619), .A2(G868), .ZN(n616) );
  NOR2_X1 U706 ( .A1(G559), .A2(n616), .ZN(n617) );
  NOR2_X1 U707 ( .A1(n618), .A2(n617), .ZN(G282) );
  NAND2_X1 U708 ( .A1(G559), .A2(n619), .ZN(n664) );
  XNOR2_X1 U709 ( .A(n955), .B(n664), .ZN(n620) );
  NOR2_X1 U710 ( .A1(n620), .A2(G860), .ZN(n628) );
  NAND2_X1 U711 ( .A1(n635), .A2(G93), .ZN(n621) );
  XNOR2_X1 U712 ( .A(n621), .B(KEYINPUT76), .ZN(n623) );
  NAND2_X1 U713 ( .A1(G67), .A2(n650), .ZN(n622) );
  NAND2_X1 U714 ( .A1(n623), .A2(n622), .ZN(n627) );
  NAND2_X1 U715 ( .A1(G80), .A2(n638), .ZN(n625) );
  NAND2_X1 U716 ( .A1(G55), .A2(n646), .ZN(n624) );
  NAND2_X1 U717 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U718 ( .A1(n627), .A2(n626), .ZN(n660) );
  XNOR2_X1 U719 ( .A(n628), .B(n660), .ZN(G145) );
  NAND2_X1 U720 ( .A1(G88), .A2(n635), .ZN(n630) );
  NAND2_X1 U721 ( .A1(G75), .A2(n638), .ZN(n629) );
  NAND2_X1 U722 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U723 ( .A1(G62), .A2(n650), .ZN(n632) );
  NAND2_X1 U724 ( .A1(G50), .A2(n646), .ZN(n631) );
  NAND2_X1 U725 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U726 ( .A1(n634), .A2(n633), .ZN(G166) );
  NAND2_X1 U727 ( .A1(G86), .A2(n635), .ZN(n637) );
  NAND2_X1 U728 ( .A1(G61), .A2(n650), .ZN(n636) );
  NAND2_X1 U729 ( .A1(n637), .A2(n636), .ZN(n641) );
  NAND2_X1 U730 ( .A1(n638), .A2(G73), .ZN(n639) );
  XOR2_X1 U731 ( .A(KEYINPUT2), .B(n639), .Z(n640) );
  NOR2_X1 U732 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U733 ( .A1(n646), .A2(G48), .ZN(n642) );
  NAND2_X1 U734 ( .A1(n643), .A2(n642), .ZN(G305) );
  NAND2_X1 U735 ( .A1(n644), .A2(G87), .ZN(n645) );
  XNOR2_X1 U736 ( .A(KEYINPUT78), .B(n645), .ZN(n653) );
  NAND2_X1 U737 ( .A1(G49), .A2(n646), .ZN(n648) );
  NAND2_X1 U738 ( .A1(G74), .A2(G651), .ZN(n647) );
  NAND2_X1 U739 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U740 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U741 ( .A(KEYINPUT77), .B(n651), .Z(n652) );
  NAND2_X1 U742 ( .A1(n653), .A2(n652), .ZN(G288) );
  NOR2_X1 U743 ( .A1(G868), .A2(n660), .ZN(n654) );
  XNOR2_X1 U744 ( .A(n654), .B(KEYINPUT81), .ZN(n667) );
  XNOR2_X1 U745 ( .A(KEYINPUT79), .B(KEYINPUT19), .ZN(n656) );
  XNOR2_X1 U746 ( .A(G290), .B(G166), .ZN(n655) );
  XNOR2_X1 U747 ( .A(n656), .B(n655), .ZN(n659) );
  INV_X1 U748 ( .A(G299), .ZN(n944) );
  XNOR2_X1 U749 ( .A(n944), .B(G305), .ZN(n657) );
  XNOR2_X1 U750 ( .A(n657), .B(G288), .ZN(n658) );
  XNOR2_X1 U751 ( .A(n659), .B(n658), .ZN(n662) );
  XNOR2_X1 U752 ( .A(n955), .B(n660), .ZN(n661) );
  XNOR2_X1 U753 ( .A(n662), .B(n661), .ZN(n900) );
  XOR2_X1 U754 ( .A(n900), .B(KEYINPUT80), .Z(n663) );
  XNOR2_X1 U755 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U756 ( .A1(G868), .A2(n665), .ZN(n666) );
  NAND2_X1 U757 ( .A1(n667), .A2(n666), .ZN(G295) );
  NAND2_X1 U758 ( .A1(G2078), .A2(G2084), .ZN(n668) );
  XOR2_X1 U759 ( .A(KEYINPUT20), .B(n668), .Z(n669) );
  NAND2_X1 U760 ( .A1(G2090), .A2(n669), .ZN(n670) );
  XNOR2_X1 U761 ( .A(KEYINPUT21), .B(n670), .ZN(n671) );
  NAND2_X1 U762 ( .A1(n671), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U763 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U764 ( .A(KEYINPUT67), .B(G57), .ZN(G237) );
  NOR2_X1 U765 ( .A1(G220), .A2(G219), .ZN(n672) );
  XNOR2_X1 U766 ( .A(KEYINPUT22), .B(n672), .ZN(n673) );
  NAND2_X1 U767 ( .A1(n673), .A2(G96), .ZN(n674) );
  NOR2_X1 U768 ( .A1(G218), .A2(n674), .ZN(n675) );
  XOR2_X1 U769 ( .A(KEYINPUT82), .B(n675), .Z(n912) );
  NAND2_X1 U770 ( .A1(n912), .A2(G2106), .ZN(n676) );
  XOR2_X1 U771 ( .A(KEYINPUT83), .B(n676), .Z(n680) );
  NAND2_X1 U772 ( .A1(G108), .A2(G120), .ZN(n677) );
  NOR2_X1 U773 ( .A1(G237), .A2(n677), .ZN(n678) );
  NAND2_X1 U774 ( .A1(G69), .A2(n678), .ZN(n911) );
  NAND2_X1 U775 ( .A1(G567), .A2(n911), .ZN(n679) );
  NAND2_X1 U776 ( .A1(n680), .A2(n679), .ZN(n835) );
  NAND2_X1 U777 ( .A1(G483), .A2(G661), .ZN(n681) );
  NOR2_X1 U778 ( .A1(n835), .A2(n681), .ZN(n834) );
  NAND2_X1 U779 ( .A1(n834), .A2(G36), .ZN(G176) );
  INV_X1 U780 ( .A(G166), .ZN(G303) );
  NAND2_X1 U781 ( .A1(G160), .A2(G40), .ZN(n780) );
  INV_X1 U782 ( .A(G1384), .ZN(n682) );
  AND2_X1 U783 ( .A1(G138), .A2(n682), .ZN(n683) );
  NAND2_X1 U784 ( .A1(n878), .A2(n683), .ZN(n686) );
  NAND2_X1 U785 ( .A1(n686), .A2(n685), .ZN(n688) );
  INV_X1 U786 ( .A(KEYINPUT64), .ZN(n687) );
  XNOR2_X1 U787 ( .A(n688), .B(n687), .ZN(n781) );
  INV_X1 U788 ( .A(n693), .ZN(n723) );
  NAND2_X1 U789 ( .A1(n723), .A2(G8), .ZN(n689) );
  XNOR2_X2 U790 ( .A(n689), .B(KEYINPUT88), .ZN(n773) );
  NOR2_X1 U791 ( .A1(G1981), .A2(G305), .ZN(n690) );
  XOR2_X1 U792 ( .A(n690), .B(KEYINPUT24), .Z(n691) );
  NOR2_X1 U793 ( .A1(n773), .A2(n691), .ZN(n692) );
  XOR2_X1 U794 ( .A(KEYINPUT89), .B(n692), .Z(n779) );
  XNOR2_X1 U795 ( .A(G1981), .B(G305), .ZN(n949) );
  BUF_X2 U796 ( .A(n693), .Z(n718) );
  XNOR2_X1 U797 ( .A(n694), .B(KEYINPUT26), .ZN(n695) );
  INV_X1 U798 ( .A(n695), .ZN(n697) );
  NAND2_X1 U799 ( .A1(n738), .A2(G1341), .ZN(n696) );
  NAND2_X1 U800 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U801 ( .A1(n955), .A2(n698), .ZN(n699) );
  XNOR2_X1 U802 ( .A(n699), .B(KEYINPUT65), .ZN(n703) );
  NAND2_X1 U803 ( .A1(G2067), .A2(n718), .ZN(n701) );
  NAND2_X1 U804 ( .A1(G1348), .A2(n738), .ZN(n700) );
  NAND2_X1 U805 ( .A1(n701), .A2(n700), .ZN(n708) );
  AND2_X1 U806 ( .A1(n937), .A2(n708), .ZN(n702) );
  NOR2_X1 U807 ( .A1(n703), .A2(n702), .ZN(n704) );
  INV_X1 U808 ( .A(n704), .ZN(n710) );
  NAND2_X1 U809 ( .A1(n718), .A2(G2072), .ZN(n705) );
  XNOR2_X1 U810 ( .A(n705), .B(KEYINPUT27), .ZN(n707) );
  INV_X1 U811 ( .A(G1956), .ZN(n913) );
  NOR2_X1 U812 ( .A1(n913), .A2(n718), .ZN(n706) );
  NOR2_X1 U813 ( .A1(n707), .A2(n706), .ZN(n711) );
  NOR2_X1 U814 ( .A1(n937), .A2(n708), .ZN(n709) );
  NAND2_X1 U815 ( .A1(n710), .A2(n511), .ZN(n715) );
  NOR2_X1 U816 ( .A1(n711), .A2(n944), .ZN(n713) );
  XNOR2_X1 U817 ( .A(KEYINPUT91), .B(KEYINPUT28), .ZN(n712) );
  XNOR2_X1 U818 ( .A(n713), .B(n712), .ZN(n714) );
  NAND2_X1 U819 ( .A1(n715), .A2(n714), .ZN(n717) );
  XNOR2_X1 U820 ( .A(G2078), .B(KEYINPUT25), .ZN(n972) );
  NOR2_X1 U821 ( .A1(n738), .A2(n972), .ZN(n720) );
  INV_X1 U822 ( .A(G1961), .ZN(n939) );
  NOR2_X1 U823 ( .A1(n718), .A2(n939), .ZN(n719) );
  NOR2_X1 U824 ( .A1(n720), .A2(n719), .ZN(n730) );
  NAND2_X1 U825 ( .A1(G171), .A2(n730), .ZN(n721) );
  NAND2_X1 U826 ( .A1(n722), .A2(n721), .ZN(n734) );
  INV_X1 U827 ( .A(KEYINPUT90), .ZN(n724) );
  XNOR2_X1 U828 ( .A(n725), .B(n724), .ZN(n752) );
  NAND2_X1 U829 ( .A1(n752), .A2(G8), .ZN(n726) );
  XNOR2_X1 U830 ( .A(n727), .B(KEYINPUT30), .ZN(n729) );
  NOR2_X1 U831 ( .A1(G171), .A2(n730), .ZN(n731) );
  NOR2_X1 U832 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U833 ( .A1(n734), .A2(n510), .ZN(n735) );
  XNOR2_X1 U834 ( .A(n735), .B(KEYINPUT92), .ZN(n748) );
  AND2_X1 U835 ( .A1(G286), .A2(G8), .ZN(n736) );
  NAND2_X1 U836 ( .A1(n748), .A2(n736), .ZN(n746) );
  INV_X1 U837 ( .A(G8), .ZN(n744) );
  NOR2_X1 U838 ( .A1(n773), .A2(G1971), .ZN(n737) );
  XOR2_X1 U839 ( .A(KEYINPUT93), .B(n737), .Z(n740) );
  NOR2_X1 U840 ( .A1(G2090), .A2(n738), .ZN(n739) );
  NOR2_X1 U841 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U842 ( .A(n741), .B(KEYINPUT94), .ZN(n742) );
  NAND2_X1 U843 ( .A1(n742), .A2(G303), .ZN(n743) );
  OR2_X1 U844 ( .A1(n744), .A2(n743), .ZN(n745) );
  BUF_X1 U845 ( .A(n748), .Z(n749) );
  INV_X1 U846 ( .A(n749), .ZN(n751) );
  NOR2_X1 U847 ( .A1(n751), .A2(n750), .ZN(n755) );
  INV_X1 U848 ( .A(n752), .ZN(n753) );
  NAND2_X1 U849 ( .A1(G8), .A2(n753), .ZN(n754) );
  NAND2_X1 U850 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U851 ( .A1(n757), .A2(n756), .ZN(n771) );
  NOR2_X1 U852 ( .A1(G1971), .A2(G303), .ZN(n758) );
  NOR2_X1 U853 ( .A1(G1976), .A2(G288), .ZN(n962) );
  NOR2_X1 U854 ( .A1(n758), .A2(n962), .ZN(n759) );
  NAND2_X1 U855 ( .A1(n771), .A2(n759), .ZN(n760) );
  NAND2_X1 U856 ( .A1(G1976), .A2(G288), .ZN(n959) );
  NAND2_X1 U857 ( .A1(n760), .A2(n959), .ZN(n761) );
  INV_X1 U858 ( .A(n773), .ZN(n763) );
  NAND2_X1 U859 ( .A1(n762), .A2(n763), .ZN(n766) );
  NAND2_X1 U860 ( .A1(n962), .A2(n763), .ZN(n764) );
  NAND2_X1 U861 ( .A1(n764), .A2(KEYINPUT33), .ZN(n765) );
  NAND2_X1 U862 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U863 ( .A(n767), .B(KEYINPUT95), .ZN(n768) );
  NOR2_X1 U864 ( .A1(n949), .A2(n768), .ZN(n776) );
  NOR2_X1 U865 ( .A1(G2090), .A2(G303), .ZN(n769) );
  NAND2_X1 U866 ( .A1(G8), .A2(n769), .ZN(n770) );
  NAND2_X1 U867 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U868 ( .A1(n773), .A2(n772), .ZN(n774) );
  XOR2_X1 U869 ( .A(KEYINPUT96), .B(n774), .Z(n775) );
  NOR2_X2 U870 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U871 ( .A(n777), .B(KEYINPUT97), .ZN(n778) );
  NOR2_X1 U872 ( .A1(n779), .A2(n778), .ZN(n815) );
  INV_X1 U873 ( .A(n781), .ZN(n782) );
  NOR2_X1 U874 ( .A1(n780), .A2(n782), .ZN(n825) );
  XNOR2_X1 U875 ( .A(KEYINPUT37), .B(G2067), .ZN(n823) );
  NAND2_X1 U876 ( .A1(G104), .A2(n877), .ZN(n784) );
  NAND2_X1 U877 ( .A1(G140), .A2(n878), .ZN(n783) );
  NAND2_X1 U878 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U879 ( .A(KEYINPUT34), .B(n785), .ZN(n790) );
  NAND2_X1 U880 ( .A1(G116), .A2(n881), .ZN(n787) );
  NAND2_X1 U881 ( .A1(G128), .A2(n882), .ZN(n786) );
  NAND2_X1 U882 ( .A1(n787), .A2(n786), .ZN(n788) );
  XOR2_X1 U883 ( .A(KEYINPUT35), .B(n788), .Z(n789) );
  NOR2_X1 U884 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U885 ( .A(KEYINPUT36), .B(n791), .ZN(n897) );
  NOR2_X1 U886 ( .A1(n823), .A2(n897), .ZN(n1009) );
  NAND2_X1 U887 ( .A1(n825), .A2(n1009), .ZN(n821) );
  NAND2_X1 U888 ( .A1(G131), .A2(n878), .ZN(n792) );
  XNOR2_X1 U889 ( .A(n792), .B(KEYINPUT86), .ZN(n799) );
  NAND2_X1 U890 ( .A1(G95), .A2(n877), .ZN(n794) );
  NAND2_X1 U891 ( .A1(G119), .A2(n882), .ZN(n793) );
  NAND2_X1 U892 ( .A1(n794), .A2(n793), .ZN(n797) );
  NAND2_X1 U893 ( .A1(G107), .A2(n881), .ZN(n795) );
  XNOR2_X1 U894 ( .A(KEYINPUT85), .B(n795), .ZN(n796) );
  NOR2_X1 U895 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U896 ( .A1(n799), .A2(n798), .ZN(n864) );
  AND2_X1 U897 ( .A1(n864), .A2(G1991), .ZN(n809) );
  NAND2_X1 U898 ( .A1(G117), .A2(n881), .ZN(n801) );
  NAND2_X1 U899 ( .A1(G141), .A2(n878), .ZN(n800) );
  NAND2_X1 U900 ( .A1(n801), .A2(n800), .ZN(n805) );
  NAND2_X1 U901 ( .A1(G105), .A2(n877), .ZN(n802) );
  XNOR2_X1 U902 ( .A(n802), .B(KEYINPUT87), .ZN(n803) );
  XNOR2_X1 U903 ( .A(n803), .B(KEYINPUT38), .ZN(n804) );
  NOR2_X1 U904 ( .A1(n805), .A2(n804), .ZN(n807) );
  NAND2_X1 U905 ( .A1(n882), .A2(G129), .ZN(n806) );
  NAND2_X1 U906 ( .A1(n807), .A2(n806), .ZN(n865) );
  AND2_X1 U907 ( .A1(n865), .A2(G1996), .ZN(n808) );
  NOR2_X1 U908 ( .A1(n809), .A2(n808), .ZN(n1000) );
  INV_X1 U909 ( .A(n825), .ZN(n810) );
  NOR2_X1 U910 ( .A1(n1000), .A2(n810), .ZN(n818) );
  INV_X1 U911 ( .A(n818), .ZN(n811) );
  NAND2_X1 U912 ( .A1(n821), .A2(n811), .ZN(n813) );
  XNOR2_X1 U913 ( .A(G1986), .B(KEYINPUT84), .ZN(n812) );
  XNOR2_X1 U914 ( .A(n812), .B(G290), .ZN(n941) );
  NOR2_X1 U915 ( .A1(G1996), .A2(n865), .ZN(n1002) );
  NOR2_X1 U916 ( .A1(G1991), .A2(n864), .ZN(n998) );
  NOR2_X1 U917 ( .A1(G1986), .A2(G290), .ZN(n816) );
  NOR2_X1 U918 ( .A1(n998), .A2(n816), .ZN(n817) );
  NOR2_X1 U919 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U920 ( .A1(n1002), .A2(n819), .ZN(n820) );
  XNOR2_X1 U921 ( .A(n820), .B(KEYINPUT39), .ZN(n822) );
  NAND2_X1 U922 ( .A1(n822), .A2(n821), .ZN(n824) );
  NAND2_X1 U923 ( .A1(n823), .A2(n897), .ZN(n1006) );
  NAND2_X1 U924 ( .A1(n824), .A2(n1006), .ZN(n826) );
  NAND2_X1 U925 ( .A1(n826), .A2(n825), .ZN(n827) );
  NAND2_X1 U926 ( .A1(n828), .A2(n827), .ZN(n830) );
  XNOR2_X1 U927 ( .A(KEYINPUT98), .B(KEYINPUT40), .ZN(n829) );
  XNOR2_X1 U928 ( .A(n830), .B(n829), .ZN(G329) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n831), .ZN(G217) );
  AND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n832) );
  NAND2_X1 U931 ( .A1(G661), .A2(n832), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n833) );
  NAND2_X1 U933 ( .A1(n834), .A2(n833), .ZN(G188) );
  XOR2_X1 U934 ( .A(G120), .B(KEYINPUT100), .Z(G236) );
  XNOR2_X1 U935 ( .A(KEYINPUT101), .B(n835), .ZN(G319) );
  XOR2_X1 U936 ( .A(KEYINPUT104), .B(G1961), .Z(n837) );
  XNOR2_X1 U937 ( .A(G1981), .B(G1966), .ZN(n836) );
  XNOR2_X1 U938 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U939 ( .A(n838), .B(KEYINPUT41), .Z(n840) );
  XNOR2_X1 U940 ( .A(G1996), .B(G1991), .ZN(n839) );
  XNOR2_X1 U941 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U942 ( .A(G1956), .B(G1971), .Z(n842) );
  XNOR2_X1 U943 ( .A(G1986), .B(G1976), .ZN(n841) );
  XNOR2_X1 U944 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U945 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U946 ( .A(KEYINPUT103), .B(G2474), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n846), .B(n845), .ZN(G229) );
  XOR2_X1 U948 ( .A(G2096), .B(KEYINPUT102), .Z(n848) );
  XNOR2_X1 U949 ( .A(G2090), .B(KEYINPUT43), .ZN(n847) );
  XNOR2_X1 U950 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U951 ( .A(n849), .B(KEYINPUT42), .Z(n851) );
  XNOR2_X1 U952 ( .A(G2067), .B(G2072), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U954 ( .A(G2678), .B(G2100), .Z(n853) );
  XNOR2_X1 U955 ( .A(G2078), .B(G2084), .ZN(n852) );
  XNOR2_X1 U956 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U957 ( .A(n855), .B(n854), .ZN(G227) );
  NAND2_X1 U958 ( .A1(G124), .A2(n882), .ZN(n856) );
  XNOR2_X1 U959 ( .A(n856), .B(KEYINPUT44), .ZN(n859) );
  NAND2_X1 U960 ( .A1(G112), .A2(n881), .ZN(n857) );
  XOR2_X1 U961 ( .A(KEYINPUT105), .B(n857), .Z(n858) );
  NAND2_X1 U962 ( .A1(n859), .A2(n858), .ZN(n863) );
  NAND2_X1 U963 ( .A1(G100), .A2(n877), .ZN(n861) );
  NAND2_X1 U964 ( .A1(G136), .A2(n878), .ZN(n860) );
  NAND2_X1 U965 ( .A1(n861), .A2(n860), .ZN(n862) );
  NOR2_X1 U966 ( .A1(n863), .A2(n862), .ZN(G162) );
  XNOR2_X1 U967 ( .A(n865), .B(n864), .ZN(n896) );
  NAND2_X1 U968 ( .A1(G106), .A2(n877), .ZN(n867) );
  NAND2_X1 U969 ( .A1(G142), .A2(n878), .ZN(n866) );
  NAND2_X1 U970 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U971 ( .A(n868), .B(KEYINPUT45), .ZN(n870) );
  NAND2_X1 U972 ( .A1(G118), .A2(n881), .ZN(n869) );
  NAND2_X1 U973 ( .A1(n870), .A2(n869), .ZN(n873) );
  NAND2_X1 U974 ( .A1(n882), .A2(G130), .ZN(n871) );
  XOR2_X1 U975 ( .A(KEYINPUT106), .B(n871), .Z(n872) );
  NOR2_X1 U976 ( .A1(n873), .A2(n872), .ZN(n892) );
  XOR2_X1 U977 ( .A(KEYINPUT46), .B(KEYINPUT107), .Z(n875) );
  XNOR2_X1 U978 ( .A(KEYINPUT109), .B(KEYINPUT48), .ZN(n874) );
  XNOR2_X1 U979 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U980 ( .A(n995), .B(n876), .ZN(n890) );
  NAND2_X1 U981 ( .A1(G103), .A2(n877), .ZN(n880) );
  NAND2_X1 U982 ( .A1(G139), .A2(n878), .ZN(n879) );
  NAND2_X1 U983 ( .A1(n880), .A2(n879), .ZN(n888) );
  NAND2_X1 U984 ( .A1(G115), .A2(n881), .ZN(n884) );
  NAND2_X1 U985 ( .A1(G127), .A2(n882), .ZN(n883) );
  NAND2_X1 U986 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U987 ( .A(KEYINPUT108), .B(n885), .Z(n886) );
  XNOR2_X1 U988 ( .A(KEYINPUT47), .B(n886), .ZN(n887) );
  NOR2_X1 U989 ( .A1(n888), .A2(n887), .ZN(n991) );
  XNOR2_X1 U990 ( .A(G164), .B(n991), .ZN(n889) );
  XNOR2_X1 U991 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U992 ( .A(n892), .B(n891), .Z(n894) );
  XNOR2_X1 U993 ( .A(G160), .B(G162), .ZN(n893) );
  XNOR2_X1 U994 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n898) );
  XOR2_X1 U996 ( .A(n898), .B(n897), .Z(n899) );
  NOR2_X1 U997 ( .A1(G37), .A2(n899), .ZN(G395) );
  XOR2_X1 U998 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n902) );
  XNOR2_X1 U999 ( .A(G171), .B(n900), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(n902), .B(n901), .ZN(n904) );
  XOR2_X1 U1001 ( .A(G286), .B(n937), .Z(n903) );
  XNOR2_X1 U1002 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n905), .ZN(G397) );
  NOR2_X1 U1004 ( .A1(G229), .A2(G227), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(n906), .ZN(n907) );
  NOR2_X1 U1006 ( .A1(G401), .A2(n907), .ZN(n909) );
  NOR2_X1 U1007 ( .A1(G395), .A2(G397), .ZN(n908) );
  AND2_X1 U1008 ( .A1(n909), .A2(n908), .ZN(n910) );
  NAND2_X1 U1009 ( .A1(G319), .A2(n910), .ZN(G225) );
  XOR2_X1 U1010 ( .A(KEYINPUT112), .B(G225), .Z(G308) );
  INV_X1 U1012 ( .A(G108), .ZN(G238) );
  INV_X1 U1013 ( .A(G96), .ZN(G221) );
  INV_X1 U1014 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1015 ( .A1(n912), .A2(n911), .ZN(G325) );
  INV_X1 U1016 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U1017 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n1025) );
  XOR2_X1 U1018 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n935) );
  XNOR2_X1 U1019 ( .A(G20), .B(n913), .ZN(n917) );
  XNOR2_X1 U1020 ( .A(G1981), .B(G6), .ZN(n915) );
  XNOR2_X1 U1021 ( .A(G19), .B(G1341), .ZN(n914) );
  NOR2_X1 U1022 ( .A1(n915), .A2(n914), .ZN(n916) );
  NAND2_X1 U1023 ( .A1(n917), .A2(n916), .ZN(n920) );
  XOR2_X1 U1024 ( .A(KEYINPUT59), .B(G1348), .Z(n918) );
  XNOR2_X1 U1025 ( .A(G4), .B(n918), .ZN(n919) );
  NOR2_X1 U1026 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1027 ( .A(KEYINPUT60), .B(n921), .Z(n923) );
  XNOR2_X1 U1028 ( .A(G1961), .B(G5), .ZN(n922) );
  NOR2_X1 U1029 ( .A1(n923), .A2(n922), .ZN(n933) );
  XNOR2_X1 U1030 ( .A(G1976), .B(G23), .ZN(n925) );
  XNOR2_X1 U1031 ( .A(G22), .B(G1971), .ZN(n924) );
  NOR2_X1 U1032 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1033 ( .A(KEYINPUT124), .B(n926), .Z(n928) );
  XNOR2_X1 U1034 ( .A(G1986), .B(G24), .ZN(n927) );
  NOR2_X1 U1035 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1036 ( .A(KEYINPUT58), .B(n929), .Z(n931) );
  XNOR2_X1 U1037 ( .A(G1966), .B(G21), .ZN(n930) );
  NOR2_X1 U1038 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1039 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1040 ( .A(n935), .B(n934), .ZN(n936) );
  NOR2_X1 U1041 ( .A1(G16), .A2(n936), .ZN(n1023) );
  XNOR2_X1 U1042 ( .A(KEYINPUT56), .B(G16), .ZN(n967) );
  XNOR2_X1 U1043 ( .A(G1348), .B(n937), .ZN(n938) );
  XNOR2_X1 U1044 ( .A(n938), .B(KEYINPUT119), .ZN(n943) );
  XNOR2_X1 U1045 ( .A(G171), .B(n939), .ZN(n940) );
  NOR2_X1 U1046 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1047 ( .A1(n943), .A2(n942), .ZN(n947) );
  XOR2_X1 U1048 ( .A(G1956), .B(n944), .Z(n945) );
  XNOR2_X1 U1049 ( .A(KEYINPUT120), .B(n945), .ZN(n946) );
  NOR2_X1 U1050 ( .A1(n947), .A2(n946), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(G1966), .B(G168), .ZN(n948) );
  XNOR2_X1 U1052 ( .A(n948), .B(KEYINPUT117), .ZN(n950) );
  NOR2_X1 U1053 ( .A1(n950), .A2(n949), .ZN(n952) );
  XOR2_X1 U1054 ( .A(KEYINPUT118), .B(KEYINPUT57), .Z(n951) );
  XNOR2_X1 U1055 ( .A(n952), .B(n951), .ZN(n953) );
  NAND2_X1 U1056 ( .A1(n954), .A2(n953), .ZN(n957) );
  XNOR2_X1 U1057 ( .A(G1341), .B(n955), .ZN(n956) );
  NOR2_X1 U1058 ( .A1(n957), .A2(n956), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(G1971), .B(G303), .ZN(n958) );
  XNOR2_X1 U1060 ( .A(n958), .B(KEYINPUT121), .ZN(n960) );
  NAND2_X1 U1061 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1062 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1063 ( .A(n963), .B(KEYINPUT122), .ZN(n964) );
  NAND2_X1 U1064 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1065 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1066 ( .A(n968), .B(KEYINPUT123), .ZN(n1020) );
  XOR2_X1 U1067 ( .A(G2090), .B(G35), .Z(n971) );
  XOR2_X1 U1068 ( .A(G34), .B(KEYINPUT54), .Z(n969) );
  XNOR2_X1 U1069 ( .A(n969), .B(G2084), .ZN(n970) );
  NAND2_X1 U1070 ( .A1(n971), .A2(n970), .ZN(n987) );
  XOR2_X1 U1071 ( .A(n972), .B(G27), .Z(n974) );
  XNOR2_X1 U1072 ( .A(G2072), .B(G33), .ZN(n973) );
  NOR2_X1 U1073 ( .A1(n974), .A2(n973), .ZN(n983) );
  XOR2_X1 U1074 ( .A(G2067), .B(G26), .Z(n977) );
  INV_X1 U1075 ( .A(G1996), .ZN(n975) );
  XNOR2_X1 U1076 ( .A(n975), .B(G32), .ZN(n976) );
  NAND2_X1 U1077 ( .A1(n977), .A2(n976), .ZN(n981) );
  XOR2_X1 U1078 ( .A(G1991), .B(G25), .Z(n978) );
  NAND2_X1 U1079 ( .A1(n978), .A2(G28), .ZN(n979) );
  XNOR2_X1 U1080 ( .A(n979), .B(KEYINPUT114), .ZN(n980) );
  NOR2_X1 U1081 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1082 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1083 ( .A(KEYINPUT53), .B(n984), .ZN(n985) );
  XNOR2_X1 U1084 ( .A(n985), .B(KEYINPUT115), .ZN(n986) );
  NOR2_X1 U1085 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1086 ( .A(KEYINPUT55), .B(n988), .Z(n989) );
  NOR2_X1 U1087 ( .A1(G29), .A2(n989), .ZN(n990) );
  XOR2_X1 U1088 ( .A(KEYINPUT116), .B(n990), .Z(n1018) );
  XOR2_X1 U1089 ( .A(G2072), .B(n991), .Z(n993) );
  XOR2_X1 U1090 ( .A(G164), .B(G2078), .Z(n992) );
  NOR2_X1 U1091 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1092 ( .A(KEYINPUT50), .B(n994), .Z(n1012) );
  XNOR2_X1 U1093 ( .A(G160), .B(G2084), .ZN(n996) );
  NAND2_X1 U1094 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1095 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1096 ( .A1(n1000), .A2(n999), .ZN(n1005) );
  XOR2_X1 U1097 ( .A(G2090), .B(G162), .Z(n1001) );
  NOR2_X1 U1098 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1099 ( .A(n1003), .B(KEYINPUT51), .ZN(n1004) );
  NOR2_X1 U1100 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  NAND2_X1 U1101 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1102 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1103 ( .A(KEYINPUT113), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1104 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1105 ( .A(KEYINPUT52), .B(n1013), .ZN(n1015) );
  INV_X1 U1106 ( .A(KEYINPUT55), .ZN(n1014) );
  NAND2_X1 U1107 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1108 ( .A1(n1016), .A2(G29), .ZN(n1017) );
  NAND2_X1 U1109 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1111 ( .A1(n1021), .A2(G11), .ZN(n1022) );
  NOR2_X1 U1112 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1113 ( .A(n1025), .B(n1024), .ZN(G311) );
  XNOR2_X1 U1114 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

