//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 0 0 0 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n841, new_n842,
    new_n843, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949;
  INV_X1    g000(.A(G169gat), .ZN(new_n202));
  INV_X1    g001(.A(G176gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT65), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT65), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G169gat), .B2(G176gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT26), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  AND2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT69), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT69), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n212), .A2(new_n216), .A3(new_n213), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT27), .B(G183gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n219), .A2(G190gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n221));
  AND3_X1   g020(.A1(new_n218), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n221), .B1(new_n218), .B2(new_n220), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n215), .A2(new_n217), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n213), .ZN(new_n226));
  AND2_X1   g025(.A1(KEYINPUT66), .A2(KEYINPUT24), .ZN(new_n227));
  NOR2_X1   g026(.A1(KEYINPUT66), .A2(KEYINPUT24), .ZN(new_n228));
  NOR3_X1   g027(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  OR2_X1    g028(.A1(G183gat), .A2(G190gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT67), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT23), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT64), .ZN(new_n235));
  NOR2_X1   g034(.A1(G169gat), .A2(G176gat), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n235), .B1(new_n236), .B2(KEYINPUT23), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT23), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n238), .B(KEYINPUT64), .C1(G169gat), .C2(G176gat), .ZN(new_n239));
  AOI22_X1  g038(.A1(new_n237), .A2(new_n239), .B1(G169gat), .B2(G176gat), .ZN(new_n240));
  OR2_X1    g039(.A1(KEYINPUT66), .A2(KEYINPUT24), .ZN(new_n241));
  NAND2_X1  g040(.A1(KEYINPUT66), .A2(KEYINPUT24), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n241), .A2(new_n213), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n243), .A2(new_n244), .A3(new_n230), .A4(new_n231), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n233), .A2(new_n234), .A3(new_n240), .A4(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(KEYINPUT25), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n237), .A2(new_n239), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n210), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT25), .B1(new_n236), .B2(KEYINPUT23), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n226), .A2(KEYINPUT24), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n250), .B1(new_n251), .B2(new_n232), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n225), .A2(new_n247), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G226gat), .A2(G233gat), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G197gat), .B(G204gat), .ZN(new_n259));
  INV_X1    g058(.A(G211gat), .ZN(new_n260));
  INV_X1    g059(.A(G218gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n259), .B1(KEYINPUT22), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G211gat), .B(G218gat), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n264), .B(new_n259), .C1(KEYINPUT22), .C2(new_n262), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n258), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT29), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n257), .B1(new_n255), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(KEYINPUT76), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n268), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n273), .B1(new_n255), .B2(new_n257), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT76), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n253), .B1(new_n246), .B2(KEYINPUT25), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT29), .B1(new_n276), .B2(new_n225), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n274), .B(new_n275), .C1(new_n257), .C2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n256), .B1(new_n276), .B2(new_n225), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n273), .B1(new_n271), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n272), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G8gat), .B(G36gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(G64gat), .B(G92gat), .ZN(new_n283));
  XOR2_X1   g082(.A(new_n282), .B(new_n283), .Z(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n272), .A2(new_n284), .A3(new_n278), .A4(new_n280), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n286), .A2(KEYINPUT30), .A3(new_n287), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n258), .B(new_n268), .C1(new_n257), .C2(new_n277), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n258), .B1(new_n257), .B2(new_n277), .ZN(new_n290));
  AOI22_X1  g089(.A1(new_n289), .A2(KEYINPUT76), .B1(new_n290), .B2(new_n273), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT30), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n291), .A2(new_n292), .A3(new_n284), .A4(new_n278), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n288), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT77), .B(G162gat), .ZN(new_n295));
  INV_X1    g094(.A(G155gat), .ZN(new_n296));
  OAI21_X1  g095(.A(KEYINPUT2), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OR2_X1    g096(.A1(G141gat), .A2(G148gat), .ZN(new_n298));
  INV_X1    g097(.A(G162gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G155gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n296), .A2(G162gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(G141gat), .A2(G148gat), .ZN(new_n302));
  AND4_X1   g101(.A1(new_n298), .A2(new_n300), .A3(new_n301), .A4(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT2), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n298), .A2(new_n304), .A3(new_n302), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n300), .A2(new_n301), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n297), .A2(new_n303), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AND2_X1   g106(.A1(G113gat), .A2(G120gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(G113gat), .A2(G120gat), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT70), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G113gat), .ZN(new_n311));
  INV_X1    g110(.A(G120gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT70), .ZN(new_n314));
  NAND2_X1  g113(.A1(G113gat), .A2(G120gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT1), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n310), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(G134gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G127gat), .ZN(new_n320));
  INV_X1    g119(.A(G127gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G134gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n320), .A2(new_n322), .A3(new_n317), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT71), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n327), .B1(new_n308), .B2(new_n309), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n313), .A2(KEYINPUT71), .A3(new_n315), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n326), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n307), .A2(new_n324), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT4), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT80), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n308), .A2(new_n309), .A3(new_n327), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n334), .A2(new_n325), .ZN(new_n335));
  AOI22_X1  g134(.A1(new_n328), .A2(new_n335), .B1(new_n318), .B2(new_n323), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT4), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n336), .A2(new_n337), .A3(new_n307), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n332), .A2(new_n333), .A3(new_n338), .ZN(new_n339));
  AND2_X1   g138(.A1(new_n298), .A2(new_n302), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n300), .A2(new_n301), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n299), .A2(KEYINPUT77), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT77), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(G162gat), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n296), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n340), .B(new_n341), .C1(new_n345), .C2(new_n304), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n305), .A2(new_n306), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT3), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n324), .A2(new_n330), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n307), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n349), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n331), .A2(KEYINPUT80), .A3(KEYINPUT4), .ZN(new_n354));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n356), .A2(KEYINPUT5), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n339), .A2(new_n353), .A3(new_n354), .A4(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT81), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n350), .A2(new_n348), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n324), .A2(new_n330), .B1(new_n346), .B2(new_n347), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n356), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT78), .ZN(new_n364));
  NOR3_X1   g163(.A1(new_n350), .A2(new_n348), .A3(KEYINPUT4), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n337), .B1(new_n336), .B2(new_n307), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n353), .B(new_n355), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT78), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n368), .B(new_n356), .C1(new_n361), .C2(new_n362), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n364), .A2(new_n367), .A3(KEYINPUT5), .A4(new_n369), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n354), .A2(new_n353), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n371), .A2(KEYINPUT81), .A3(new_n339), .A4(new_n357), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n360), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  XOR2_X1   g172(.A(G1gat), .B(G29gat), .Z(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G57gat), .B(G85gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT6), .ZN(new_n380));
  INV_X1    g179(.A(new_n378), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n360), .A2(new_n370), .A3(new_n381), .A4(new_n372), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n379), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n373), .A2(KEYINPUT6), .A3(new_n378), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n294), .A2(new_n385), .ZN(new_n386));
  AND2_X1   g185(.A1(G228gat), .A2(G233gat), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT29), .B1(new_n266), .B2(new_n267), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n348), .B1(new_n388), .B2(KEYINPUT3), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n387), .B1(new_n389), .B2(KEYINPUT82), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT29), .B1(new_n307), .B2(new_n351), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n389), .B1(new_n391), .B2(new_n268), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  OAI221_X1 g192(.A(new_n389), .B1(KEYINPUT82), .B2(new_n387), .C1(new_n391), .C2(new_n268), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT83), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(G22gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(G78gat), .B(G106gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT31), .B(G50gat), .ZN(new_n400));
  XOR2_X1   g199(.A(new_n399), .B(new_n400), .Z(new_n401));
  NAND3_X1  g200(.A1(new_n397), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n395), .A2(new_n396), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT83), .B1(new_n393), .B2(new_n394), .ZN(new_n404));
  INV_X1    g203(.A(new_n401), .ZN(new_n405));
  OAI21_X1  g204(.A(G22gat), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n402), .A2(new_n403), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n403), .B1(new_n402), .B2(new_n406), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n386), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT36), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT73), .ZN(new_n413));
  NAND2_X1  g212(.A1(G227gat), .A2(G233gat), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n336), .B1(new_n276), .B2(new_n225), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT72), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n276), .A2(new_n225), .A3(new_n336), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n276), .A2(KEYINPUT72), .A3(new_n225), .A4(new_n336), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n414), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT32), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n413), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n417), .A2(new_n416), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n255), .A2(new_n350), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n423), .A2(new_n419), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n414), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n427), .A2(KEYINPUT73), .A3(KEYINPUT32), .ZN(new_n428));
  XNOR2_X1  g227(.A(G15gat), .B(G43gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(KEYINPUT74), .ZN(new_n430));
  XOR2_X1   g229(.A(G71gat), .B(G99gat), .Z(new_n431));
  XNOR2_X1  g230(.A(new_n430), .B(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT33), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n433), .B1(new_n427), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n422), .A2(new_n428), .A3(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n423), .A2(new_n414), .A3(new_n424), .A4(new_n419), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT75), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT34), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n439), .B1(new_n437), .B2(new_n438), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n427), .B(KEYINPUT32), .C1(new_n434), .C2(new_n433), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n436), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n442), .B1(new_n436), .B2(new_n443), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n412), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n436), .A2(new_n443), .ZN(new_n447));
  INV_X1    g246(.A(new_n442), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n436), .A2(new_n442), .A3(new_n443), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(KEYINPUT36), .A3(new_n450), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n411), .A2(new_n446), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n294), .ZN(new_n453));
  XNOR2_X1  g252(.A(KEYINPUT84), .B(KEYINPUT39), .ZN(new_n454));
  INV_X1    g253(.A(new_n339), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n354), .A2(new_n353), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n356), .B(new_n454), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n381), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n355), .B1(new_n371), .B2(new_n339), .ZN(new_n459));
  OR2_X1    g258(.A1(new_n361), .A2(new_n362), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT39), .B1(new_n460), .B2(new_n356), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT85), .B1(new_n458), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT40), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n379), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n463), .A2(KEYINPUT40), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n410), .B1(new_n453), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT37), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n272), .A2(new_n469), .A3(new_n278), .A4(new_n280), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT87), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n291), .A2(KEYINPUT87), .A3(new_n469), .A4(new_n278), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT38), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n285), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT86), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n280), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n290), .A2(KEYINPUT86), .A3(new_n273), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(new_n289), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n476), .B1(new_n480), .B2(KEYINPUT37), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n474), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT88), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n474), .A2(KEYINPUT88), .A3(new_n481), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n383), .A2(new_n384), .A3(new_n287), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT89), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n284), .B1(new_n281), .B2(KEYINPUT37), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n488), .A2(new_n489), .B1(new_n472), .B2(new_n473), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n489), .A2(new_n488), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n475), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n468), .B1(new_n487), .B2(new_n492), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n288), .A2(new_n293), .B1(new_n384), .B2(new_n383), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n494), .B(new_n409), .C1(new_n444), .C2(new_n445), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT35), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n449), .A2(new_n450), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT35), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n497), .A2(new_n498), .A3(new_n409), .A4(new_n494), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n452), .A2(new_n493), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  XOR2_X1   g299(.A(G43gat), .B(G50gat), .Z(new_n501));
  INV_X1    g300(.A(KEYINPUT92), .ZN(new_n502));
  OR2_X1    g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(G29gat), .A2(G36gat), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  NOR3_X1   g305(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n501), .A2(new_n502), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n503), .A2(KEYINPUT15), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n507), .A2(KEYINPUT95), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n507), .A2(KEYINPUT95), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n505), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT96), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n503), .A2(KEYINPUT15), .A3(new_n509), .ZN(new_n516));
  XOR2_X1   g315(.A(KEYINPUT93), .B(KEYINPUT15), .Z(new_n517));
  INV_X1    g316(.A(KEYINPUT94), .ZN(new_n518));
  INV_X1    g317(.A(G50gat), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n518), .B1(new_n519), .B2(G43gat), .ZN(new_n520));
  INV_X1    g319(.A(G43gat), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n520), .B1(new_n521), .B2(G50gat), .ZN(new_n522));
  NOR3_X1   g321(.A1(new_n518), .A2(new_n519), .A3(G43gat), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n517), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n504), .B(KEYINPUT97), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n516), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n510), .B1(new_n515), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT17), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G15gat), .B(G22gat), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT16), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n530), .B1(new_n531), .B2(G1gat), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n532), .B1(G1gat), .B2(new_n530), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n533), .B(G8gat), .Z(new_n534));
  OAI211_X1 g333(.A(KEYINPUT17), .B(new_n510), .C1(new_n515), .C2(new_n526), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n529), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(G229gat), .A2(G233gat), .ZN(new_n537));
  INV_X1    g336(.A(new_n534), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n527), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT18), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n536), .A2(KEYINPUT18), .A3(new_n537), .A4(new_n539), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n537), .B(KEYINPUT13), .Z(new_n544));
  INV_X1    g343(.A(new_n539), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n538), .A2(new_n527), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n542), .A2(new_n543), .A3(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G113gat), .B(G141gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G169gat), .B(G197gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(KEYINPUT91), .B(KEYINPUT12), .Z(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n548), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n542), .A2(new_n555), .A3(new_n543), .A4(new_n547), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n500), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n385), .ZN(new_n562));
  NAND2_X1  g361(.A1(G85gat), .A2(G92gat), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT7), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(KEYINPUT101), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT8), .ZN(new_n566));
  AND2_X1   g365(.A1(G99gat), .A2(G106gat), .ZN(new_n567));
  OAI221_X1 g366(.A(new_n565), .B1(G85gat), .B2(G92gat), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT7), .B1(new_n563), .B2(KEYINPUT101), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n569), .B1(KEYINPUT101), .B2(new_n563), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(G99gat), .A2(G106gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n573), .B1(new_n568), .B2(new_n570), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n529), .A2(new_n535), .A3(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n577), .ZN(new_n579));
  AND2_X1   g378(.A1(G232gat), .A2(G233gat), .ZN(new_n580));
  AOI22_X1  g379(.A1(new_n527), .A2(new_n579), .B1(KEYINPUT41), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G190gat), .B(G218gat), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT102), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G134gat), .B(G162gat), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n582), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n587), .B1(new_n582), .B2(new_n585), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n583), .A2(new_n584), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n580), .A2(KEYINPUT41), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n590), .B(new_n591), .Z(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  OR3_X1    g392(.A1(new_n588), .A2(new_n589), .A3(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n593), .B1(new_n588), .B2(new_n589), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AND2_X1   g395(.A1(G71gat), .A2(G78gat), .ZN(new_n597));
  NOR2_X1   g396(.A1(G71gat), .A2(G78gat), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AND2_X1   g398(.A1(G57gat), .A2(G64gat), .ZN(new_n600));
  OAI21_X1  g399(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n597), .B1(KEYINPUT9), .B2(new_n598), .ZN(new_n603));
  NAND2_X1  g402(.A1(KEYINPUT98), .A2(G57gat), .ZN(new_n604));
  INV_X1    g403(.A(G64gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n602), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n608), .A2(KEYINPUT21), .ZN(new_n609));
  AND2_X1   g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(new_n321), .ZN(new_n612));
  XOR2_X1   g411(.A(G183gat), .B(G211gat), .Z(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n611), .B(G127gat), .ZN(new_n615));
  INV_X1    g414(.A(new_n613), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n608), .A2(KEYINPUT21), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n534), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(new_n296), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n622), .A2(new_n625), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n618), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n628), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n630), .A2(new_n614), .A3(new_n617), .A4(new_n626), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT104), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n579), .A2(KEYINPUT10), .A3(new_n608), .ZN(new_n634));
  OAI21_X1  g433(.A(KEYINPUT103), .B1(new_n568), .B2(new_n570), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n607), .B1(new_n635), .B2(new_n573), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n636), .B1(new_n573), .B2(new_n635), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n575), .A2(new_n607), .A3(new_n576), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OAI211_X1 g438(.A(new_n633), .B(new_n634), .C1(new_n639), .C2(KEYINPUT10), .ZN(new_n640));
  AOI21_X1  g439(.A(KEYINPUT10), .B1(new_n637), .B2(new_n638), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n579), .A2(KEYINPUT10), .A3(new_n608), .ZN(new_n642));
  OAI21_X1  g441(.A(KEYINPUT104), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(G230gat), .A2(G233gat), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n644), .B(KEYINPUT105), .Z(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n640), .A2(new_n643), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G120gat), .B(G148gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(G176gat), .B(G204gat), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n648), .B(new_n649), .Z(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n651), .B1(new_n639), .B2(new_n645), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n646), .B1(new_n641), .B2(new_n642), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n645), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n650), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n596), .A2(new_n632), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n561), .A2(new_n562), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(G1gat), .ZN(G1324gat));
  NOR3_X1   g461(.A1(new_n500), .A2(new_n560), .A3(new_n659), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT16), .B(G8gat), .Z(new_n664));
  NAND3_X1  g463(.A1(new_n663), .A2(new_n453), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n663), .ZN(new_n666));
  OAI21_X1  g465(.A(G8gat), .B1(new_n666), .B2(new_n294), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(new_n665), .ZN(new_n668));
  MUX2_X1   g467(.A(new_n665), .B(new_n668), .S(KEYINPUT42), .Z(G1325gat));
  AND2_X1   g468(.A1(new_n446), .A2(new_n451), .ZN(new_n670));
  OAI21_X1  g469(.A(G15gat), .B1(new_n666), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n497), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n672), .A2(new_n659), .A3(G15gat), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n561), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n671), .A2(new_n674), .ZN(G1326gat));
  NAND2_X1  g474(.A1(new_n663), .A2(new_n410), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT106), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT43), .B(G22gat), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n677), .B(new_n678), .Z(G1327gat));
  NOR2_X1   g478(.A1(new_n500), .A2(new_n596), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n680), .A2(KEYINPUT44), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(KEYINPUT44), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n632), .B(KEYINPUT108), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT107), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n559), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n557), .A2(KEYINPUT107), .A3(new_n558), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n658), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n685), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n683), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(G29gat), .B1(new_n693), .B2(new_n385), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n596), .A2(new_n691), .A3(new_n632), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n561), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(G29gat), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n696), .A2(new_n697), .A3(new_n562), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT45), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n694), .A2(new_n699), .ZN(G1328gat));
  OAI21_X1  g499(.A(G36gat), .B1(new_n693), .B2(new_n294), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT109), .ZN(new_n702));
  AOI21_X1  g501(.A(G36gat), .B1(new_n702), .B2(KEYINPUT46), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n696), .A2(new_n453), .A3(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n702), .A2(KEYINPUT46), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n701), .A2(new_n706), .ZN(G1329gat));
  NAND3_X1  g506(.A1(new_n696), .A2(new_n521), .A3(new_n497), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT110), .ZN(new_n709));
  INV_X1    g508(.A(new_n670), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n681), .A2(new_n710), .A3(new_n682), .A4(new_n692), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n711), .A2(G43gat), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT47), .ZN(new_n713));
  OR3_X1    g512(.A1(new_n709), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n713), .B1(new_n709), .B2(new_n712), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(G1330gat));
  NAND4_X1  g515(.A1(new_n681), .A2(new_n410), .A3(new_n682), .A4(new_n692), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(G50gat), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n696), .A2(new_n519), .A3(new_n410), .ZN(new_n719));
  AOI21_X1  g518(.A(KEYINPUT111), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT48), .Z(G1331gat));
  NAND3_X1  g520(.A1(new_n596), .A2(new_n632), .A3(new_n691), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n500), .A2(new_n689), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n562), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n453), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n726), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n727));
  XOR2_X1   g526(.A(KEYINPUT49), .B(G64gat), .Z(new_n728));
  OAI21_X1  g527(.A(new_n727), .B1(new_n726), .B2(new_n728), .ZN(G1333gat));
  NAND2_X1  g528(.A1(new_n723), .A2(new_n710), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n672), .A2(G71gat), .ZN(new_n731));
  AOI22_X1  g530(.A1(new_n730), .A2(G71gat), .B1(new_n723), .B2(new_n731), .ZN(new_n732));
  XOR2_X1   g531(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(G1334gat));
  NAND2_X1  g533(.A1(new_n723), .A2(new_n410), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G78gat), .ZN(G1335gat));
  INV_X1    g535(.A(G85gat), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n689), .A2(new_n632), .A3(new_n658), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n683), .A2(new_n562), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n737), .B1(new_n739), .B2(KEYINPUT113), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n740), .B1(KEYINPUT113), .B2(new_n739), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT114), .B1(new_n500), .B2(new_n596), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT114), .ZN(new_n743));
  INV_X1    g542(.A(new_n596), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n411), .A2(new_n446), .A3(new_n451), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n490), .A2(new_n491), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT38), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n747), .A2(new_n485), .A3(new_n484), .A4(new_n486), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n745), .B1(new_n748), .B2(new_n468), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n496), .A2(new_n499), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n743), .B(new_n744), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n689), .A2(new_n632), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n742), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n742), .A2(new_n751), .A3(KEYINPUT51), .A4(new_n752), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n691), .A2(new_n562), .A3(new_n737), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n741), .B1(new_n758), .B2(new_n759), .ZN(G1336gat));
  INV_X1    g559(.A(new_n758), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n294), .A2(G92gat), .A3(new_n658), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n681), .A2(new_n453), .A3(new_n682), .A4(new_n738), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n764), .A2(G92gat), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n765), .A2(KEYINPUT52), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n753), .A2(KEYINPUT115), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT115), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n742), .A2(new_n751), .A3(new_n769), .A4(new_n752), .ZN(new_n770));
  AND4_X1   g569(.A1(KEYINPUT116), .A2(new_n768), .A3(new_n754), .A4(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT116), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT51), .B1(new_n753), .B2(KEYINPUT115), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n773), .B1(new_n774), .B2(new_n770), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n765), .B1(new_n776), .B2(new_n762), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n767), .B1(new_n777), .B2(new_n778), .ZN(G1337gat));
  NAND3_X1  g578(.A1(new_n683), .A2(new_n710), .A3(new_n738), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(G99gat), .ZN(new_n781));
  OR3_X1    g580(.A1(new_n672), .A2(G99gat), .A3(new_n658), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n781), .B1(new_n758), .B2(new_n782), .ZN(G1338gat));
  NOR3_X1   g582(.A1(new_n409), .A2(new_n658), .A3(G106gat), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n761), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n681), .A2(new_n410), .A3(new_n682), .A4(new_n738), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n786), .A2(G106gat), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(KEYINPUT53), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n787), .B1(new_n776), .B2(new_n784), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(G1339gat));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n645), .B(new_n634), .C1(new_n639), .C2(KEYINPUT10), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT54), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n643), .A2(new_n646), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n795), .B1(new_n796), .B2(new_n640), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n651), .B1(new_n655), .B2(KEYINPUT54), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n793), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n795), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n798), .B1(new_n800), .B2(new_n647), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT55), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n799), .A2(new_n802), .A3(new_n653), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n803), .B1(new_n687), .B2(new_n688), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n537), .B1(new_n536), .B2(new_n539), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n545), .A2(new_n546), .A3(new_n544), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n553), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n558), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n658), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n596), .B1(new_n804), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n653), .B1(new_n801), .B2(KEYINPUT55), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n797), .A2(new_n793), .A3(new_n798), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n744), .A2(new_n813), .A3(new_n558), .A4(new_n807), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n685), .B1(new_n810), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n689), .A2(new_n659), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n672), .A2(new_n410), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n453), .A2(new_n385), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(G113gat), .B1(new_n822), .B2(new_n560), .ZN(new_n823));
  INV_X1    g622(.A(new_n688), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT107), .B1(new_n557), .B2(new_n558), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n813), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n809), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n744), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n814), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n684), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n816), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n385), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n818), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(new_n453), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(new_n311), .A3(new_n689), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n823), .A2(new_n835), .ZN(new_n836));
  XOR2_X1   g635(.A(new_n836), .B(KEYINPUT117), .Z(G1340gat));
  AOI21_X1  g636(.A(G120gat), .B1(new_n834), .B2(new_n691), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n822), .A2(new_n312), .A3(new_n658), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(G1341gat));
  NOR3_X1   g639(.A1(new_n822), .A2(new_n321), .A3(new_n684), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT118), .ZN(new_n842));
  AOI21_X1  g641(.A(G127gat), .B1(new_n834), .B2(new_n632), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(new_n843), .ZN(G1342gat));
  OR4_X1    g643(.A1(G134gat), .A2(new_n833), .A3(new_n453), .A4(new_n596), .ZN(new_n845));
  OR2_X1    g644(.A1(new_n845), .A2(KEYINPUT56), .ZN(new_n846));
  OAI21_X1  g645(.A(G134gat), .B1(new_n822), .B2(new_n596), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(KEYINPUT56), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(G1343gat));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n850), .B(new_n410), .C1(new_n815), .C2(new_n816), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n809), .B1(new_n813), .B2(new_n559), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n814), .B1(new_n852), .B2(new_n744), .ZN(new_n853));
  INV_X1    g652(.A(new_n632), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n816), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(KEYINPUT57), .B1(new_n855), .B2(new_n409), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n670), .A2(new_n821), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n851), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(G141gat), .B1(new_n858), .B2(new_n690), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n830), .A2(new_n831), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n670), .A2(new_n410), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(new_n453), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n560), .A2(G141gat), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n860), .A2(new_n862), .A3(new_n562), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(KEYINPUT58), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n851), .A2(new_n856), .A3(new_n559), .A4(new_n857), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT58), .B1(new_n867), .B2(G141gat), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n864), .A2(KEYINPUT119), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT119), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n832), .A2(new_n870), .A3(new_n862), .A4(new_n863), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n868), .A2(new_n872), .A3(KEYINPUT120), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT120), .B1(new_n868), .B2(new_n872), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n866), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT121), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n877), .B(new_n866), .C1(new_n873), .C2(new_n874), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n878), .ZN(G1344gat));
  AND2_X1   g678(.A1(new_n832), .A2(new_n862), .ZN(new_n880));
  INV_X1    g679(.A(G148gat), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n880), .A2(new_n881), .A3(new_n691), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT57), .B1(new_n817), .B2(new_n409), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n803), .A2(new_n596), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n808), .B1(new_n885), .B2(KEYINPUT122), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n886), .B1(KEYINPUT122), .B2(new_n885), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n852), .A2(new_n744), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n632), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n659), .A2(new_n559), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n850), .B(new_n410), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n884), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(new_n691), .A3(new_n857), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n883), .B1(new_n893), .B2(G148gat), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n858), .A2(new_n658), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n895), .A2(KEYINPUT59), .A3(new_n881), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n882), .B1(new_n894), .B2(new_n896), .ZN(G1345gat));
  OAI21_X1  g696(.A(G155gat), .B1(new_n858), .B2(new_n684), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n880), .A2(new_n296), .A3(new_n632), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1346gat));
  NAND3_X1  g699(.A1(new_n880), .A2(new_n295), .A3(new_n744), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n858), .A2(new_n596), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n902), .B2(new_n295), .ZN(G1347gat));
  NOR2_X1   g702(.A1(new_n562), .A2(new_n294), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n820), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(G169gat), .B1(new_n905), .B2(new_n560), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT123), .ZN(new_n907));
  NOR4_X1   g706(.A1(new_n817), .A2(new_n562), .A3(new_n294), .A4(new_n819), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n202), .A3(new_n689), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(G1348gat));
  AOI21_X1  g709(.A(G176gat), .B1(new_n908), .B2(new_n691), .ZN(new_n911));
  XOR2_X1   g710(.A(new_n911), .B(KEYINPUT124), .Z(new_n912));
  NOR3_X1   g711(.A1(new_n905), .A2(new_n203), .A3(new_n658), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n912), .A2(new_n913), .ZN(G1349gat));
  OAI21_X1  g713(.A(G183gat), .B1(new_n905), .B2(new_n684), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT125), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n908), .A2(new_n218), .A3(new_n632), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g718(.A(G190gat), .B1(new_n905), .B2(new_n596), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT61), .ZN(new_n921));
  INV_X1    g720(.A(G190gat), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n908), .A2(new_n922), .A3(new_n744), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(G1351gat));
  AND2_X1   g723(.A1(new_n670), .A2(new_n904), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n892), .A2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(G197gat), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n926), .A2(new_n927), .A3(new_n560), .ZN(new_n928));
  NOR4_X1   g727(.A1(new_n817), .A2(new_n562), .A3(new_n294), .A4(new_n861), .ZN(new_n929));
  AOI21_X1  g728(.A(G197gat), .B1(new_n929), .B2(new_n689), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n928), .A2(new_n930), .ZN(G1352gat));
  INV_X1    g730(.A(G204gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n929), .A2(new_n932), .A3(new_n691), .ZN(new_n933));
  XOR2_X1   g732(.A(new_n933), .B(KEYINPUT62), .Z(new_n934));
  OAI21_X1  g733(.A(G204gat), .B1(new_n926), .B2(new_n658), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1353gat));
  NAND3_X1  g735(.A1(new_n929), .A2(new_n260), .A3(new_n632), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n892), .A2(new_n632), .A3(new_n925), .ZN(new_n938));
  AND4_X1   g737(.A1(KEYINPUT126), .A2(new_n938), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n939));
  OAI21_X1  g738(.A(G211gat), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  AOI22_X1  g740(.A1(new_n938), .A2(new_n941), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n937), .B1(new_n939), .B2(new_n942), .ZN(G1354gat));
  OAI21_X1  g742(.A(G218gat), .B1(new_n926), .B2(new_n596), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n929), .A2(new_n261), .A3(new_n744), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(KEYINPUT127), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT127), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n944), .A2(new_n948), .A3(new_n945), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n949), .ZN(G1355gat));
endmodule


