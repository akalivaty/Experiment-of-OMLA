//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 0 1 0 0 1 0 0 0 0 0 0 0 1 1 1 1 1 0 1 1 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n844, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT16), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(new_n204), .B2(G1gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G1gat), .B2(new_n203), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(G8gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(G29gat), .A2(G36gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n209), .A2(KEYINPUT90), .ZN(new_n210));
  XOR2_X1   g009(.A(G43gat), .B(G50gat), .Z(new_n211));
  INV_X1    g010(.A(KEYINPUT15), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(G29gat), .A2(G36gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n214), .B(KEYINPUT14), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G43gat), .B(G50gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT15), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n209), .A2(KEYINPUT90), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n213), .A2(new_n216), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  OAI211_X1 g019(.A(KEYINPUT15), .B(new_n217), .C1(new_n215), .C2(new_n209), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n207), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT17), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n222), .B(new_n224), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n202), .B(new_n223), .C1(new_n225), .C2(new_n207), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT18), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT91), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n202), .B(KEYINPUT13), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n207), .A2(new_n222), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n229), .B1(new_n230), .B2(new_n223), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n231), .B1(new_n226), .B2(new_n227), .ZN(new_n232));
  INV_X1    g031(.A(new_n223), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n222), .B(KEYINPUT17), .ZN(new_n234));
  XOR2_X1   g033(.A(new_n206), .B(G8gat), .Z(new_n235));
  AOI21_X1  g034(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT91), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n236), .A2(new_n237), .A3(KEYINPUT18), .A4(new_n202), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n228), .A2(new_n232), .A3(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(G169gat), .B(G197gat), .Z(new_n240));
  XNOR2_X1  g039(.A(G113gat), .B(G141gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g041(.A(KEYINPUT89), .B(KEYINPUT11), .Z(new_n243));
  XNOR2_X1  g042(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(KEYINPUT12), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n239), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n228), .A2(new_n232), .A3(new_n238), .A4(new_n245), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  OR2_X1    g048(.A1(G155gat), .A2(G162gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(G155gat), .A2(G162gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT2), .ZN(new_n253));
  INV_X1    g052(.A(G148gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(G141gat), .ZN(new_n255));
  INV_X1    g054(.A(G141gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(G148gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n252), .B1(new_n253), .B2(new_n258), .ZN(new_n259));
  AND2_X1   g058(.A1(KEYINPUT74), .A2(G148gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(KEYINPUT74), .A2(G148gat), .ZN(new_n261));
  OAI21_X1  g060(.A(G141gat), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT75), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT73), .B(G141gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G148gat), .ZN(new_n266));
  OAI211_X1 g065(.A(KEYINPUT75), .B(G141gat), .C1(new_n260), .C2(new_n261), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n264), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n251), .B1(new_n250), .B2(KEYINPUT2), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n259), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G113gat), .B(G120gat), .ZN(new_n272));
  INV_X1    g071(.A(G127gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n273), .A2(G134gat), .ZN(new_n274));
  OAI22_X1  g073(.A1(new_n272), .A2(KEYINPUT1), .B1(KEYINPUT67), .B2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G127gat), .B(G134gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  OR3_X1    g076(.A1(new_n271), .A2(new_n277), .A3(KEYINPUT4), .ZN(new_n278));
  INV_X1    g077(.A(new_n277), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(new_n270), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT4), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n271), .A2(KEYINPUT3), .ZN(new_n282));
  AOI211_X1 g081(.A(KEYINPUT3), .B(new_n259), .C1(new_n268), .C2(new_n269), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n283), .A2(new_n279), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n278), .A2(new_n281), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G225gat), .A2(G233gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(KEYINPUT5), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n277), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT76), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n280), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n271), .A2(KEYINPUT76), .A3(new_n277), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n286), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n287), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(G1gat), .B(G29gat), .Z(new_n297));
  XNOR2_X1  g096(.A(KEYINPUT78), .B(KEYINPUT79), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G57gat), .B(G85gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT5), .B1(new_n285), .B2(new_n286), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n296), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT6), .ZN(new_n307));
  INV_X1    g106(.A(new_n303), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(new_n295), .B2(new_n304), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n306), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n296), .A2(KEYINPUT6), .A3(new_n303), .A4(new_n305), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(G226gat), .ZN(new_n313));
  INV_X1    g112(.A(G233gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT25), .ZN(new_n316));
  NAND2_X1  g115(.A1(G183gat), .A2(G190gat), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT24), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n320));
  INV_X1    g119(.A(G183gat), .ZN(new_n321));
  INV_X1    g120(.A(G190gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n319), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(G169gat), .ZN(new_n325));
  INV_X1    g124(.A(G176gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(new_n326), .A3(KEYINPUT23), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT64), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G169gat), .A2(G176gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(G169gat), .A2(G176gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n331), .A2(KEYINPUT64), .A3(KEYINPUT23), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n324), .A2(new_n329), .A3(new_n330), .A4(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n331), .A2(KEYINPUT23), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n316), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT65), .ZN(new_n336));
  INV_X1    g135(.A(new_n330), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT23), .ZN(new_n338));
  NOR3_X1   g137(.A1(new_n338), .A2(G169gat), .A3(G176gat), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n337), .B1(new_n339), .B2(KEYINPUT64), .ZN(new_n340));
  INV_X1    g139(.A(new_n334), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n340), .A2(new_n341), .A3(new_n324), .A4(new_n329), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT65), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n342), .A2(new_n343), .A3(new_n316), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n341), .A2(new_n324), .A3(KEYINPUT25), .A4(new_n327), .ZN(new_n345));
  XOR2_X1   g144(.A(new_n330), .B(KEYINPUT66), .Z(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n336), .A2(new_n344), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT26), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n331), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(new_n330), .A3(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT27), .B(G183gat), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(KEYINPUT28), .A3(new_n322), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT28), .B1(new_n354), .B2(new_n322), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n353), .B(new_n317), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n349), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT29), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n315), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n359), .A2(KEYINPUT71), .A3(new_n315), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT71), .B1(new_n359), .B2(new_n315), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n362), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G211gat), .B(G218gat), .ZN(new_n367));
  INV_X1    g166(.A(G211gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT70), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT70), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(G211gat), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n369), .A2(new_n371), .A3(G218gat), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT22), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G197gat), .B(G204gat), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n367), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n374), .A2(new_n375), .A3(new_n367), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n366), .A2(new_n379), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n374), .A2(new_n375), .A3(new_n367), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n381), .A2(new_n376), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n359), .A2(new_n315), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n362), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(G8gat), .B(G36gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(G64gat), .B(G92gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n385), .B(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n380), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n387), .B1(new_n380), .B2(new_n384), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT72), .ZN(new_n390));
  OAI21_X1  g189(.A(KEYINPUT30), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT71), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n383), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n361), .B1(new_n393), .B2(new_n363), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n384), .B1(new_n394), .B2(new_n382), .ZN(new_n395));
  INV_X1    g194(.A(new_n387), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT30), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(KEYINPUT72), .A3(new_n398), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n312), .A2(new_n388), .A3(new_n391), .A4(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT80), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT83), .ZN(new_n403));
  INV_X1    g202(.A(G228gat), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n404), .A2(new_n314), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n268), .A2(new_n269), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT3), .ZN(new_n407));
  INV_X1    g206(.A(new_n259), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n379), .B1(new_n409), .B2(new_n360), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n405), .B1(new_n410), .B2(KEYINPUT82), .ZN(new_n411));
  OAI211_X1 g210(.A(KEYINPUT82), .B(new_n382), .C1(new_n283), .C2(KEYINPUT29), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n360), .B1(new_n381), .B2(new_n376), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n407), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n271), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n403), .B1(new_n411), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n405), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n382), .B1(new_n283), .B2(KEYINPUT29), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT82), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n270), .B1(new_n413), .B2(new_n407), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n422), .B1(new_n410), .B2(KEYINPUT82), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n421), .A2(new_n423), .A3(KEYINPUT83), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n417), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(G22gat), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n405), .B1(new_n415), .B2(new_n419), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n425), .A2(KEYINPUT84), .A3(new_n426), .A4(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(G78gat), .B(G106gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(G50gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n432));
  XOR2_X1   g231(.A(new_n431), .B(new_n432), .Z(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n429), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n426), .B1(new_n425), .B2(new_n428), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n436), .A2(KEYINPUT84), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n427), .B1(new_n417), .B2(new_n424), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n426), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n435), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n411), .A2(new_n416), .A3(new_n403), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT83), .B1(new_n421), .B2(new_n423), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n428), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n444), .A2(KEYINPUT85), .A3(G22gat), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT85), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n446), .B1(new_n438), .B2(new_n426), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n445), .A2(new_n447), .A3(new_n433), .A4(new_n439), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT86), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI211_X1 g249(.A(G22gat), .B(new_n427), .C1(new_n417), .C2(new_n424), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n444), .A2(G22gat), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n451), .B1(new_n452), .B2(new_n446), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n434), .B1(new_n436), .B2(KEYINPUT85), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT86), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n441), .B1(new_n450), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT88), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n349), .A2(new_n277), .A3(new_n358), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n277), .B1(new_n349), .B2(new_n358), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(G227gat), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n461), .A2(new_n314), .ZN(new_n462));
  AND2_X1   g261(.A1(KEYINPUT69), .A2(KEYINPUT34), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(G15gat), .B(G43gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(G71gat), .B(G99gat), .ZN(new_n466));
  XOR2_X1   g265(.A(new_n465), .B(new_n466), .Z(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n342), .A2(new_n343), .A3(new_n316), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n343), .B1(new_n342), .B2(new_n316), .ZN(new_n470));
  NOR3_X1   g269(.A1(new_n469), .A2(new_n470), .A3(new_n347), .ZN(new_n471));
  INV_X1    g270(.A(new_n358), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n279), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n349), .A2(new_n277), .A3(new_n358), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(new_n462), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT33), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n468), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT68), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n477), .A2(new_n478), .B1(KEYINPUT32), .B2(new_n475), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n468), .A2(new_n476), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n475), .A2(KEYINPUT32), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n481), .B1(new_n477), .B2(KEYINPUT68), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n464), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n462), .ZN(new_n484));
  NOR3_X1   g283(.A1(new_n458), .A2(new_n459), .A3(new_n484), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n478), .B(new_n467), .C1(new_n485), .C2(KEYINPUT33), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n475), .A2(KEYINPUT32), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g287(.A(KEYINPUT68), .B(new_n467), .C1(new_n485), .C2(KEYINPUT33), .ZN(new_n489));
  INV_X1    g288(.A(new_n481), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n464), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n488), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(KEYINPUT69), .A2(KEYINPUT34), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n483), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n494), .B1(new_n483), .B2(new_n493), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n456), .A2(new_n457), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n448), .A2(new_n449), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n454), .A2(KEYINPUT86), .A3(new_n447), .A4(new_n439), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n440), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n494), .ZN(new_n502));
  NOR3_X1   g301(.A1(new_n479), .A2(new_n482), .A3(new_n464), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n492), .B1(new_n488), .B2(new_n491), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n483), .A2(new_n493), .A3(new_n494), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT88), .B1(new_n501), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n498), .A2(new_n508), .A3(KEYINPUT35), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT36), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n505), .A2(KEYINPUT36), .A3(new_n506), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(new_n501), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n402), .B1(new_n509), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n391), .A2(new_n388), .A3(new_n399), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n292), .A2(new_n293), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n285), .A2(new_n286), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT39), .ZN(new_n519));
  OR3_X1    g318(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  OR2_X1    g319(.A1(KEYINPUT87), .A2(KEYINPUT40), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n303), .B1(new_n518), .B2(new_n519), .ZN(new_n522));
  AND3_X1   g321(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n521), .B1(new_n520), .B2(new_n522), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n516), .A2(new_n525), .A3(new_n306), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT38), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n380), .A2(new_n527), .A3(new_n384), .A4(new_n396), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT37), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n395), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n380), .A2(KEYINPUT37), .A3(new_n384), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n396), .B1(new_n533), .B2(KEYINPUT38), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n362), .A2(new_n383), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n379), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n536), .B(KEYINPUT37), .C1(new_n379), .C2(new_n366), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n531), .A2(new_n537), .A3(new_n527), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n529), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n526), .B1(new_n539), .B2(new_n312), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n513), .A2(new_n540), .A3(new_n456), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT35), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n456), .A2(new_n497), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n542), .B1(new_n543), .B2(new_n400), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n249), .B1(new_n515), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT92), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(G230gat), .A2(G233gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(G99gat), .A2(G106gat), .ZN(new_n550));
  INV_X1    g349(.A(G85gat), .ZN(new_n551));
  INV_X1    g350(.A(G92gat), .ZN(new_n552));
  AOI22_X1  g351(.A1(KEYINPUT8), .A2(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT7), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n554), .B1(new_n551), .B2(new_n552), .ZN(new_n555));
  NAND3_X1  g354(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n553), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(G99gat), .B(G106gat), .Z(new_n558));
  AND2_X1   g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n557), .A2(new_n558), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT97), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n557), .B(new_n558), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT97), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  XOR2_X1   g364(.A(G57gat), .B(G64gat), .Z(new_n566));
  INV_X1    g365(.A(G71gat), .ZN(new_n567));
  INV_X1    g366(.A(G78gat), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n566), .B1(KEYINPUT9), .B2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G71gat), .B(G78gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n562), .A2(new_n565), .A3(KEYINPUT10), .A4(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT101), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n574), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n561), .A2(KEYINPUT100), .ZN(new_n578));
  INV_X1    g377(.A(new_n572), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT100), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n572), .A2(new_n563), .A3(new_n580), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT10), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n549), .B1(new_n577), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G120gat), .B(G148gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT103), .ZN(new_n587));
  XNOR2_X1  g386(.A(G176gat), .B(G204gat), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n587), .B(new_n588), .Z(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n582), .A2(new_n583), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n591), .A2(new_n549), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n590), .B1(new_n592), .B2(KEYINPUT102), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n585), .B(new_n593), .C1(KEYINPUT102), .C2(new_n592), .ZN(new_n594));
  INV_X1    g393(.A(new_n549), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n573), .B(KEYINPUT101), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT10), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n591), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n595), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n590), .B1(new_n599), .B2(new_n592), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  OAI211_X1 g401(.A(KEYINPUT92), .B(new_n249), .C1(new_n515), .C2(new_n545), .ZN(new_n603));
  AND3_X1   g402(.A1(new_n548), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT93), .ZN(new_n606));
  XOR2_X1   g405(.A(G127gat), .B(G155gat), .Z(new_n607));
  XOR2_X1   g406(.A(new_n606), .B(new_n607), .Z(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT21), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n235), .B1(new_n610), .B2(new_n579), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT94), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(G231gat), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n614), .A2(new_n314), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n613), .A2(new_n615), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n579), .A2(new_n610), .ZN(new_n619));
  XOR2_X1   g418(.A(G183gat), .B(G211gat), .Z(new_n620));
  XOR2_X1   g419(.A(new_n619), .B(new_n620), .Z(new_n621));
  NOR3_X1   g420(.A1(new_n617), .A2(new_n618), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n621), .ZN(new_n623));
  OR2_X1    g422(.A1(new_n613), .A2(new_n615), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n623), .B1(new_n624), .B2(new_n616), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n609), .B1(new_n622), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n621), .B1(new_n617), .B2(new_n618), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n624), .A2(new_n616), .A3(new_n623), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n627), .A2(new_n608), .A3(new_n628), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n562), .A2(new_n565), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(new_n222), .ZN(new_n632));
  NAND2_X1  g431(.A1(G232gat), .A2(G233gat), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n633), .B(KEYINPUT95), .Z(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(KEYINPUT41), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n632), .B(new_n636), .C1(new_n225), .C2(new_n631), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n635), .A2(KEYINPUT41), .ZN(new_n638));
  XNOR2_X1  g437(.A(KEYINPUT96), .B(KEYINPUT98), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n637), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G134gat), .B(G162gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(G190gat), .B(G218gat), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n642), .B(new_n643), .Z(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n641), .B(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n630), .A2(KEYINPUT99), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n626), .A2(new_n646), .A3(new_n629), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT99), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n604), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n312), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g454(.A(KEYINPUT16), .B(G8gat), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT104), .ZN(new_n657));
  AOI21_X1  g456(.A(KEYINPUT42), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n658), .B1(new_n657), .B2(new_n656), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n652), .A2(new_n516), .A3(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n660), .B1(new_n661), .B2(G8gat), .ZN(new_n662));
  INV_X1    g461(.A(new_n656), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n652), .A2(KEYINPUT42), .A3(new_n516), .A4(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n664), .A2(KEYINPUT105), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT105), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n604), .A2(new_n651), .ZN(new_n667));
  INV_X1    g466(.A(new_n516), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n667), .A2(new_n661), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n666), .B1(new_n669), .B2(new_n663), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n662), .B1(new_n665), .B2(new_n670), .ZN(G1325gat));
  AOI21_X1  g470(.A(G15gat), .B1(new_n652), .B2(new_n497), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n513), .A2(KEYINPUT106), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n513), .A2(KEYINPUT106), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n667), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n672), .B1(G15gat), .B2(new_n677), .ZN(G1326gat));
  NOR2_X1   g477(.A1(new_n667), .A2(new_n456), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT43), .B(G22gat), .Z(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1327gat));
  INV_X1    g480(.A(new_n630), .ZN(new_n682));
  INV_X1    g481(.A(new_n646), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n604), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n684), .A2(G29gat), .A3(new_n312), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(KEYINPUT45), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT45), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n601), .B(KEYINPUT107), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n683), .B1(new_n515), .B2(new_n545), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(KEYINPUT44), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n691), .B(new_n683), .C1(new_n515), .C2(new_n545), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n688), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n249), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n630), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n693), .A2(new_n653), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n687), .B1(new_n696), .B2(G29gat), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n686), .B1(new_n697), .B2(new_n685), .ZN(G1328gat));
  INV_X1    g497(.A(G36gat), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n516), .A2(new_n699), .ZN(new_n700));
  OR3_X1    g499(.A1(new_n684), .A2(KEYINPUT46), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT46), .B1(new_n684), .B2(new_n700), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n693), .A2(new_n516), .A3(new_n695), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n701), .B(new_n702), .C1(new_n699), .C2(new_n703), .ZN(G1329gat));
  INV_X1    g503(.A(new_n513), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n693), .A2(new_n705), .A3(new_n695), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(G43gat), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n507), .A2(G43gat), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n604), .A2(new_n682), .A3(new_n683), .A4(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n707), .A2(new_n709), .A3(KEYINPUT47), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n690), .A2(new_n692), .ZN(new_n712));
  INV_X1    g511(.A(new_n688), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n712), .A2(new_n675), .A3(new_n695), .A4(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(G43gat), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n711), .B1(new_n715), .B2(new_n709), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT109), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI211_X1 g517(.A(KEYINPUT109), .B(new_n711), .C1(new_n715), .C2(new_n709), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n710), .B1(new_n718), .B2(new_n719), .ZN(G1330gat));
  INV_X1    g519(.A(G50gat), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(new_n684), .B2(new_n456), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n693), .A2(G50gat), .A3(new_n501), .A4(new_n695), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT48), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT48), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n722), .A2(new_n723), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(G1331gat));
  NAND2_X1  g527(.A1(new_n509), .A2(new_n514), .ZN(new_n729));
  INV_X1    g528(.A(new_n402), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n545), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n249), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n651), .A2(new_n688), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n653), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g537(.A1(new_n735), .A2(new_n668), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  AND2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n739), .B2(new_n740), .ZN(G1333gat));
  NAND3_X1  g542(.A1(new_n736), .A2(new_n567), .A3(new_n497), .ZN(new_n744));
  OAI21_X1  g543(.A(G71gat), .B1(new_n735), .B2(new_n676), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g546(.A1(new_n735), .A2(new_n456), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(new_n568), .ZN(G1335gat));
  NOR2_X1   g548(.A1(new_n630), .A2(new_n249), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n751), .A2(new_n602), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n753), .B1(new_n690), .B2(new_n692), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(G85gat), .B1(new_n755), .B2(new_n312), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n731), .A2(new_n732), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n757), .A2(KEYINPUT51), .A3(new_n683), .A4(new_n750), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n683), .B(new_n750), .C1(new_n515), .C2(new_n545), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n602), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n762), .A2(new_n551), .A3(new_n653), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n756), .A2(new_n763), .ZN(G1336gat));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n691), .B1(new_n757), .B2(new_n683), .ZN(new_n766));
  INV_X1    g565(.A(new_n692), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n516), .B(new_n752), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G92gat), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n765), .B1(new_n769), .B2(KEYINPUT110), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n552), .B1(new_n754), .B2(new_n516), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n668), .A2(G92gat), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  AOI211_X1 g572(.A(new_n713), .B(new_n773), .C1(new_n758), .C2(new_n761), .ZN(new_n774));
  OAI21_X1  g573(.A(KEYINPUT111), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n776));
  INV_X1    g575(.A(new_n761), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n759), .A2(new_n760), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n688), .B(new_n772), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n769), .A2(new_n776), .A3(new_n779), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n770), .A2(new_n775), .A3(new_n780), .ZN(new_n781));
  AOI211_X1 g580(.A(new_n668), .B(new_n753), .C1(new_n690), .C2(new_n692), .ZN(new_n782));
  OAI21_X1  g581(.A(KEYINPUT110), .B1(new_n782), .B2(new_n552), .ZN(new_n783));
  AOI22_X1  g582(.A1(new_n775), .A2(new_n780), .B1(KEYINPUT52), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n781), .A2(new_n784), .ZN(G1337gat));
  OAI21_X1  g584(.A(G99gat), .B1(new_n755), .B2(new_n676), .ZN(new_n786));
  INV_X1    g585(.A(G99gat), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n762), .A2(new_n787), .A3(new_n497), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(G1338gat));
  NOR2_X1   g588(.A1(new_n755), .A2(new_n456), .ZN(new_n790));
  INV_X1    g589(.A(G106gat), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n688), .B1(new_n777), .B2(new_n778), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n501), .A2(new_n791), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(KEYINPUT53), .B1(new_n792), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797));
  OAI221_X1 g596(.A(new_n797), .B1(new_n793), .B2(new_n794), .C1(new_n790), .C2(new_n791), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(G1339gat));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n590), .B1(new_n585), .B2(KEYINPUT54), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n598), .A2(new_n575), .A3(new_n595), .A4(new_n576), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(KEYINPUT54), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n803), .A2(new_n599), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n800), .B1(new_n801), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n589), .B1(new_n599), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n585), .A2(KEYINPUT54), .A3(new_n802), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(new_n808), .A3(KEYINPUT55), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n805), .A2(new_n249), .A3(new_n594), .A4(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n236), .A2(new_n202), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n230), .A2(new_n223), .A3(new_n229), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n244), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT112), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OR2_X1    g614(.A1(new_n813), .A2(new_n814), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n601), .A2(new_n248), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n810), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT113), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT113), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n810), .A2(new_n820), .A3(new_n817), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n819), .A2(new_n646), .A3(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n805), .A2(new_n594), .A3(new_n809), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n816), .A2(new_n248), .A3(new_n815), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n823), .A2(new_n646), .A3(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n630), .B1(new_n822), .B2(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n647), .A2(new_n650), .A3(new_n602), .A4(new_n694), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(new_n312), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n668), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n498), .A2(new_n508), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OR3_X1    g634(.A1(new_n835), .A2(G113gat), .A3(new_n694), .ZN(new_n836));
  INV_X1    g635(.A(new_n543), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(G113gat), .B1(new_n838), .B2(new_n694), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n836), .A2(new_n839), .ZN(G1340gat));
  OR3_X1    g639(.A1(new_n835), .A2(G120gat), .A3(new_n602), .ZN(new_n841));
  OAI21_X1  g640(.A(G120gat), .B1(new_n838), .B2(new_n713), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(G1341gat));
  NOR3_X1   g642(.A1(new_n838), .A2(new_n273), .A3(new_n682), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n835), .A2(new_n682), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(KEYINPUT114), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n844), .B1(new_n846), .B2(new_n273), .ZN(G1342gat));
  OAI21_X1  g646(.A(G134gat), .B1(new_n838), .B2(new_n646), .ZN(new_n848));
  INV_X1    g647(.A(G134gat), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n516), .A2(new_n646), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(KEYINPUT115), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n831), .A2(new_n849), .A3(new_n834), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT56), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n852), .A2(KEYINPUT56), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n848), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT116), .ZN(G1343gat));
  OAI21_X1  g655(.A(new_n501), .B1(new_n827), .B2(new_n829), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n857), .A2(KEYINPUT57), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n683), .B1(new_n810), .B2(new_n817), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n825), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n861), .B1(new_n859), .B2(new_n860), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n829), .B1(new_n862), .B2(new_n682), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT57), .B1(new_n863), .B2(new_n456), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n705), .A2(new_n312), .A3(new_n516), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n858), .A2(new_n249), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n265), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n866), .A2(new_n867), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n676), .A2(new_n501), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n832), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n256), .A3(new_n249), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n871), .A2(new_n872), .A3(new_n875), .ZN(new_n876));
  AND3_X1   g675(.A1(new_n866), .A2(KEYINPUT118), .A3(new_n869), .ZN(new_n877));
  AOI21_X1  g676(.A(KEYINPUT118), .B1(new_n866), .B2(new_n869), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n879), .A2(new_n875), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n876), .B1(new_n880), .B2(new_n872), .ZN(G1344gat));
  NOR2_X1   g680(.A1(new_n260), .A2(new_n261), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n874), .A2(new_n883), .A3(new_n601), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n682), .B1(new_n860), .B2(new_n825), .ZN(new_n885));
  AOI211_X1 g684(.A(KEYINPUT57), .B(new_n456), .C1(new_n828), .C2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n886), .B1(new_n857), .B2(KEYINPUT57), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n601), .A3(new_n865), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n858), .A2(new_n864), .A3(new_n865), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n883), .B1(new_n891), .B2(new_n601), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n884), .B(new_n889), .C1(new_n892), .C2(KEYINPUT59), .ZN(G1345gat));
  AND3_X1   g692(.A1(new_n891), .A2(G155gat), .A3(new_n630), .ZN(new_n894));
  AOI21_X1  g693(.A(G155gat), .B1(new_n874), .B2(new_n630), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n894), .A2(new_n895), .ZN(G1346gat));
  NAND2_X1  g695(.A1(new_n831), .A2(new_n851), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n897), .A2(G162gat), .A3(new_n873), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT120), .ZN(new_n899));
  OAI21_X1  g698(.A(G162gat), .B1(new_n890), .B2(new_n646), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(G1347gat));
  NOR2_X1   g700(.A1(new_n830), .A2(new_n653), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n902), .A2(new_n516), .A3(new_n834), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n325), .A3(new_n249), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n902), .A2(new_n837), .A3(new_n516), .ZN(new_n905));
  OAI21_X1  g704(.A(G169gat), .B1(new_n905), .B2(new_n694), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(G1348gat));
  AOI21_X1  g706(.A(G176gat), .B1(new_n903), .B2(new_n601), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n905), .A2(new_n326), .A3(new_n713), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(G1349gat));
  OR3_X1    g709(.A1(new_n905), .A2(KEYINPUT121), .A3(new_n682), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT121), .B1(new_n905), .B2(new_n682), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(G183gat), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n903), .A2(new_n630), .A3(new_n354), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  OR2_X1    g715(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n916), .B(new_n917), .ZN(G1350gat));
  OAI21_X1  g717(.A(G190gat), .B1(new_n905), .B2(new_n646), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT61), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n903), .A2(new_n322), .A3(new_n683), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1351gat));
  NAND4_X1  g721(.A1(new_n673), .A2(new_n501), .A3(new_n516), .A4(new_n674), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n923), .A2(KEYINPUT123), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(KEYINPUT123), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n924), .A2(new_n902), .A3(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(G197gat), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n926), .A2(new_n927), .A3(new_n249), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n675), .A2(new_n668), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n887), .A2(new_n312), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(G197gat), .B1(new_n930), .B2(new_n694), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n928), .A2(new_n931), .ZN(G1352gat));
  INV_X1    g731(.A(G204gat), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n926), .A2(new_n933), .A3(new_n601), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n934), .A2(KEYINPUT62), .ZN(new_n935));
  OAI21_X1  g734(.A(G204gat), .B1(new_n930), .B2(new_n713), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(KEYINPUT62), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(G1353gat));
  NAND4_X1  g737(.A1(new_n887), .A2(new_n312), .A3(new_n630), .A4(new_n929), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(G211gat), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT63), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n939), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n942), .A2(KEYINPUT125), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n369), .A2(new_n371), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n926), .A2(KEYINPUT124), .A3(new_n630), .A4(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT124), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n924), .A2(new_n630), .A3(new_n902), .A4(new_n925), .ZN(new_n948));
  INV_X1    g747(.A(new_n945), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT125), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n940), .A2(new_n952), .A3(new_n941), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n944), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n944), .A2(KEYINPUT126), .A3(new_n951), .A4(new_n953), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(G1354gat));
  OAI21_X1  g757(.A(G218gat), .B1(new_n930), .B2(new_n646), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n926), .A2(new_n683), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n959), .B1(new_n960), .B2(G218gat), .ZN(new_n961));
  XOR2_X1   g760(.A(new_n961), .B(KEYINPUT127), .Z(G1355gat));
endmodule


