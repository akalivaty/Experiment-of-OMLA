

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U556 ( .A(n567), .Z(n521) );
  BUF_X1 U557 ( .A(n602), .Z(n524) );
  XNOR2_X1 U558 ( .A(n804), .B(n803), .ZN(n811) );
  AND2_X1 U559 ( .A1(n802), .A2(n801), .ZN(n804) );
  AND2_X1 U560 ( .A1(n759), .A2(n758), .ZN(n760) );
  INV_X1 U561 ( .A(n761), .ZN(n780) );
  AND2_X2 U562 ( .A1(n530), .A2(G2104), .ZN(n899) );
  XNOR2_X1 U563 ( .A(n523), .B(n522), .ZN(n832) );
  INV_X1 U564 ( .A(KEYINPUT110), .ZN(n522) );
  NAND2_X1 U565 ( .A1(n831), .A2(n830), .ZN(n523) );
  XNOR2_X1 U566 ( .A(n526), .B(n525), .ZN(n567) );
  XNOR2_X1 U567 ( .A(KEYINPUT1), .B(n537), .ZN(n602) );
  NOR2_X1 U568 ( .A1(n739), .A2(n738), .ZN(n741) );
  NOR2_X1 U569 ( .A1(G543), .A2(n542), .ZN(n536) );
  NOR2_X1 U570 ( .A1(n535), .A2(n534), .ZN(G160) );
  NOR2_X2 U571 ( .A1(G651), .A2(n645), .ZN(n656) );
  AND2_X1 U572 ( .A1(n1021), .A2(G1348), .ZN(n745) );
  INV_X1 U573 ( .A(G8), .ZN(n734) );
  OR2_X1 U574 ( .A1(n794), .A2(n734), .ZN(n735) );
  XNOR2_X1 U575 ( .A(n773), .B(KEYINPUT29), .ZN(n774) );
  INV_X1 U576 ( .A(KEYINPUT31), .ZN(n740) );
  NOR2_X1 U577 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U578 ( .A(n733), .B(KEYINPUT95), .ZN(n817) );
  INV_X1 U579 ( .A(KEYINPUT108), .ZN(n803) );
  NAND2_X1 U580 ( .A1(G160), .A2(G40), .ZN(n725) );
  NOR2_X1 U581 ( .A1(n833), .A2(n832), .ZN(n835) );
  AND2_X1 U582 ( .A1(n608), .A2(n607), .ZN(n610) );
  NOR2_X2 U583 ( .A1(n645), .A2(n542), .ZN(n659) );
  XOR2_X1 U584 ( .A(KEYINPUT70), .B(n548), .Z(G299) );
  XNOR2_X1 U585 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n526) );
  NOR2_X1 U586 ( .A1(G2105), .A2(G2104), .ZN(n525) );
  NAND2_X1 U587 ( .A1(n521), .A2(G137), .ZN(n529) );
  INV_X1 U588 ( .A(G2105), .ZN(n530) );
  NAND2_X1 U589 ( .A1(G101), .A2(n899), .ZN(n527) );
  XOR2_X1 U590 ( .A(KEYINPUT23), .B(n527), .Z(n528) );
  NAND2_X1 U591 ( .A1(n529), .A2(n528), .ZN(n535) );
  NOR2_X1 U592 ( .A1(G2104), .A2(n530), .ZN(n563) );
  BUF_X1 U593 ( .A(n563), .Z(n895) );
  NAND2_X1 U594 ( .A1(G125), .A2(n895), .ZN(n533) );
  NAND2_X1 U595 ( .A1(G2104), .A2(G2105), .ZN(n531) );
  XOR2_X1 U596 ( .A(KEYINPUT64), .B(n531), .Z(n627) );
  NAND2_X1 U597 ( .A1(G113), .A2(n627), .ZN(n532) );
  NAND2_X1 U598 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U599 ( .A(KEYINPUT0), .B(G543), .Z(n645) );
  NAND2_X1 U600 ( .A1(n656), .A2(G53), .ZN(n539) );
  XOR2_X1 U601 ( .A(n536), .B(KEYINPUT66), .Z(n537) );
  NAND2_X1 U602 ( .A1(G65), .A2(n524), .ZN(n538) );
  NAND2_X1 U603 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U604 ( .A(n540), .B(KEYINPUT69), .Z(n541) );
  INV_X1 U605 ( .A(n541), .ZN(n544) );
  INV_X1 U606 ( .A(G651), .ZN(n542) );
  NAND2_X1 U607 ( .A1(G78), .A2(n659), .ZN(n543) );
  NAND2_X1 U608 ( .A1(n544), .A2(n543), .ZN(n547) );
  NOR2_X1 U609 ( .A1(G651), .A2(G543), .ZN(n663) );
  NAND2_X1 U610 ( .A1(n663), .A2(G91), .ZN(n545) );
  XOR2_X1 U611 ( .A(KEYINPUT68), .B(n545), .Z(n546) );
  NOR2_X1 U612 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U613 ( .A1(G76), .A2(n659), .ZN(n552) );
  XOR2_X1 U614 ( .A(KEYINPUT4), .B(KEYINPUT75), .Z(n550) );
  NAND2_X1 U615 ( .A1(G89), .A2(n663), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(n551) );
  NAND2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n553), .B(KEYINPUT76), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n554), .B(KEYINPUT5), .ZN(n561) );
  XNOR2_X1 U620 ( .A(KEYINPUT6), .B(KEYINPUT78), .ZN(n559) );
  NAND2_X1 U621 ( .A1(n656), .A2(G51), .ZN(n557) );
  NAND2_X1 U622 ( .A1(G63), .A2(n524), .ZN(n555) );
  XOR2_X1 U623 ( .A(KEYINPUT77), .B(n555), .Z(n556) );
  NAND2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U625 ( .A(n559), .B(n558), .Z(n560) );
  NAND2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n562), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U628 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U629 ( .A1(G114), .A2(n627), .ZN(n565) );
  NAND2_X1 U630 ( .A1(G126), .A2(n563), .ZN(n564) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U632 ( .A(KEYINPUT90), .B(n566), .Z(n573) );
  NAND2_X1 U633 ( .A1(n567), .A2(G138), .ZN(n571) );
  NAND2_X1 U634 ( .A1(G102), .A2(n899), .ZN(n568) );
  XNOR2_X1 U635 ( .A(KEYINPUT91), .B(n568), .ZN(n569) );
  INV_X1 U636 ( .A(n569), .ZN(n570) );
  AND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  AND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(G164) );
  NAND2_X1 U639 ( .A1(G85), .A2(n663), .ZN(n575) );
  NAND2_X1 U640 ( .A1(G60), .A2(n524), .ZN(n574) );
  NAND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n579) );
  NAND2_X1 U642 ( .A1(G72), .A2(n659), .ZN(n577) );
  NAND2_X1 U643 ( .A1(G47), .A2(n656), .ZN(n576) );
  NAND2_X1 U644 ( .A1(n577), .A2(n576), .ZN(n578) );
  OR2_X1 U645 ( .A1(n579), .A2(n578), .ZN(G290) );
  AND2_X1 U646 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U647 ( .A(G132), .ZN(G219) );
  INV_X1 U648 ( .A(G82), .ZN(G220) );
  INV_X1 U649 ( .A(G120), .ZN(G236) );
  INV_X1 U650 ( .A(G69), .ZN(G235) );
  INV_X1 U651 ( .A(G108), .ZN(G238) );
  NAND2_X1 U652 ( .A1(n524), .A2(G64), .ZN(n580) );
  XNOR2_X1 U653 ( .A(n580), .B(KEYINPUT67), .ZN(n587) );
  NAND2_X1 U654 ( .A1(G90), .A2(n663), .ZN(n582) );
  NAND2_X1 U655 ( .A1(G77), .A2(n659), .ZN(n581) );
  NAND2_X1 U656 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U657 ( .A(n583), .B(KEYINPUT9), .ZN(n585) );
  NAND2_X1 U658 ( .A1(G52), .A2(n656), .ZN(n584) );
  NAND2_X1 U659 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U660 ( .A1(n587), .A2(n586), .ZN(G171) );
  XOR2_X1 U661 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n589) );
  NAND2_X1 U662 ( .A1(G7), .A2(G661), .ZN(n588) );
  XNOR2_X1 U663 ( .A(n589), .B(n588), .ZN(G223) );
  INV_X1 U664 ( .A(G223), .ZN(n853) );
  NAND2_X1 U665 ( .A1(n853), .A2(G567), .ZN(n590) );
  XOR2_X1 U666 ( .A(KEYINPUT11), .B(n590), .Z(G234) );
  NAND2_X1 U667 ( .A1(n663), .A2(G81), .ZN(n591) );
  XNOR2_X1 U668 ( .A(n591), .B(KEYINPUT12), .ZN(n593) );
  NAND2_X1 U669 ( .A1(G68), .A2(n659), .ZN(n592) );
  NAND2_X1 U670 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U671 ( .A(KEYINPUT13), .B(n594), .ZN(n601) );
  XOR2_X1 U672 ( .A(KEYINPUT72), .B(KEYINPUT14), .Z(n596) );
  NAND2_X1 U673 ( .A1(G56), .A2(n524), .ZN(n595) );
  XNOR2_X1 U674 ( .A(n596), .B(n595), .ZN(n599) );
  NAND2_X1 U675 ( .A1(G43), .A2(n656), .ZN(n597) );
  XNOR2_X1 U676 ( .A(KEYINPUT73), .B(n597), .ZN(n598) );
  NOR2_X1 U677 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U678 ( .A1(n601), .A2(n600), .ZN(n1014) );
  INV_X1 U679 ( .A(G860), .ZN(n636) );
  OR2_X1 U680 ( .A1(n1014), .A2(n636), .ZN(G153) );
  INV_X1 U681 ( .A(G171), .ZN(G301) );
  NAND2_X1 U682 ( .A1(G66), .A2(n602), .ZN(n608) );
  AND2_X1 U683 ( .A1(n656), .A2(G54), .ZN(n606) );
  NAND2_X1 U684 ( .A1(G79), .A2(n659), .ZN(n604) );
  NAND2_X1 U685 ( .A1(G92), .A2(n663), .ZN(n603) );
  NAND2_X1 U686 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U687 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U688 ( .A(KEYINPUT74), .B(KEYINPUT15), .ZN(n609) );
  XNOR2_X2 U689 ( .A(n610), .B(n609), .ZN(n1021) );
  NOR2_X1 U690 ( .A1(n1021), .A2(G868), .ZN(n612) );
  INV_X1 U691 ( .A(G868), .ZN(n676) );
  NOR2_X1 U692 ( .A1(n676), .A2(G301), .ZN(n611) );
  NOR2_X1 U693 ( .A1(n612), .A2(n611), .ZN(G284) );
  XNOR2_X1 U694 ( .A(KEYINPUT79), .B(G868), .ZN(n613) );
  NOR2_X1 U695 ( .A1(G286), .A2(n613), .ZN(n615) );
  NOR2_X1 U696 ( .A1(G299), .A2(G868), .ZN(n614) );
  NOR2_X1 U697 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U698 ( .A(KEYINPUT80), .B(n616), .ZN(G297) );
  NAND2_X1 U699 ( .A1(n636), .A2(G559), .ZN(n617) );
  INV_X1 U700 ( .A(n1021), .ZN(n634) );
  NAND2_X1 U701 ( .A1(n617), .A2(n634), .ZN(n618) );
  XNOR2_X1 U702 ( .A(n618), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U703 ( .A1(n1021), .A2(n676), .ZN(n619) );
  XNOR2_X1 U704 ( .A(n619), .B(KEYINPUT81), .ZN(n620) );
  NOR2_X1 U705 ( .A1(G559), .A2(n620), .ZN(n621) );
  XNOR2_X1 U706 ( .A(n621), .B(KEYINPUT82), .ZN(n623) );
  NOR2_X1 U707 ( .A1(n1014), .A2(G868), .ZN(n622) );
  NOR2_X1 U708 ( .A1(n623), .A2(n622), .ZN(G282) );
  NAND2_X1 U709 ( .A1(n895), .A2(G123), .ZN(n624) );
  XNOR2_X1 U710 ( .A(n624), .B(KEYINPUT18), .ZN(n626) );
  NAND2_X1 U711 ( .A1(G99), .A2(n899), .ZN(n625) );
  NAND2_X1 U712 ( .A1(n626), .A2(n625), .ZN(n631) );
  NAND2_X1 U713 ( .A1(n521), .A2(G135), .ZN(n629) );
  BUF_X1 U714 ( .A(n627), .Z(n896) );
  NAND2_X1 U715 ( .A1(G111), .A2(n896), .ZN(n628) );
  NAND2_X1 U716 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U717 ( .A1(n631), .A2(n630), .ZN(n949) );
  XNOR2_X1 U718 ( .A(n949), .B(G2096), .ZN(n633) );
  INV_X1 U719 ( .A(G2100), .ZN(n632) );
  NAND2_X1 U720 ( .A1(n633), .A2(n632), .ZN(G156) );
  NAND2_X1 U721 ( .A1(n634), .A2(G559), .ZN(n635) );
  XOR2_X1 U722 ( .A(n1014), .B(n635), .Z(n674) );
  NAND2_X1 U723 ( .A1(n636), .A2(n674), .ZN(n644) );
  NAND2_X1 U724 ( .A1(G93), .A2(n663), .ZN(n638) );
  NAND2_X1 U725 ( .A1(G67), .A2(n524), .ZN(n637) );
  NAND2_X1 U726 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U727 ( .A1(G80), .A2(n659), .ZN(n639) );
  XNOR2_X1 U728 ( .A(KEYINPUT83), .B(n639), .ZN(n640) );
  NOR2_X1 U729 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U730 ( .A1(n656), .A2(G55), .ZN(n642) );
  NAND2_X1 U731 ( .A1(n643), .A2(n642), .ZN(n677) );
  XNOR2_X1 U732 ( .A(n644), .B(n677), .ZN(G145) );
  NAND2_X1 U733 ( .A1(G87), .A2(n645), .ZN(n647) );
  NAND2_X1 U734 ( .A1(G74), .A2(G651), .ZN(n646) );
  NAND2_X1 U735 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U736 ( .A1(n524), .A2(n648), .ZN(n650) );
  NAND2_X1 U737 ( .A1(n656), .A2(G49), .ZN(n649) );
  NAND2_X1 U738 ( .A1(n650), .A2(n649), .ZN(G288) );
  NAND2_X1 U739 ( .A1(G88), .A2(n663), .ZN(n652) );
  NAND2_X1 U740 ( .A1(G62), .A2(n524), .ZN(n651) );
  NAND2_X1 U741 ( .A1(n652), .A2(n651), .ZN(n655) );
  NAND2_X1 U742 ( .A1(G75), .A2(n659), .ZN(n653) );
  XNOR2_X1 U743 ( .A(KEYINPUT85), .B(n653), .ZN(n654) );
  NOR2_X1 U744 ( .A1(n655), .A2(n654), .ZN(n658) );
  NAND2_X1 U745 ( .A1(n656), .A2(G50), .ZN(n657) );
  NAND2_X1 U746 ( .A1(n658), .A2(n657), .ZN(G303) );
  INV_X1 U747 ( .A(G303), .ZN(G166) );
  NAND2_X1 U748 ( .A1(G73), .A2(n659), .ZN(n660) );
  XNOR2_X1 U749 ( .A(n660), .B(KEYINPUT2), .ZN(n668) );
  NAND2_X1 U750 ( .A1(n656), .A2(G48), .ZN(n662) );
  NAND2_X1 U751 ( .A1(G61), .A2(n524), .ZN(n661) );
  NAND2_X1 U752 ( .A1(n662), .A2(n661), .ZN(n666) );
  NAND2_X1 U753 ( .A1(n663), .A2(G86), .ZN(n664) );
  XOR2_X1 U754 ( .A(KEYINPUT84), .B(n664), .Z(n665) );
  NOR2_X1 U755 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U756 ( .A1(n668), .A2(n667), .ZN(G305) );
  XNOR2_X1 U757 ( .A(KEYINPUT19), .B(G288), .ZN(n673) );
  XNOR2_X1 U758 ( .A(G299), .B(G305), .ZN(n669) );
  XNOR2_X1 U759 ( .A(n669), .B(n677), .ZN(n670) );
  XNOR2_X1 U760 ( .A(G166), .B(n670), .ZN(n671) );
  XNOR2_X1 U761 ( .A(n671), .B(G290), .ZN(n672) );
  XNOR2_X1 U762 ( .A(n673), .B(n672), .ZN(n920) );
  XOR2_X1 U763 ( .A(n920), .B(n674), .Z(n675) );
  NOR2_X1 U764 ( .A1(n676), .A2(n675), .ZN(n679) );
  NOR2_X1 U765 ( .A1(G868), .A2(n677), .ZN(n678) );
  NOR2_X1 U766 ( .A1(n679), .A2(n678), .ZN(G295) );
  NAND2_X1 U767 ( .A1(G2084), .A2(G2078), .ZN(n681) );
  XOR2_X1 U768 ( .A(KEYINPUT20), .B(KEYINPUT86), .Z(n680) );
  XNOR2_X1 U769 ( .A(n681), .B(n680), .ZN(n682) );
  NAND2_X1 U770 ( .A1(n682), .A2(G2090), .ZN(n683) );
  XOR2_X1 U771 ( .A(KEYINPUT87), .B(n683), .Z(n684) );
  XNOR2_X1 U772 ( .A(KEYINPUT21), .B(n684), .ZN(n685) );
  NAND2_X1 U773 ( .A1(n685), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U774 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U775 ( .A1(G235), .A2(G236), .ZN(n686) );
  XNOR2_X1 U776 ( .A(n686), .B(KEYINPUT89), .ZN(n687) );
  NOR2_X1 U777 ( .A1(G238), .A2(n687), .ZN(n688) );
  NAND2_X1 U778 ( .A1(G57), .A2(n688), .ZN(n857) );
  NAND2_X1 U779 ( .A1(n857), .A2(G567), .ZN(n694) );
  NOR2_X1 U780 ( .A1(G220), .A2(G219), .ZN(n689) );
  XNOR2_X1 U781 ( .A(KEYINPUT22), .B(n689), .ZN(n690) );
  NAND2_X1 U782 ( .A1(n690), .A2(G96), .ZN(n691) );
  NOR2_X1 U783 ( .A1(G218), .A2(n691), .ZN(n692) );
  XOR2_X1 U784 ( .A(KEYINPUT88), .B(n692), .Z(n858) );
  NAND2_X1 U785 ( .A1(n858), .A2(G2106), .ZN(n693) );
  NAND2_X1 U786 ( .A1(n694), .A2(n693), .ZN(n859) );
  NAND2_X1 U787 ( .A1(G483), .A2(G661), .ZN(n695) );
  NOR2_X1 U788 ( .A1(n859), .A2(n695), .ZN(n856) );
  NAND2_X1 U789 ( .A1(n856), .A2(G36), .ZN(G176) );
  NAND2_X1 U790 ( .A1(G105), .A2(n899), .ZN(n696) );
  XOR2_X1 U791 ( .A(KEYINPUT38), .B(n696), .Z(n701) );
  NAND2_X1 U792 ( .A1(G129), .A2(n895), .ZN(n698) );
  NAND2_X1 U793 ( .A1(G117), .A2(n896), .ZN(n697) );
  NAND2_X1 U794 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U795 ( .A(KEYINPUT93), .B(n699), .Z(n700) );
  NOR2_X1 U796 ( .A1(n701), .A2(n700), .ZN(n703) );
  NAND2_X1 U797 ( .A1(n521), .A2(G141), .ZN(n702) );
  NAND2_X1 U798 ( .A1(n703), .A2(n702), .ZN(n914) );
  NAND2_X1 U799 ( .A1(G1996), .A2(n914), .ZN(n704) );
  XOR2_X1 U800 ( .A(KEYINPUT94), .B(n704), .Z(n712) );
  NAND2_X1 U801 ( .A1(G119), .A2(n895), .ZN(n706) );
  NAND2_X1 U802 ( .A1(G131), .A2(n521), .ZN(n705) );
  NAND2_X1 U803 ( .A1(n706), .A2(n705), .ZN(n710) );
  NAND2_X1 U804 ( .A1(n899), .A2(G95), .ZN(n708) );
  NAND2_X1 U805 ( .A1(G107), .A2(n896), .ZN(n707) );
  NAND2_X1 U806 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U807 ( .A1(n710), .A2(n709), .ZN(n910) );
  INV_X1 U808 ( .A(G1991), .ZN(n836) );
  NOR2_X1 U809 ( .A1(n910), .A2(n836), .ZN(n711) );
  NOR2_X1 U810 ( .A1(n712), .A2(n711), .ZN(n960) );
  NOR2_X1 U811 ( .A1(G164), .A2(G1384), .ZN(n727) );
  NOR2_X1 U812 ( .A1(n727), .A2(n725), .ZN(n847) );
  INV_X1 U813 ( .A(n847), .ZN(n713) );
  NOR2_X1 U814 ( .A1(n960), .A2(n713), .ZN(n839) );
  INV_X1 U815 ( .A(n839), .ZN(n724) );
  NAND2_X1 U816 ( .A1(G104), .A2(n899), .ZN(n715) );
  NAND2_X1 U817 ( .A1(G140), .A2(n521), .ZN(n714) );
  NAND2_X1 U818 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U819 ( .A(KEYINPUT34), .B(n716), .ZN(n722) );
  NAND2_X1 U820 ( .A1(n895), .A2(G128), .ZN(n717) );
  XNOR2_X1 U821 ( .A(n717), .B(KEYINPUT92), .ZN(n719) );
  NAND2_X1 U822 ( .A1(G116), .A2(n896), .ZN(n718) );
  NAND2_X1 U823 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U824 ( .A(KEYINPUT35), .B(n720), .Z(n721) );
  NOR2_X1 U825 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U826 ( .A(KEYINPUT36), .B(n723), .ZN(n894) );
  XNOR2_X1 U827 ( .A(G2067), .B(KEYINPUT37), .ZN(n845) );
  NOR2_X1 U828 ( .A1(n894), .A2(n845), .ZN(n947) );
  NAND2_X1 U829 ( .A1(n847), .A2(n947), .ZN(n843) );
  NAND2_X1 U830 ( .A1(n724), .A2(n843), .ZN(n833) );
  INV_X1 U831 ( .A(n725), .ZN(n726) );
  AND2_X4 U832 ( .A1(n727), .A2(n726), .ZN(n761) );
  XNOR2_X1 U833 ( .A(G2078), .B(KEYINPUT25), .ZN(n728) );
  XNOR2_X1 U834 ( .A(n728), .B(KEYINPUT96), .ZN(n967) );
  NAND2_X1 U835 ( .A1(n761), .A2(n967), .ZN(n729) );
  XNOR2_X1 U836 ( .A(n729), .B(KEYINPUT97), .ZN(n731) );
  NOR2_X1 U837 ( .A1(n761), .A2(G1961), .ZN(n730) );
  NOR2_X1 U838 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U839 ( .A(KEYINPUT98), .B(n732), .Z(n742) );
  NOR2_X1 U840 ( .A1(G171), .A2(n742), .ZN(n739) );
  NAND2_X1 U841 ( .A1(n780), .A2(G8), .ZN(n733) );
  INV_X1 U842 ( .A(n817), .ZN(n819) );
  NOR2_X1 U843 ( .A1(G1966), .A2(n819), .ZN(n791) );
  NOR2_X1 U844 ( .A1(G2084), .A2(n780), .ZN(n794) );
  OR2_X1 U845 ( .A1(n791), .A2(n735), .ZN(n736) );
  XNOR2_X1 U846 ( .A(n736), .B(KEYINPUT30), .ZN(n737) );
  NOR2_X1 U847 ( .A1(G168), .A2(n737), .ZN(n738) );
  XNOR2_X1 U848 ( .A(n741), .B(n740), .ZN(n789) );
  NAND2_X1 U849 ( .A1(G171), .A2(n742), .ZN(n777) );
  INV_X1 U850 ( .A(G1341), .ZN(n743) );
  NAND2_X1 U851 ( .A1(KEYINPUT26), .A2(n743), .ZN(n744) );
  NOR2_X1 U852 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U853 ( .A1(n746), .A2(n761), .ZN(n747) );
  NOR2_X1 U854 ( .A1(n747), .A2(n1014), .ZN(n754) );
  OR2_X1 U855 ( .A1(G1996), .A2(KEYINPUT26), .ZN(n752) );
  NAND2_X1 U856 ( .A1(n1021), .A2(G2067), .ZN(n749) );
  NAND2_X1 U857 ( .A1(KEYINPUT26), .A2(G1996), .ZN(n748) );
  NAND2_X1 U858 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U859 ( .A1(n750), .A2(n761), .ZN(n751) );
  AND2_X1 U860 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U861 ( .A1(n754), .A2(n753), .ZN(n759) );
  NAND2_X1 U862 ( .A1(G1348), .A2(n780), .ZN(n756) );
  NAND2_X1 U863 ( .A1(G2067), .A2(n761), .ZN(n755) );
  NAND2_X1 U864 ( .A1(n756), .A2(n755), .ZN(n757) );
  OR2_X1 U865 ( .A1(n1021), .A2(n757), .ZN(n758) );
  XOR2_X1 U866 ( .A(n760), .B(KEYINPUT100), .Z(n767) );
  NAND2_X1 U867 ( .A1(G1956), .A2(n780), .ZN(n764) );
  NAND2_X1 U868 ( .A1(n761), .A2(G2072), .ZN(n762) );
  XOR2_X1 U869 ( .A(KEYINPUT27), .B(n762), .Z(n763) );
  NAND2_X1 U870 ( .A1(n764), .A2(n763), .ZN(n765) );
  XOR2_X1 U871 ( .A(KEYINPUT99), .B(n765), .Z(n769) );
  NOR2_X1 U872 ( .A1(G299), .A2(n769), .ZN(n766) );
  NOR2_X1 U873 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U874 ( .A(KEYINPUT101), .B(n768), .ZN(n772) );
  NAND2_X1 U875 ( .A1(G299), .A2(n769), .ZN(n770) );
  XNOR2_X1 U876 ( .A(KEYINPUT28), .B(n770), .ZN(n771) );
  NAND2_X1 U877 ( .A1(n772), .A2(n771), .ZN(n775) );
  XNOR2_X1 U878 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n773) );
  XNOR2_X1 U879 ( .A(n775), .B(n774), .ZN(n776) );
  NAND2_X1 U880 ( .A1(n777), .A2(n776), .ZN(n790) );
  NAND2_X1 U881 ( .A1(n789), .A2(n790), .ZN(n778) );
  NAND2_X1 U882 ( .A1(n778), .A2(G286), .ZN(n785) );
  NOR2_X1 U883 ( .A1(G1971), .A2(n819), .ZN(n779) );
  XOR2_X1 U884 ( .A(KEYINPUT105), .B(n779), .Z(n782) );
  NOR2_X1 U885 ( .A1(G2090), .A2(n780), .ZN(n781) );
  NOR2_X1 U886 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U887 ( .A1(n783), .A2(G303), .ZN(n784) );
  NAND2_X1 U888 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U889 ( .A(n786), .B(KEYINPUT106), .ZN(n787) );
  NAND2_X1 U890 ( .A1(n787), .A2(G8), .ZN(n788) );
  XNOR2_X1 U891 ( .A(n788), .B(KEYINPUT32), .ZN(n821) );
  AND2_X1 U892 ( .A1(n790), .A2(n789), .ZN(n792) );
  XNOR2_X1 U893 ( .A(n793), .B(KEYINPUT104), .ZN(n796) );
  NAND2_X1 U894 ( .A1(n794), .A2(G8), .ZN(n795) );
  NAND2_X1 U895 ( .A1(n796), .A2(n795), .ZN(n820) );
  NAND2_X1 U896 ( .A1(G1976), .A2(G288), .ZN(n1018) );
  AND2_X1 U897 ( .A1(n820), .A2(n1018), .ZN(n797) );
  NAND2_X1 U898 ( .A1(n821), .A2(n797), .ZN(n802) );
  INV_X1 U899 ( .A(n1018), .ZN(n800) );
  NOR2_X1 U900 ( .A1(G1976), .A2(G288), .ZN(n805) );
  NOR2_X1 U901 ( .A1(G1971), .A2(G303), .ZN(n798) );
  OR2_X1 U902 ( .A1(n805), .A2(n798), .ZN(n1020) );
  XNOR2_X1 U903 ( .A(n1020), .B(KEYINPUT107), .ZN(n799) );
  OR2_X1 U904 ( .A1(n800), .A2(n799), .ZN(n801) );
  INV_X1 U905 ( .A(KEYINPUT33), .ZN(n813) );
  NAND2_X1 U906 ( .A1(n817), .A2(n805), .ZN(n806) );
  NOR2_X1 U907 ( .A1(n813), .A2(n806), .ZN(n807) );
  XNOR2_X1 U908 ( .A(n807), .B(KEYINPUT109), .ZN(n812) );
  AND2_X1 U909 ( .A1(n817), .A2(n812), .ZN(n809) );
  XNOR2_X1 U910 ( .A(G1981), .B(G305), .ZN(n1028) );
  INV_X1 U911 ( .A(n1028), .ZN(n808) );
  AND2_X1 U912 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U913 ( .A1(n811), .A2(n810), .ZN(n831) );
  INV_X1 U914 ( .A(n812), .ZN(n814) );
  OR2_X1 U915 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U916 ( .A1(n1028), .A2(n815), .ZN(n829) );
  NOR2_X1 U917 ( .A1(G1981), .A2(G305), .ZN(n816) );
  XNOR2_X1 U918 ( .A(KEYINPUT24), .B(n816), .ZN(n818) );
  NAND2_X1 U919 ( .A1(n818), .A2(n817), .ZN(n827) );
  NAND2_X1 U920 ( .A1(n821), .A2(n820), .ZN(n824) );
  NOR2_X1 U921 ( .A1(G2090), .A2(G303), .ZN(n822) );
  NAND2_X1 U922 ( .A1(G8), .A2(n822), .ZN(n823) );
  NAND2_X1 U923 ( .A1(n824), .A2(n823), .ZN(n825) );
  NAND2_X1 U924 ( .A1(n819), .A2(n825), .ZN(n826) );
  NAND2_X1 U925 ( .A1(n827), .A2(n826), .ZN(n828) );
  NOR2_X1 U926 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U927 ( .A(G1986), .B(G290), .ZN(n1019) );
  NAND2_X1 U928 ( .A1(n1019), .A2(n847), .ZN(n834) );
  NAND2_X1 U929 ( .A1(n835), .A2(n834), .ZN(n850) );
  XOR2_X1 U930 ( .A(KEYINPUT39), .B(KEYINPUT111), .Z(n842) );
  NOR2_X1 U931 ( .A1(G1996), .A2(n914), .ZN(n944) );
  AND2_X1 U932 ( .A1(n836), .A2(n910), .ZN(n953) );
  NOR2_X1 U933 ( .A1(G1986), .A2(G290), .ZN(n837) );
  NOR2_X1 U934 ( .A1(n953), .A2(n837), .ZN(n838) );
  NOR2_X1 U935 ( .A1(n839), .A2(n838), .ZN(n840) );
  NOR2_X1 U936 ( .A1(n944), .A2(n840), .ZN(n841) );
  XNOR2_X1 U937 ( .A(n842), .B(n841), .ZN(n844) );
  NAND2_X1 U938 ( .A1(n844), .A2(n843), .ZN(n846) );
  NAND2_X1 U939 ( .A1(n894), .A2(n845), .ZN(n950) );
  NAND2_X1 U940 ( .A1(n846), .A2(n950), .ZN(n848) );
  NAND2_X1 U941 ( .A1(n848), .A2(n847), .ZN(n849) );
  NAND2_X1 U942 ( .A1(n850), .A2(n849), .ZN(n852) );
  XNOR2_X1 U943 ( .A(KEYINPUT40), .B(KEYINPUT112), .ZN(n851) );
  XNOR2_X1 U944 ( .A(n852), .B(n851), .ZN(G329) );
  NAND2_X1 U945 ( .A1(G2106), .A2(n853), .ZN(G217) );
  AND2_X1 U946 ( .A1(G15), .A2(G2), .ZN(n854) );
  NAND2_X1 U947 ( .A1(G661), .A2(n854), .ZN(G259) );
  NAND2_X1 U948 ( .A1(G3), .A2(G1), .ZN(n855) );
  NAND2_X1 U949 ( .A1(n856), .A2(n855), .ZN(G188) );
  XNOR2_X1 U950 ( .A(G96), .B(KEYINPUT115), .ZN(G221) );
  NOR2_X1 U952 ( .A1(n858), .A2(n857), .ZN(G325) );
  INV_X1 U953 ( .A(G325), .ZN(G261) );
  INV_X1 U954 ( .A(n859), .ZN(G319) );
  XOR2_X1 U955 ( .A(G2100), .B(G2096), .Z(n861) );
  XNOR2_X1 U956 ( .A(KEYINPUT42), .B(G2678), .ZN(n860) );
  XNOR2_X1 U957 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U958 ( .A(KEYINPUT43), .B(G2090), .Z(n863) );
  XNOR2_X1 U959 ( .A(G2067), .B(G2072), .ZN(n862) );
  XNOR2_X1 U960 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U961 ( .A(n865), .B(n864), .Z(n867) );
  XNOR2_X1 U962 ( .A(G2084), .B(G2078), .ZN(n866) );
  XNOR2_X1 U963 ( .A(n867), .B(n866), .ZN(G227) );
  XOR2_X1 U964 ( .A(KEYINPUT117), .B(G1976), .Z(n869) );
  XNOR2_X1 U965 ( .A(G1966), .B(G1961), .ZN(n868) );
  XNOR2_X1 U966 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U967 ( .A(n870), .B(KEYINPUT41), .Z(n872) );
  XNOR2_X1 U968 ( .A(G1996), .B(G1991), .ZN(n871) );
  XNOR2_X1 U969 ( .A(n872), .B(n871), .ZN(n876) );
  XOR2_X1 U970 ( .A(G1981), .B(G1971), .Z(n874) );
  XNOR2_X1 U971 ( .A(G1986), .B(G1956), .ZN(n873) );
  XNOR2_X1 U972 ( .A(n874), .B(n873), .ZN(n875) );
  XOR2_X1 U973 ( .A(n876), .B(n875), .Z(n878) );
  XNOR2_X1 U974 ( .A(KEYINPUT116), .B(G2474), .ZN(n877) );
  XNOR2_X1 U975 ( .A(n878), .B(n877), .ZN(G229) );
  NAND2_X1 U976 ( .A1(n895), .A2(G124), .ZN(n879) );
  XNOR2_X1 U977 ( .A(n879), .B(KEYINPUT44), .ZN(n881) );
  NAND2_X1 U978 ( .A1(G100), .A2(n899), .ZN(n880) );
  NAND2_X1 U979 ( .A1(n881), .A2(n880), .ZN(n885) );
  NAND2_X1 U980 ( .A1(n521), .A2(G136), .ZN(n883) );
  NAND2_X1 U981 ( .A1(G112), .A2(n896), .ZN(n882) );
  NAND2_X1 U982 ( .A1(n883), .A2(n882), .ZN(n884) );
  NOR2_X1 U983 ( .A1(n885), .A2(n884), .ZN(G162) );
  NAND2_X1 U984 ( .A1(G103), .A2(n899), .ZN(n887) );
  NAND2_X1 U985 ( .A1(G139), .A2(n521), .ZN(n886) );
  NAND2_X1 U986 ( .A1(n887), .A2(n886), .ZN(n893) );
  NAND2_X1 U987 ( .A1(G115), .A2(n896), .ZN(n888) );
  XOR2_X1 U988 ( .A(KEYINPUT119), .B(n888), .Z(n890) );
  NAND2_X1 U989 ( .A1(n895), .A2(G127), .ZN(n889) );
  NAND2_X1 U990 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U991 ( .A(KEYINPUT47), .B(n891), .Z(n892) );
  NOR2_X1 U992 ( .A1(n893), .A2(n892), .ZN(n956) );
  XNOR2_X1 U993 ( .A(n956), .B(n894), .ZN(n909) );
  NAND2_X1 U994 ( .A1(G130), .A2(n895), .ZN(n898) );
  NAND2_X1 U995 ( .A1(G118), .A2(n896), .ZN(n897) );
  NAND2_X1 U996 ( .A1(n898), .A2(n897), .ZN(n905) );
  NAND2_X1 U997 ( .A1(n899), .A2(G106), .ZN(n900) );
  XNOR2_X1 U998 ( .A(n900), .B(KEYINPUT118), .ZN(n902) );
  NAND2_X1 U999 ( .A1(G142), .A2(n521), .ZN(n901) );
  NAND2_X1 U1000 ( .A1(n902), .A2(n901), .ZN(n903) );
  XOR2_X1 U1001 ( .A(KEYINPUT45), .B(n903), .Z(n904) );
  NOR2_X1 U1002 ( .A1(n905), .A2(n904), .ZN(n907) );
  XOR2_X1 U1003 ( .A(G160), .B(n949), .Z(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n918) );
  XOR2_X1 U1006 ( .A(KEYINPUT48), .B(KEYINPUT120), .Z(n912) );
  XNOR2_X1 U1007 ( .A(n910), .B(KEYINPUT46), .ZN(n911) );
  XNOR2_X1 U1008 ( .A(n912), .B(n911), .ZN(n916) );
  XOR2_X1 U1009 ( .A(G164), .B(G162), .Z(n913) );
  XNOR2_X1 U1010 ( .A(n914), .B(n913), .ZN(n915) );
  XNOR2_X1 U1011 ( .A(n916), .B(n915), .ZN(n917) );
  XNOR2_X1 U1012 ( .A(n918), .B(n917), .ZN(n919) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n919), .ZN(G395) );
  XNOR2_X1 U1014 ( .A(n1014), .B(n920), .ZN(n922) );
  XNOR2_X1 U1015 ( .A(G171), .B(n1021), .ZN(n921) );
  XNOR2_X1 U1016 ( .A(n922), .B(n921), .ZN(n923) );
  XNOR2_X1 U1017 ( .A(n923), .B(G286), .ZN(n924) );
  NOR2_X1 U1018 ( .A1(G37), .A2(n924), .ZN(G397) );
  XNOR2_X1 U1019 ( .A(G2454), .B(G2427), .ZN(n934) );
  XOR2_X1 U1020 ( .A(G2430), .B(KEYINPUT114), .Z(n926) );
  XNOR2_X1 U1021 ( .A(G2443), .B(G2451), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(n926), .B(n925), .ZN(n930) );
  XOR2_X1 U1023 ( .A(G2446), .B(KEYINPUT113), .Z(n928) );
  XNOR2_X1 U1024 ( .A(G1348), .B(G1341), .ZN(n927) );
  XNOR2_X1 U1025 ( .A(n928), .B(n927), .ZN(n929) );
  XOR2_X1 U1026 ( .A(n930), .B(n929), .Z(n932) );
  XNOR2_X1 U1027 ( .A(G2435), .B(G2438), .ZN(n931) );
  XNOR2_X1 U1028 ( .A(n932), .B(n931), .ZN(n933) );
  XNOR2_X1 U1029 ( .A(n934), .B(n933), .ZN(n935) );
  NAND2_X1 U1030 ( .A1(n935), .A2(G14), .ZN(n942) );
  NAND2_X1 U1031 ( .A1(G319), .A2(n942), .ZN(n939) );
  NOR2_X1 U1032 ( .A1(G227), .A2(G229), .ZN(n936) );
  XOR2_X1 U1033 ( .A(KEYINPUT49), .B(n936), .Z(n937) );
  XNOR2_X1 U1034 ( .A(n937), .B(KEYINPUT121), .ZN(n938) );
  NOR2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n941) );
  NOR2_X1 U1036 ( .A1(G395), .A2(G397), .ZN(n940) );
  NAND2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(G225) );
  INV_X1 U1038 ( .A(G225), .ZN(G308) );
  INV_X1 U1039 ( .A(G57), .ZN(G237) );
  INV_X1 U1040 ( .A(n942), .ZN(G401) );
  XOR2_X1 U1041 ( .A(G2090), .B(G162), .Z(n943) );
  NOR2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1043 ( .A(n945), .B(KEYINPUT51), .ZN(n946) );
  NOR2_X1 U1044 ( .A1(n947), .A2(n946), .ZN(n955) );
  XOR2_X1 U1045 ( .A(G2084), .B(G160), .Z(n948) );
  NOR2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n951) );
  NAND2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n963) );
  XOR2_X1 U1050 ( .A(G2072), .B(n956), .Z(n958) );
  XOR2_X1 U1051 ( .A(G164), .B(G2078), .Z(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1053 ( .A(KEYINPUT50), .B(n959), .ZN(n961) );
  NAND2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(KEYINPUT52), .B(n964), .ZN(n965) );
  INV_X1 U1057 ( .A(KEYINPUT55), .ZN(n986) );
  NAND2_X1 U1058 ( .A1(n965), .A2(n986), .ZN(n966) );
  NAND2_X1 U1059 ( .A1(n966), .A2(G29), .ZN(n1043) );
  XOR2_X1 U1060 ( .A(KEYINPUT123), .B(KEYINPUT53), .Z(n979) );
  XNOR2_X1 U1061 ( .A(n967), .B(G27), .ZN(n971) );
  XNOR2_X1 U1062 ( .A(G2067), .B(G26), .ZN(n969) );
  XNOR2_X1 U1063 ( .A(G1996), .B(G32), .ZN(n968) );
  NOR2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n973) );
  XNOR2_X1 U1066 ( .A(G33), .B(G2072), .ZN(n972) );
  NOR2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  XOR2_X1 U1068 ( .A(KEYINPUT122), .B(n974), .Z(n976) );
  XNOR2_X1 U1069 ( .A(G1991), .B(G25), .ZN(n975) );
  NOR2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1071 ( .A1(n977), .A2(G28), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(n979), .B(n978), .ZN(n984) );
  XNOR2_X1 U1073 ( .A(G2084), .B(G34), .ZN(n980) );
  XNOR2_X1 U1074 ( .A(n980), .B(KEYINPUT54), .ZN(n982) );
  XNOR2_X1 U1075 ( .A(G35), .B(G2090), .ZN(n981) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(n986), .B(n985), .ZN(n988) );
  INV_X1 U1079 ( .A(G29), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1081 ( .A1(G11), .A2(n989), .ZN(n1041) );
  XOR2_X1 U1082 ( .A(G1348), .B(G4), .Z(n990) );
  XNOR2_X1 U1083 ( .A(KEYINPUT59), .B(n990), .ZN(n997) );
  XOR2_X1 U1084 ( .A(G1981), .B(G6), .Z(n994) );
  XNOR2_X1 U1085 ( .A(G1956), .B(G20), .ZN(n992) );
  XNOR2_X1 U1086 ( .A(G19), .B(G1341), .ZN(n991) );
  NOR2_X1 U1087 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1089 ( .A(KEYINPUT125), .B(n995), .Z(n996) );
  NOR2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1091 ( .A(KEYINPUT60), .B(n998), .ZN(n999) );
  XNOR2_X1 U1092 ( .A(n999), .B(KEYINPUT126), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(G1966), .B(G21), .ZN(n1001) );
  XNOR2_X1 U1094 ( .A(G1961), .B(G5), .ZN(n1000) );
  NOR2_X1 U1095 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1096 ( .A1(n1003), .A2(n1002), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(G1971), .B(G22), .ZN(n1005) );
  XNOR2_X1 U1098 ( .A(G23), .B(G1976), .ZN(n1004) );
  NOR2_X1 U1099 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  XOR2_X1 U1100 ( .A(G1986), .B(G24), .Z(n1006) );
  NAND2_X1 U1101 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1102 ( .A(KEYINPUT58), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1103 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1104 ( .A(KEYINPUT61), .B(n1011), .Z(n1012) );
  NOR2_X1 U1105 ( .A1(G16), .A2(n1012), .ZN(n1013) );
  XNOR2_X1 U1106 ( .A(KEYINPUT127), .B(n1013), .ZN(n1039) );
  XNOR2_X1 U1107 ( .A(KEYINPUT56), .B(G16), .ZN(n1037) );
  XNOR2_X1 U1108 ( .A(G301), .B(G1961), .ZN(n1016) );
  XNOR2_X1 U1109 ( .A(n1014), .B(G1341), .ZN(n1015) );
  NOR2_X1 U1110 ( .A1(n1016), .A2(n1015), .ZN(n1035) );
  NAND2_X1 U1111 ( .A1(G1971), .A2(G303), .ZN(n1017) );
  NAND2_X1 U1112 ( .A1(n1018), .A2(n1017), .ZN(n1025) );
  NOR2_X1 U1113 ( .A1(n1020), .A2(n1019), .ZN(n1023) );
  XOR2_X1 U1114 ( .A(n1021), .B(G1348), .Z(n1022) );
  NAND2_X1 U1115 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1116 ( .A1(n1025), .A2(n1024), .ZN(n1031) );
  XOR2_X1 U1117 ( .A(G1966), .B(G168), .Z(n1026) );
  XNOR2_X1 U1118 ( .A(KEYINPUT124), .B(n1026), .ZN(n1027) );
  NOR2_X1 U1119 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1120 ( .A(KEYINPUT57), .B(n1029), .Z(n1030) );
  NAND2_X1 U1121 ( .A1(n1031), .A2(n1030), .ZN(n1033) );
  XNOR2_X1 U1122 ( .A(G1956), .B(G299), .ZN(n1032) );
  NOR2_X1 U1123 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1124 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1125 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NAND2_X1 U1126 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  NOR2_X1 U1127 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  NAND2_X1 U1128 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  XOR2_X1 U1129 ( .A(KEYINPUT62), .B(n1044), .Z(G311) );
  INV_X1 U1130 ( .A(G311), .ZN(G150) );
endmodule

