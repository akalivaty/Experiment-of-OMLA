//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n626, new_n627, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n797, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT93), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G1gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n204), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n208), .B1(new_n207), .B2(new_n206), .ZN(new_n209));
  INV_X1    g008(.A(G8gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G57gat), .ZN(new_n213));
  OR3_X1    g012(.A1(new_n213), .A2(KEYINPUT95), .A3(G64gat), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT95), .B1(new_n213), .B2(G64gat), .ZN(new_n215));
  INV_X1    g014(.A(G64gat), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n214), .B(new_n215), .C1(G57gat), .C2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G71gat), .A2(G78gat), .ZN(new_n218));
  OR2_X1    g017(.A1(G71gat), .A2(G78gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT9), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  XOR2_X1   g021(.A(new_n222), .B(KEYINPUT96), .Z(new_n223));
  XNOR2_X1  g022(.A(G57gat), .B(G64gat), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n218), .B(new_n219), .C1(new_n224), .C2(new_n220), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(KEYINPUT21), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n212), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G183gat), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n227), .B(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G231gat), .A2(G233gat), .ZN(new_n230));
  XOR2_X1   g029(.A(new_n229), .B(new_n230), .Z(new_n231));
  XNOR2_X1  g030(.A(G127gat), .B(G155gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n232), .B(G211gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n231), .B(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT21), .B1(new_n223), .B2(new_n225), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g036(.A(new_n234), .B(new_n237), .Z(new_n238));
  INV_X1    g037(.A(KEYINPUT92), .ZN(new_n239));
  OR3_X1    g038(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G43gat), .B(G50gat), .ZN(new_n243));
  INV_X1    g042(.A(G36gat), .ZN(new_n244));
  XOR2_X1   g043(.A(KEYINPUT91), .B(G29gat), .Z(new_n245));
  OAI221_X1 g044(.A(new_n242), .B1(KEYINPUT15), .B2(new_n243), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n243), .A2(KEYINPUT15), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n246), .B(new_n247), .Z(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT17), .ZN(new_n249));
  NAND2_X1  g048(.A1(G85gat), .A2(G92gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT99), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(KEYINPUT7), .ZN(new_n252));
  NAND2_X1  g051(.A1(G99gat), .A2(G106gat), .ZN(new_n253));
  INV_X1    g052(.A(G85gat), .ZN(new_n254));
  INV_X1    g053(.A(G92gat), .ZN(new_n255));
  AOI22_X1  g054(.A1(KEYINPUT8), .A2(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G99gat), .B(G106gat), .ZN(new_n258));
  XOR2_X1   g057(.A(new_n257), .B(new_n258), .Z(new_n259));
  NAND2_X1  g058(.A1(new_n249), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n259), .ZN(new_n261));
  AND2_X1   g060(.A1(G232gat), .A2(G233gat), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n261), .A2(new_n248), .B1(KEYINPUT41), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(KEYINPUT97), .ZN(new_n265));
  XOR2_X1   g064(.A(KEYINPUT98), .B(KEYINPUT100), .Z(new_n266));
  XNOR2_X1  g065(.A(G134gat), .B(G162gat), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n266), .B(new_n267), .Z(new_n268));
  XNOR2_X1  g067(.A(new_n265), .B(new_n268), .ZN(new_n269));
  XOR2_X1   g068(.A(G190gat), .B(G218gat), .Z(new_n270));
  NOR2_X1   g069(.A1(new_n262), .A2(KEYINPUT41), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n269), .B(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n223), .A2(new_n225), .ZN(new_n274));
  OR2_X1    g073(.A1(new_n259), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT101), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT10), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n259), .A2(new_n274), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n275), .A2(new_n276), .A3(KEYINPUT10), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  AND2_X1   g081(.A1(G230gat), .A2(G233gat), .ZN(new_n283));
  OR2_X1    g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n275), .A2(new_n280), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(new_n283), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G120gat), .B(G148gat), .ZN(new_n288));
  INV_X1    g087(.A(G176gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  XOR2_X1   g089(.A(new_n290), .B(G204gat), .Z(new_n291));
  AND2_X1   g090(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n287), .A2(new_n291), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NOR3_X1   g093(.A1(new_n238), .A2(new_n273), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT3), .ZN(new_n296));
  XNOR2_X1  g095(.A(G197gat), .B(G204gat), .ZN(new_n297));
  INV_X1    g096(.A(G211gat), .ZN(new_n298));
  INV_X1    g097(.A(G218gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n297), .B1(KEYINPUT22), .B2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G211gat), .B(G218gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n296), .B1(new_n303), .B2(KEYINPUT29), .ZN(new_n304));
  INV_X1    g103(.A(G141gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G148gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT74), .ZN(new_n307));
  INV_X1    g106(.A(G148gat), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n307), .B1(G141gat), .B2(new_n308), .ZN(new_n309));
  NOR3_X1   g108(.A1(new_n305), .A2(KEYINPUT74), .A3(G148gat), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n306), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT75), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OAI211_X1 g112(.A(KEYINPUT75), .B(new_n306), .C1(new_n309), .C2(new_n310), .ZN(new_n314));
  NAND2_X1  g113(.A1(G155gat), .A2(G162gat), .ZN(new_n315));
  OR2_X1    g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n315), .B1(new_n316), .B2(KEYINPUT2), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n313), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n308), .A2(G141gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n306), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT73), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n315), .A2(KEYINPUT2), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n306), .A2(new_n319), .A3(KEYINPUT73), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  OR2_X1    g124(.A1(new_n315), .A2(KEYINPUT72), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n315), .A2(KEYINPUT72), .ZN(new_n327));
  AND3_X1   g126(.A1(new_n326), .A2(new_n316), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n318), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n304), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n318), .A2(new_n296), .A3(new_n329), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT76), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n318), .A2(KEYINPUT76), .A3(new_n329), .A4(new_n296), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT29), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n303), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n331), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G228gat), .A2(G233gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n339), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n341), .B(new_n331), .C1(new_n336), .C2(new_n337), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  XOR2_X1   g142(.A(G78gat), .B(G106gat), .Z(new_n344));
  XNOR2_X1  g143(.A(new_n344), .B(KEYINPUT31), .ZN(new_n345));
  INV_X1    g144(.A(G50gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n345), .B(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(G22gat), .B1(new_n343), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT83), .B1(new_n343), .B2(new_n347), .ZN(new_n349));
  INV_X1    g148(.A(G22gat), .ZN(new_n350));
  INV_X1    g149(.A(new_n347), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n340), .A2(new_n350), .A3(new_n342), .A4(new_n351), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n348), .A2(new_n349), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n349), .B1(new_n348), .B2(new_n352), .ZN(new_n354));
  OR2_X1    g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G15gat), .B(G43gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(G71gat), .B(G99gat), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n356), .B(new_n357), .Z(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G183gat), .A2(G190gat), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(G169gat), .A2(G176gat), .ZN(new_n362));
  OR3_X1    g161(.A1(new_n361), .A2(new_n362), .A3(KEYINPUT67), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT26), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT67), .B1(new_n361), .B2(new_n362), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n363), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT66), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT27), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n369), .A2(G183gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n228), .A2(KEYINPUT27), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n368), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n228), .A2(KEYINPUT27), .ZN(new_n373));
  AOI21_X1  g172(.A(G190gat), .B1(new_n373), .B2(KEYINPUT66), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT28), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT27), .B(G183gat), .ZN(new_n376));
  INV_X1    g175(.A(G190gat), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n376), .A2(KEYINPUT28), .A3(new_n377), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n360), .B(new_n367), .C1(new_n375), .C2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NOR3_X1   g180(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT25), .B1(new_n383), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT23), .ZN(new_n389));
  INV_X1    g188(.A(G169gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(new_n390), .A3(new_n289), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(G169gat), .A2(G176gat), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT24), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n360), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n228), .A2(new_n377), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(new_n398), .A3(new_n384), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n399), .A2(new_n393), .A3(new_n394), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n388), .A2(new_n395), .B1(new_n400), .B2(KEYINPUT25), .ZN(new_n401));
  AND2_X1   g200(.A1(new_n379), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT68), .ZN(new_n403));
  XNOR2_X1  g202(.A(G113gat), .B(G120gat), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n403), .B1(new_n404), .B2(KEYINPUT1), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT1), .ZN(new_n406));
  INV_X1    g205(.A(G113gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n407), .A2(G120gat), .ZN(new_n408));
  INV_X1    g207(.A(G120gat), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n409), .A2(G113gat), .ZN(new_n410));
  OAI211_X1 g209(.A(KEYINPUT68), .B(new_n406), .C1(new_n408), .C2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G127gat), .B(G134gat), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n405), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n403), .B(new_n412), .C1(new_n404), .C2(KEYINPUT1), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(G227gat), .A2(G233gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT64), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n379), .A2(new_n401), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n416), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n418), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT33), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n359), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n423), .A2(KEYINPUT32), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n418), .A2(new_n422), .ZN(new_n428));
  INV_X1    g227(.A(new_n420), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(KEYINPUT34), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT69), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n427), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n432), .B1(new_n427), .B2(new_n433), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n355), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G1gat), .B(G29gat), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT79), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  XOR2_X1   g239(.A(G57gat), .B(G85gat), .Z(new_n441));
  XNOR2_X1  g240(.A(new_n440), .B(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n442), .B(new_n443), .ZN(new_n444));
  XOR2_X1   g243(.A(KEYINPUT77), .B(KEYINPUT5), .Z(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n330), .A2(new_n417), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n416), .A2(new_n318), .A3(new_n329), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(G225gat), .A2(G233gat), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n446), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n334), .A2(new_n335), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n330), .A2(KEYINPUT3), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n453), .A2(new_n417), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n448), .A2(KEYINPUT4), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT4), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n416), .A2(new_n318), .A3(new_n457), .A4(new_n329), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n450), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n452), .B1(new_n455), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n458), .A2(KEYINPUT80), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT81), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n448), .A2(new_n464), .A3(KEYINPUT4), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n464), .B1(new_n448), .B2(KEYINPUT4), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n456), .A2(KEYINPUT81), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n448), .A2(new_n464), .A3(KEYINPUT4), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(new_n462), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n453), .A2(new_n417), .A3(new_n454), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n445), .A2(new_n451), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n467), .A2(new_n470), .A3(new_n471), .A4(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n444), .B1(new_n461), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT6), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n461), .A2(new_n473), .A3(new_n444), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT6), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n475), .B1(new_n478), .B2(new_n474), .ZN(new_n479));
  XNOR2_X1  g278(.A(G8gat), .B(G36gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n480), .B(new_n216), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n481), .B(new_n255), .ZN(new_n482));
  NAND2_X1  g281(.A1(G226gat), .A2(G233gat), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT70), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n421), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n379), .A2(new_n401), .A3(KEYINPUT70), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n483), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n488), .A2(KEYINPUT29), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n421), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n303), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n485), .A2(new_n486), .A3(new_n489), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n402), .A2(new_n488), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n492), .A2(new_n337), .A3(new_n493), .ZN(new_n494));
  AOI211_X1 g293(.A(KEYINPUT30), .B(new_n482), .C1(new_n491), .C2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n482), .B(KEYINPUT71), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n491), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT30), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n482), .B1(new_n491), .B2(new_n494), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n496), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n479), .A2(KEYINPUT82), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT82), .B1(new_n479), .B2(new_n501), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n437), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT35), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n444), .B(KEYINPUT84), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n507), .B1(new_n461), .B2(new_n473), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT87), .B1(new_n478), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n461), .A2(new_n473), .ZN(new_n510));
  INV_X1    g309(.A(new_n507), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT87), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n512), .A2(new_n513), .A3(new_n477), .A4(new_n476), .ZN(new_n514));
  AND3_X1   g313(.A1(new_n509), .A2(new_n475), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT30), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n492), .A2(new_n337), .A3(new_n493), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n379), .A2(new_n401), .A3(KEYINPUT70), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT70), .B1(new_n379), .B2(new_n401), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n488), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n421), .A2(new_n489), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n337), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n516), .B1(new_n523), .B2(new_n497), .ZN(new_n524));
  INV_X1    g323(.A(new_n500), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n495), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR3_X1   g325(.A1(new_n515), .A2(KEYINPUT35), .A3(new_n526), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n432), .A2(new_n427), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n432), .A2(new_n427), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n355), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n506), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n353), .A2(new_n354), .ZN(new_n535));
  NOR3_X1   g334(.A1(new_n502), .A2(new_n535), .A3(new_n503), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT85), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n537), .A2(KEYINPUT40), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT39), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n449), .A2(new_n451), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n467), .A2(new_n470), .A3(new_n471), .ZN(new_n541));
  AOI211_X1 g340(.A(new_n539), .B(new_n540), .C1(new_n541), .C2(new_n451), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(new_n539), .A3(new_n451), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(new_n507), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n538), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n541), .A2(new_n451), .ZN(new_n546));
  INV_X1    g345(.A(new_n540), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(KEYINPUT39), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n538), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n548), .A2(new_n549), .A3(new_n543), .A4(new_n507), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n545), .A2(new_n550), .A3(new_n526), .A4(new_n512), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT86), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n548), .A2(new_n543), .A3(new_n507), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n508), .B1(new_n553), .B2(new_n538), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT86), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n554), .A2(new_n555), .A3(new_n526), .A4(new_n550), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n485), .A2(new_n486), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n490), .B1(new_n557), .B2(new_n488), .ZN(new_n558));
  OAI211_X1 g357(.A(KEYINPUT37), .B(new_n494), .C1(new_n558), .C2(new_n337), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n559), .A2(KEYINPUT88), .A3(new_n482), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT37), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n561), .B1(new_n517), .B2(new_n522), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT88), .B1(new_n559), .B2(new_n482), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT38), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT89), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g366(.A(KEYINPUT89), .B(KEYINPUT38), .C1(new_n563), .C2(new_n564), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n558), .A2(new_n337), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n492), .A2(new_n493), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n570), .B(KEYINPUT37), .C1(new_n337), .C2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT38), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n572), .A2(new_n573), .A3(new_n497), .A4(new_n562), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n574), .A2(new_n525), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n575), .A2(new_n475), .A3(new_n509), .A4(new_n514), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n552), .B(new_n556), .C1(new_n569), .C2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n536), .B1(new_n577), .B2(new_n535), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT36), .B1(new_n434), .B2(new_n435), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT36), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n528), .A2(new_n580), .A3(new_n529), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n534), .B1(new_n578), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n211), .A2(new_n248), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT94), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n249), .A2(new_n212), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G229gat), .A2(G233gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT18), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n586), .B1(new_n211), .B2(new_n248), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n589), .B(KEYINPUT13), .Z(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G113gat), .B(G141gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(G169gat), .B(G197gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n600), .B(KEYINPUT12), .Z(new_n601));
  OR2_X1    g400(.A1(new_n595), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n595), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n295), .A2(new_n583), .A3(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n605), .A2(new_n479), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(new_n207), .ZN(G1324gat));
  OR2_X1    g406(.A1(new_n605), .A2(new_n501), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n203), .A2(new_n210), .ZN(new_n609));
  NOR2_X1   g408(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n610));
  NOR3_X1   g409(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n611), .A2(KEYINPUT42), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT102), .ZN(new_n613));
  AOI22_X1  g412(.A1(new_n611), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n608), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(G1325gat));
  INV_X1    g414(.A(G15gat), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n616), .B1(new_n605), .B2(new_n531), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n617), .B(KEYINPUT103), .Z(new_n618));
  INV_X1    g417(.A(KEYINPUT104), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n579), .A2(new_n619), .A3(new_n581), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n619), .B1(new_n579), .B2(new_n581), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NOR3_X1   g422(.A1(new_n605), .A2(new_n616), .A3(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n618), .A2(new_n624), .ZN(G1326gat));
  NOR2_X1   g424(.A1(new_n605), .A2(new_n535), .ZN(new_n626));
  XOR2_X1   g425(.A(KEYINPUT43), .B(G22gat), .Z(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(G1327gat));
  INV_X1    g427(.A(new_n238), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n629), .A2(new_n294), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n604), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n583), .A2(new_n273), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n479), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n637), .A2(new_n638), .A3(new_n245), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT45), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT108), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n634), .A2(KEYINPUT44), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n577), .A2(new_n535), .ZN(new_n644));
  INV_X1    g443(.A(new_n536), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT106), .B1(new_n646), .B2(new_n623), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT106), .ZN(new_n648));
  NOR3_X1   g447(.A1(new_n578), .A2(new_n648), .A3(new_n622), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n534), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT44), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n650), .A2(new_n651), .A3(new_n273), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT107), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n273), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n552), .A2(new_n556), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n515), .A2(new_n575), .A3(new_n567), .A4(new_n568), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n355), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI211_X1 g457(.A(KEYINPUT106), .B(new_n623), .C1(new_n658), .C2(new_n536), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n648), .B1(new_n578), .B2(new_n622), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n655), .B1(new_n661), .B2(new_n534), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n662), .A2(KEYINPUT107), .A3(new_n651), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n643), .B1(new_n654), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n604), .B(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n631), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n641), .B1(new_n664), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(KEYINPUT107), .B1(new_n662), .B2(new_n651), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n506), .A2(new_n533), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n672), .B1(new_n659), .B2(new_n660), .ZN(new_n673));
  NOR4_X1   g472(.A1(new_n673), .A2(new_n653), .A3(KEYINPUT44), .A4(new_n655), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n642), .B1(new_n671), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n675), .A2(KEYINPUT108), .A3(new_n668), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n670), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n678), .A2(new_n479), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n640), .B1(new_n679), .B2(new_n245), .ZN(G1328gat));
  NAND3_X1  g479(.A1(new_n637), .A2(new_n244), .A3(new_n526), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT109), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT46), .ZN(new_n683));
  OAI21_X1  g482(.A(G36gat), .B1(new_n678), .B2(new_n501), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(G1329gat));
  AOI21_X1  g484(.A(new_n623), .B1(new_n670), .B2(new_n676), .ZN(new_n686));
  INV_X1    g485(.A(G43gat), .ZN(new_n687));
  OAI21_X1  g486(.A(KEYINPUT110), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n664), .A2(new_n641), .A3(new_n669), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT108), .B1(new_n675), .B2(new_n668), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n622), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT110), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(new_n692), .A3(G43gat), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n636), .A2(G43gat), .A3(new_n531), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n694), .A2(KEYINPUT47), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n688), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT111), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n664), .A2(new_n669), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n687), .B1(new_n698), .B2(new_n622), .ZN(new_n699));
  OAI21_X1  g498(.A(KEYINPUT47), .B1(new_n699), .B2(new_n694), .ZN(new_n700));
  AND3_X1   g499(.A1(new_n696), .A2(new_n697), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n697), .B1(new_n696), .B2(new_n700), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(G1330gat));
  NOR3_X1   g502(.A1(new_n636), .A2(G50gat), .A3(new_n535), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n698), .A2(new_n355), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n704), .B1(new_n705), .B2(G50gat), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(KEYINPUT48), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n677), .A2(new_n355), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n704), .B1(new_n708), .B2(G50gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n707), .B1(new_n709), .B2(new_n710), .ZN(G1331gat));
  INV_X1    g510(.A(new_n294), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n666), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n713), .A2(new_n650), .A3(new_n629), .A4(new_n655), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n714), .A2(new_n479), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(new_n213), .ZN(G1332gat));
  AOI211_X1 g515(.A(new_n501), .B(new_n714), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT113), .ZN(new_n718));
  NOR2_X1   g517(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1333gat));
  OAI21_X1  g519(.A(G71gat), .B1(new_n714), .B2(new_n623), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n714), .A2(G71gat), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n722), .B2(new_n531), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n723), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g523(.A1(new_n714), .A2(new_n535), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n725), .B(G78gat), .Z(G1335gat));
  NAND2_X1  g525(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n727));
  XNOR2_X1  g526(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n728));
  NOR4_X1   g527(.A1(new_n673), .A2(new_n666), .A3(new_n629), .A4(new_n655), .ZN(new_n729));
  MUX2_X1   g528(.A(new_n727), .B(new_n728), .S(new_n729), .Z(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT115), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n294), .A2(new_n254), .A3(new_n638), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n675), .A2(new_n238), .A3(new_n713), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n733), .A2(new_n638), .ZN(new_n734));
  OAI22_X1  g533(.A1(new_n731), .A2(new_n732), .B1(new_n254), .B2(new_n734), .ZN(G1336gat));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n526), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G92gat), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n712), .A2(G92gat), .A3(new_n501), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT52), .B1(new_n730), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n729), .A2(KEYINPUT116), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n741), .B(KEYINPUT51), .Z(new_n742));
  AOI22_X1  g541(.A1(G92gat), .A2(new_n736), .B1(new_n742), .B2(new_n738), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT52), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n740), .B1(new_n743), .B2(new_n744), .ZN(G1337gat));
  NAND2_X1  g544(.A1(new_n733), .A2(new_n622), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(G99gat), .ZN(new_n747));
  OR3_X1    g546(.A1(new_n712), .A2(G99gat), .A3(new_n531), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n731), .B2(new_n748), .ZN(G1338gat));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n355), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(G106gat), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n712), .A2(G106gat), .A3(new_n535), .ZN(new_n752));
  AOI21_X1  g551(.A(KEYINPUT53), .B1(new_n730), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  AOI22_X1  g553(.A1(G106gat), .A2(new_n750), .B1(new_n742), .B2(new_n752), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT53), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(G1339gat));
  NAND2_X1  g556(.A1(new_n282), .A2(new_n283), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n284), .A2(KEYINPUT54), .A3(new_n758), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n759), .B(new_n291), .C1(KEYINPUT54), .C2(new_n284), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT55), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n762), .A2(new_n763), .A3(new_n293), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n666), .A2(new_n764), .ZN(new_n765));
  OAI22_X1  g564(.A1(new_n588), .A2(new_n589), .B1(new_n592), .B2(new_n593), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n600), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n294), .A2(new_n602), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT117), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n273), .B1(new_n765), .B2(new_n769), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n602), .A2(new_n767), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n764), .A2(new_n273), .A3(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n238), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n667), .A2(new_n295), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT118), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n479), .A2(new_n526), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n774), .A2(KEYINPUT118), .A3(new_n775), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n532), .ZN(new_n782));
  OAI21_X1  g581(.A(G113gat), .B1(new_n782), .B2(new_n632), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n437), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n666), .A2(new_n407), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(KEYINPUT119), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n783), .B1(new_n784), .B2(new_n786), .ZN(G1340gat));
  NAND3_X1  g586(.A1(new_n781), .A2(new_n532), .A3(new_n294), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT120), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n788), .A2(new_n789), .A3(G120gat), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n789), .B1(new_n788), .B2(G120gat), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n294), .A2(new_n409), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT121), .ZN(new_n794));
  OAI22_X1  g593(.A1(new_n791), .A2(new_n792), .B1(new_n784), .B2(new_n794), .ZN(G1341gat));
  INV_X1    g594(.A(G127gat), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n796), .B1(new_n784), .B2(new_n238), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n781), .A2(G127gat), .A3(new_n532), .A4(new_n629), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(G1342gat));
  NOR3_X1   g598(.A1(new_n784), .A2(G134gat), .A3(new_n655), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT56), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  OAI21_X1  g602(.A(G134gat), .B1(new_n782), .B2(new_n655), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(G1343gat));
  NAND2_X1  g604(.A1(new_n623), .A2(new_n779), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n764), .A2(new_n604), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n273), .B1(new_n807), .B2(new_n768), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n238), .B1(new_n808), .B2(new_n773), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n775), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n355), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n806), .B1(new_n811), .B2(KEYINPUT57), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n778), .A2(new_n355), .A3(new_n780), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n812), .B1(new_n813), .B2(KEYINPUT57), .ZN(new_n814));
  OAI21_X1  g613(.A(G141gat), .B1(new_n814), .B2(new_n632), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT58), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n813), .A2(new_n806), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(new_n305), .A3(new_n604), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n815), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(G141gat), .B1(new_n814), .B2(new_n667), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n820), .A2(new_n818), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n821), .B2(new_n816), .ZN(G1344gat));
  INV_X1    g621(.A(KEYINPUT59), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(new_n814), .B2(new_n712), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n295), .A2(new_n632), .ZN(new_n825));
  AOI211_X1 g624(.A(KEYINPUT57), .B(new_n535), .C1(new_n809), .C2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n826), .B1(new_n813), .B2(KEYINPUT57), .ZN(new_n827));
  INV_X1    g626(.A(new_n806), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n823), .B1(new_n828), .B2(KEYINPUT122), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n827), .A2(new_n294), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n828), .A2(KEYINPUT122), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n824), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(G148gat), .B1(new_n817), .B2(new_n294), .ZN(new_n833));
  AOI22_X1  g632(.A1(new_n832), .A2(G148gat), .B1(KEYINPUT59), .B2(new_n833), .ZN(G1345gat));
  AOI21_X1  g633(.A(G155gat), .B1(new_n817), .B2(new_n629), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n814), .A2(new_n238), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n835), .B1(new_n836), .B2(G155gat), .ZN(G1346gat));
  INV_X1    g636(.A(G162gat), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n814), .A2(new_n838), .A3(new_n655), .ZN(new_n839));
  AOI21_X1  g638(.A(G162gat), .B1(new_n817), .B2(new_n273), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(G1347gat));
  AND3_X1   g640(.A1(new_n774), .A2(KEYINPUT118), .A3(new_n775), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT118), .B1(new_n774), .B2(new_n775), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n355), .A2(new_n501), .A3(new_n436), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n844), .A2(KEYINPUT123), .A3(new_n479), .A4(new_n845), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n778), .A2(new_n479), .A3(new_n780), .A4(new_n845), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT123), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n846), .A2(new_n849), .A3(new_n390), .A4(new_n666), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n844), .A2(new_n479), .A3(new_n526), .A4(new_n532), .ZN(new_n851));
  OAI21_X1  g650(.A(G169gat), .B1(new_n851), .B2(new_n632), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(G1348gat));
  NAND4_X1  g652(.A1(new_n846), .A2(new_n849), .A3(new_n289), .A4(new_n294), .ZN(new_n854));
  OAI21_X1  g653(.A(G176gat), .B1(new_n851), .B2(new_n712), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(KEYINPUT124), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT124), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n854), .A2(new_n855), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(G1349gat));
  OAI21_X1  g659(.A(G183gat), .B1(new_n851), .B2(new_n238), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n629), .A2(new_n376), .ZN(new_n862));
  OR2_X1    g661(.A1(new_n847), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  AND2_X1   g663(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n864), .B(new_n865), .ZN(G1350gat));
  OAI21_X1  g665(.A(G190gat), .B1(new_n851), .B2(new_n655), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT61), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT61), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n869), .B(G190gat), .C1(new_n851), .C2(new_n655), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n846), .A2(new_n849), .A3(new_n377), .A4(new_n273), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n872), .A2(KEYINPUT126), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n872), .A2(KEYINPUT126), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n871), .B1(new_n873), .B2(new_n874), .ZN(G1351gat));
  NOR3_X1   g674(.A1(new_n622), .A2(new_n638), .A3(new_n501), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n827), .A2(new_n604), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(G197gat), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n842), .A2(new_n843), .A3(new_n535), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n876), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n880), .A2(G197gat), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n878), .B1(new_n667), .B2(new_n881), .ZN(G1352gat));
  XNOR2_X1  g681(.A(KEYINPUT127), .B(G204gat), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n880), .A2(new_n712), .A3(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT62), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n827), .A2(new_n294), .A3(new_n876), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(new_n883), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n884), .A2(new_n885), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n886), .A2(new_n888), .A3(new_n889), .ZN(G1353gat));
  INV_X1    g689(.A(new_n880), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n298), .A3(new_n629), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n827), .A2(new_n629), .A3(new_n876), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n893), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT63), .B1(new_n893), .B2(G211gat), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(G1354gat));
  NAND3_X1  g695(.A1(new_n891), .A2(new_n299), .A3(new_n273), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n827), .A2(new_n273), .A3(new_n876), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n897), .B1(new_n898), .B2(new_n299), .ZN(G1355gat));
endmodule


