

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582;

  AND2_X1 U324 ( .A1(G230GAT), .A2(G233GAT), .ZN(n292) );
  XOR2_X1 U325 ( .A(G183GAT), .B(KEYINPUT17), .Z(n293) );
  NOR2_X1 U326 ( .A1(n449), .A2(n553), .ZN(n450) );
  OR2_X1 U327 ( .A1(n541), .A2(n569), .ZN(n357) );
  XNOR2_X1 U328 ( .A(n368), .B(n292), .ZN(n329) );
  XNOR2_X1 U329 ( .A(n329), .B(n408), .ZN(n331) );
  INV_X1 U330 ( .A(KEYINPUT95), .ZN(n300) );
  XNOR2_X1 U331 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U332 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U333 ( .A(n335), .B(n334), .ZN(n337) );
  XNOR2_X1 U334 ( .A(n484), .B(KEYINPUT105), .ZN(n485) );
  NOR2_X1 U335 ( .A1(n552), .A2(n454), .ZN(n445) );
  NOR2_X1 U336 ( .A1(n513), .A2(n487), .ZN(n489) );
  INV_X1 U337 ( .A(G218GAT), .ZN(n446) );
  XOR2_X1 U338 ( .A(KEYINPUT41), .B(n574), .Z(n541) );
  XNOR2_X1 U339 ( .A(n489), .B(n488), .ZN(n496) );
  XNOR2_X1 U340 ( .A(n446), .B(KEYINPUT62), .ZN(n447) );
  XNOR2_X1 U341 ( .A(n448), .B(n447), .ZN(G1355GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT21), .B(KEYINPUT90), .Z(n295) );
  XNOR2_X1 U343 ( .A(G218GAT), .B(KEYINPUT91), .ZN(n294) );
  XNOR2_X1 U344 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U345 ( .A(n296), .B(G211GAT), .Z(n298) );
  XNOR2_X1 U346 ( .A(G197GAT), .B(G204GAT), .ZN(n297) );
  XNOR2_X1 U347 ( .A(n298), .B(n297), .ZN(n422) );
  XNOR2_X1 U348 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n299) );
  XNOR2_X1 U349 ( .A(n293), .B(n299), .ZN(n434) );
  NAND2_X1 U350 ( .A1(G226GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U351 ( .A(n434), .B(n302), .ZN(n306) );
  XOR2_X1 U352 ( .A(G92GAT), .B(G8GAT), .Z(n304) );
  XNOR2_X1 U353 ( .A(G169GAT), .B(G36GAT), .ZN(n303) );
  XNOR2_X1 U354 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U355 ( .A(n306), .B(n305), .Z(n308) );
  XOR2_X1 U356 ( .A(G190GAT), .B(KEYINPUT71), .Z(n364) );
  XOR2_X1 U357 ( .A(G176GAT), .B(G64GAT), .Z(n330) );
  XNOR2_X1 U358 ( .A(n364), .B(n330), .ZN(n307) );
  XNOR2_X1 U359 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U360 ( .A(n422), .B(n309), .ZN(n515) );
  XOR2_X1 U361 ( .A(G64GAT), .B(G57GAT), .Z(n311) );
  XNOR2_X1 U362 ( .A(G1GAT), .B(G8GAT), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U364 ( .A(KEYINPUT15), .B(KEYINPUT75), .Z(n313) );
  XNOR2_X1 U365 ( .A(KEYINPUT12), .B(KEYINPUT14), .ZN(n312) );
  XNOR2_X1 U366 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U367 ( .A(n315), .B(n314), .ZN(n328) );
  XOR2_X1 U368 ( .A(G183GAT), .B(G71GAT), .Z(n317) );
  XNOR2_X1 U369 ( .A(G15GAT), .B(G127GAT), .ZN(n316) );
  XNOR2_X1 U370 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U371 ( .A(G78GAT), .B(G155GAT), .Z(n319) );
  XNOR2_X1 U372 ( .A(G22GAT), .B(G211GAT), .ZN(n318) );
  XNOR2_X1 U373 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U374 ( .A(n321), .B(n320), .Z(n326) );
  XOR2_X1 U375 ( .A(KEYINPUT13), .B(KEYINPUT68), .Z(n332) );
  XOR2_X1 U376 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n323) );
  NAND2_X1 U377 ( .A1(G231GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U378 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U379 ( .A(n332), .B(n324), .ZN(n325) );
  XNOR2_X1 U380 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U381 ( .A(n328), .B(n327), .Z(n578) );
  XNOR2_X1 U382 ( .A(KEYINPUT46), .B(KEYINPUT114), .ZN(n358) );
  XOR2_X1 U383 ( .A(G85GAT), .B(G92GAT), .Z(n368) );
  XOR2_X1 U384 ( .A(G106GAT), .B(G78GAT), .Z(n408) );
  XNOR2_X1 U385 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U386 ( .A(G99GAT), .B(G71GAT), .Z(n435) );
  XOR2_X1 U387 ( .A(G148GAT), .B(G57GAT), .Z(n390) );
  XOR2_X1 U388 ( .A(n435), .B(n390), .Z(n333) );
  XOR2_X1 U389 ( .A(G120GAT), .B(G204GAT), .Z(n336) );
  XNOR2_X1 U390 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U391 ( .A(KEYINPUT33), .B(KEYINPUT69), .Z(n339) );
  XNOR2_X1 U392 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n338) );
  XNOR2_X1 U393 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U394 ( .A(n341), .B(n340), .ZN(n574) );
  XOR2_X1 U395 ( .A(KEYINPUT64), .B(KEYINPUT30), .Z(n343) );
  XNOR2_X1 U396 ( .A(KEYINPUT65), .B(KEYINPUT29), .ZN(n342) );
  XNOR2_X1 U397 ( .A(n343), .B(n342), .ZN(n352) );
  XOR2_X1 U398 ( .A(G15GAT), .B(G113GAT), .Z(n345) );
  XNOR2_X1 U399 ( .A(G169GAT), .B(G43GAT), .ZN(n344) );
  XNOR2_X1 U400 ( .A(n345), .B(n344), .ZN(n431) );
  XOR2_X1 U401 ( .A(G141GAT), .B(G22GAT), .Z(n409) );
  XOR2_X1 U402 ( .A(n431), .B(n409), .Z(n347) );
  NAND2_X1 U403 ( .A1(G229GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U404 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U405 ( .A(n348), .B(G8GAT), .Z(n350) );
  XOR2_X1 U406 ( .A(G29GAT), .B(G1GAT), .Z(n391) );
  XNOR2_X1 U407 ( .A(G197GAT), .B(n391), .ZN(n349) );
  XNOR2_X1 U408 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U409 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U410 ( .A(KEYINPUT8), .B(KEYINPUT66), .Z(n354) );
  XNOR2_X1 U411 ( .A(G50GAT), .B(G36GAT), .ZN(n353) );
  XNOR2_X1 U412 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U413 ( .A(KEYINPUT7), .B(n355), .Z(n373) );
  XOR2_X1 U414 ( .A(n356), .B(n373), .Z(n569) );
  XNOR2_X1 U415 ( .A(n358), .B(n357), .ZN(n359) );
  AND2_X1 U416 ( .A1(n578), .A2(n359), .ZN(n379) );
  XOR2_X1 U417 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n361) );
  XNOR2_X1 U418 ( .A(G134GAT), .B(G162GAT), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n361), .B(n360), .ZN(n378) );
  XOR2_X1 U420 ( .A(KEYINPUT72), .B(KEYINPUT11), .Z(n363) );
  XNOR2_X1 U421 ( .A(G218GAT), .B(KEYINPUT70), .ZN(n362) );
  XNOR2_X1 U422 ( .A(n363), .B(n362), .ZN(n365) );
  XOR2_X1 U423 ( .A(n365), .B(n364), .Z(n367) );
  XNOR2_X1 U424 ( .A(G99GAT), .B(G106GAT), .ZN(n366) );
  XNOR2_X1 U425 ( .A(n367), .B(n366), .ZN(n372) );
  XOR2_X1 U426 ( .A(n368), .B(G43GAT), .Z(n370) );
  NAND2_X1 U427 ( .A1(G232GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U428 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U429 ( .A(n372), .B(n371), .Z(n376) );
  INV_X1 U430 ( .A(n373), .ZN(n374) );
  XOR2_X1 U431 ( .A(n374), .B(G29GAT), .Z(n375) );
  XNOR2_X1 U432 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U433 ( .A(n378), .B(n377), .ZN(n565) );
  INV_X1 U434 ( .A(n565), .ZN(n549) );
  NAND2_X1 U435 ( .A1(n379), .A2(n549), .ZN(n380) );
  XNOR2_X1 U436 ( .A(n380), .B(KEYINPUT47), .ZN(n385) );
  XOR2_X1 U437 ( .A(n565), .B(KEYINPUT36), .Z(n481) );
  NOR2_X1 U438 ( .A1(n481), .A2(n578), .ZN(n381) );
  XNOR2_X1 U439 ( .A(n381), .B(KEYINPUT45), .ZN(n382) );
  NAND2_X1 U440 ( .A1(n382), .A2(n574), .ZN(n383) );
  XNOR2_X1 U441 ( .A(KEYINPUT67), .B(n569), .ZN(n557) );
  NOR2_X1 U442 ( .A1(n383), .A2(n557), .ZN(n384) );
  NOR2_X1 U443 ( .A1(n385), .A2(n384), .ZN(n386) );
  XNOR2_X1 U444 ( .A(KEYINPUT48), .B(n386), .ZN(n522) );
  NOR2_X1 U445 ( .A1(n515), .A2(n522), .ZN(n387) );
  XNOR2_X1 U446 ( .A(n387), .B(KEYINPUT54), .ZN(n407) );
  XOR2_X1 U447 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n389) );
  XNOR2_X1 U448 ( .A(G141GAT), .B(KEYINPUT5), .ZN(n388) );
  XNOR2_X1 U449 ( .A(n389), .B(n388), .ZN(n395) );
  XOR2_X1 U450 ( .A(G85GAT), .B(n390), .Z(n393) );
  XNOR2_X1 U451 ( .A(n391), .B(G113GAT), .ZN(n392) );
  XNOR2_X1 U452 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U453 ( .A(n395), .B(n394), .Z(n397) );
  NAND2_X1 U454 ( .A1(G225GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U455 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U456 ( .A(n398), .B(KEYINPUT4), .Z(n402) );
  XOR2_X1 U457 ( .A(G155GAT), .B(KEYINPUT2), .Z(n400) );
  XNOR2_X1 U458 ( .A(G162GAT), .B(KEYINPUT3), .ZN(n399) );
  XNOR2_X1 U459 ( .A(n400), .B(n399), .ZN(n413) );
  XNOR2_X1 U460 ( .A(n413), .B(KEYINPUT93), .ZN(n401) );
  XNOR2_X1 U461 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U462 ( .A(KEYINPUT0), .B(G134GAT), .Z(n404) );
  XNOR2_X1 U463 ( .A(G127GAT), .B(G120GAT), .ZN(n403) );
  XNOR2_X1 U464 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U465 ( .A(KEYINPUT78), .B(n405), .ZN(n443) );
  XNOR2_X1 U466 ( .A(n406), .B(n443), .ZN(n457) );
  XNOR2_X1 U467 ( .A(KEYINPUT94), .B(n457), .ZN(n536) );
  NAND2_X1 U468 ( .A1(n407), .A2(n536), .ZN(n552) );
  XOR2_X1 U469 ( .A(KEYINPUT24), .B(KEYINPUT92), .Z(n411) );
  XNOR2_X1 U470 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U471 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U472 ( .A(n412), .B(KEYINPUT70), .Z(n418) );
  XOR2_X1 U473 ( .A(n413), .B(KEYINPUT22), .Z(n415) );
  NAND2_X1 U474 ( .A1(G228GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U476 ( .A(G50GAT), .B(n416), .ZN(n417) );
  XNOR2_X1 U477 ( .A(n418), .B(n417), .ZN(n424) );
  XOR2_X1 U478 ( .A(KEYINPUT89), .B(KEYINPUT88), .Z(n420) );
  XNOR2_X1 U479 ( .A(G148GAT), .B(KEYINPUT23), .ZN(n419) );
  XNOR2_X1 U480 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U481 ( .A(n422), .B(n421), .Z(n423) );
  XNOR2_X1 U482 ( .A(n424), .B(n423), .ZN(n553) );
  XOR2_X1 U483 ( .A(KEYINPUT82), .B(KEYINPUT80), .Z(n426) );
  XNOR2_X1 U484 ( .A(KEYINPUT84), .B(KEYINPUT83), .ZN(n425) );
  XNOR2_X1 U485 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U486 ( .A(KEYINPUT20), .B(KEYINPUT79), .Z(n428) );
  XNOR2_X1 U487 ( .A(KEYINPUT81), .B(KEYINPUT85), .ZN(n427) );
  XNOR2_X1 U488 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U489 ( .A(n430), .B(n429), .Z(n441) );
  XOR2_X1 U490 ( .A(n431), .B(G176GAT), .Z(n433) );
  NAND2_X1 U491 ( .A1(G227GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U492 ( .A(n433), .B(n432), .ZN(n439) );
  XOR2_X1 U493 ( .A(KEYINPUT86), .B(n434), .Z(n437) );
  XNOR2_X1 U494 ( .A(G190GAT), .B(n435), .ZN(n436) );
  XNOR2_X1 U495 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U496 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U497 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X2 U498 ( .A(n443), .B(n442), .Z(n555) );
  NAND2_X1 U499 ( .A1(n553), .A2(n555), .ZN(n444) );
  XNOR2_X1 U500 ( .A(n444), .B(KEYINPUT26), .ZN(n454) );
  XOR2_X1 U501 ( .A(KEYINPUT122), .B(n445), .Z(n579) );
  NOR2_X1 U502 ( .A1(n579), .A2(n481), .ZN(n448) );
  NAND2_X1 U503 ( .A1(n557), .A2(n574), .ZN(n487) );
  NOR2_X1 U504 ( .A1(n555), .A2(n515), .ZN(n449) );
  XOR2_X1 U505 ( .A(n450), .B(KEYINPUT98), .Z(n451) );
  XNOR2_X1 U506 ( .A(KEYINPUT25), .B(n451), .ZN(n455) );
  XNOR2_X1 U507 ( .A(KEYINPUT27), .B(KEYINPUT96), .ZN(n452) );
  XOR2_X1 U508 ( .A(n452), .B(n515), .Z(n461) );
  INV_X1 U509 ( .A(n461), .ZN(n453) );
  NOR2_X1 U510 ( .A1(n454), .A2(n453), .ZN(n538) );
  NOR2_X1 U511 ( .A1(n455), .A2(n538), .ZN(n456) );
  XNOR2_X1 U512 ( .A(n456), .B(KEYINPUT99), .ZN(n458) );
  NAND2_X1 U513 ( .A1(n458), .A2(n457), .ZN(n465) );
  XOR2_X1 U514 ( .A(KEYINPUT28), .B(n553), .Z(n519) );
  INV_X1 U515 ( .A(n519), .ZN(n459) );
  NOR2_X1 U516 ( .A1(n459), .A2(n536), .ZN(n460) );
  NAND2_X1 U517 ( .A1(n461), .A2(n460), .ZN(n523) );
  XNOR2_X1 U518 ( .A(KEYINPUT97), .B(n523), .ZN(n463) );
  XOR2_X1 U519 ( .A(KEYINPUT87), .B(n555), .Z(n462) );
  NAND2_X1 U520 ( .A1(n463), .A2(n462), .ZN(n464) );
  NAND2_X1 U521 ( .A1(n465), .A2(n464), .ZN(n466) );
  XNOR2_X1 U522 ( .A(KEYINPUT100), .B(n466), .ZN(n483) );
  NOR2_X1 U523 ( .A1(n565), .A2(n578), .ZN(n469) );
  XOR2_X1 U524 ( .A(KEYINPUT76), .B(KEYINPUT16), .Z(n467) );
  XNOR2_X1 U525 ( .A(KEYINPUT77), .B(n467), .ZN(n468) );
  XNOR2_X1 U526 ( .A(n469), .B(n468), .ZN(n470) );
  NAND2_X1 U527 ( .A1(n483), .A2(n470), .ZN(n498) );
  NOR2_X1 U528 ( .A1(n487), .A2(n498), .ZN(n471) );
  XNOR2_X1 U529 ( .A(KEYINPUT101), .B(n471), .ZN(n479) );
  NOR2_X1 U530 ( .A1(n536), .A2(n479), .ZN(n473) );
  XNOR2_X1 U531 ( .A(KEYINPUT102), .B(KEYINPUT34), .ZN(n472) );
  XNOR2_X1 U532 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U533 ( .A(G1GAT), .B(n474), .Z(G1324GAT) );
  NOR2_X1 U534 ( .A1(n515), .A2(n479), .ZN(n476) );
  XNOR2_X1 U535 ( .A(G8GAT), .B(KEYINPUT103), .ZN(n475) );
  XNOR2_X1 U536 ( .A(n476), .B(n475), .ZN(G1325GAT) );
  NOR2_X1 U537 ( .A1(n555), .A2(n479), .ZN(n478) );
  XNOR2_X1 U538 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n478), .B(n477), .ZN(G1326GAT) );
  NOR2_X1 U540 ( .A1(n519), .A2(n479), .ZN(n480) );
  XOR2_X1 U541 ( .A(G22GAT), .B(n480), .Z(G1327GAT) );
  XNOR2_X1 U542 ( .A(KEYINPUT106), .B(KEYINPUT37), .ZN(n486) );
  INV_X1 U543 ( .A(n578), .ZN(n563) );
  NOR2_X1 U544 ( .A1(n481), .A2(n563), .ZN(n482) );
  NAND2_X1 U545 ( .A1(n483), .A2(n482), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(n513) );
  XNOR2_X1 U547 ( .A(KEYINPUT107), .B(KEYINPUT38), .ZN(n488) );
  NOR2_X1 U548 ( .A1(n496), .A2(n536), .ZN(n491) );
  XNOR2_X1 U549 ( .A(KEYINPUT104), .B(KEYINPUT39), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U551 ( .A(G29GAT), .B(n492), .ZN(G1328GAT) );
  NOR2_X1 U552 ( .A1(n496), .A2(n515), .ZN(n493) );
  XOR2_X1 U553 ( .A(G36GAT), .B(n493), .Z(G1329GAT) );
  NOR2_X1 U554 ( .A1(n496), .A2(n555), .ZN(n494) );
  XOR2_X1 U555 ( .A(KEYINPUT40), .B(n494), .Z(n495) );
  XNOR2_X1 U556 ( .A(n495), .B(G43GAT), .ZN(G1330GAT) );
  NOR2_X1 U557 ( .A1(n496), .A2(n519), .ZN(n497) );
  XOR2_X1 U558 ( .A(G50GAT), .B(n497), .Z(G1331GAT) );
  INV_X1 U559 ( .A(n541), .ZN(n559) );
  NAND2_X1 U560 ( .A1(n559), .A2(n569), .ZN(n512) );
  NOR2_X1 U561 ( .A1(n512), .A2(n498), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n499), .B(KEYINPUT109), .ZN(n508) );
  NOR2_X1 U563 ( .A1(n508), .A2(n536), .ZN(n503) );
  XOR2_X1 U564 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n501) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(KEYINPUT110), .ZN(n500) );
  XNOR2_X1 U566 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n503), .B(n502), .ZN(G1332GAT) );
  NOR2_X1 U568 ( .A1(n515), .A2(n508), .ZN(n505) );
  XNOR2_X1 U569 ( .A(G64GAT), .B(KEYINPUT111), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n505), .B(n504), .ZN(G1333GAT) );
  NOR2_X1 U571 ( .A1(n555), .A2(n508), .ZN(n506) );
  XOR2_X1 U572 ( .A(KEYINPUT112), .B(n506), .Z(n507) );
  XNOR2_X1 U573 ( .A(G71GAT), .B(n507), .ZN(G1334GAT) );
  NOR2_X1 U574 ( .A1(n519), .A2(n508), .ZN(n510) );
  XNOR2_X1 U575 ( .A(KEYINPUT43), .B(KEYINPUT113), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U577 ( .A(G78GAT), .B(n511), .Z(G1335GAT) );
  OR2_X1 U578 ( .A1(n513), .A2(n512), .ZN(n518) );
  NOR2_X1 U579 ( .A1(n536), .A2(n518), .ZN(n514) );
  XOR2_X1 U580 ( .A(G85GAT), .B(n514), .Z(G1336GAT) );
  NOR2_X1 U581 ( .A1(n515), .A2(n518), .ZN(n516) );
  XOR2_X1 U582 ( .A(G92GAT), .B(n516), .Z(G1337GAT) );
  NOR2_X1 U583 ( .A1(n555), .A2(n518), .ZN(n517) );
  XOR2_X1 U584 ( .A(G99GAT), .B(n517), .Z(G1338GAT) );
  NOR2_X1 U585 ( .A1(n519), .A2(n518), .ZN(n520) );
  XOR2_X1 U586 ( .A(KEYINPUT44), .B(n520), .Z(n521) );
  XNOR2_X1 U587 ( .A(G106GAT), .B(n521), .ZN(G1339GAT) );
  XOR2_X1 U588 ( .A(G113GAT), .B(KEYINPUT115), .Z(n526) );
  OR2_X1 U589 ( .A1(n555), .A2(n523), .ZN(n524) );
  NOR2_X1 U590 ( .A1(n522), .A2(n524), .ZN(n532) );
  NAND2_X1 U591 ( .A1(n532), .A2(n557), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n526), .B(n525), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(G120GAT), .B(KEYINPUT49), .Z(n528) );
  NAND2_X1 U594 ( .A1(n532), .A2(n559), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(G1341GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n530) );
  NAND2_X1 U597 ( .A1(n532), .A2(n563), .ZN(n529) );
  XNOR2_X1 U598 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U599 ( .A(G127GAT), .B(n531), .Z(G1342GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT51), .B(KEYINPUT117), .Z(n534) );
  NAND2_X1 U601 ( .A1(n532), .A2(n565), .ZN(n533) );
  XNOR2_X1 U602 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U603 ( .A(G134GAT), .B(n535), .Z(G1343GAT) );
  NOR2_X1 U604 ( .A1(n536), .A2(n522), .ZN(n537) );
  NAND2_X1 U605 ( .A1(n538), .A2(n537), .ZN(n548) );
  NOR2_X1 U606 ( .A1(n569), .A2(n548), .ZN(n539) );
  XOR2_X1 U607 ( .A(KEYINPUT118), .B(n539), .Z(n540) );
  XNOR2_X1 U608 ( .A(G141GAT), .B(n540), .ZN(G1344GAT) );
  NOR2_X1 U609 ( .A1(n548), .A2(n541), .ZN(n545) );
  XOR2_X1 U610 ( .A(KEYINPUT119), .B(KEYINPUT52), .Z(n543) );
  XNOR2_X1 U611 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n542) );
  XNOR2_X1 U612 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(G1345GAT) );
  NOR2_X1 U614 ( .A1(n578), .A2(n548), .ZN(n546) );
  XOR2_X1 U615 ( .A(KEYINPUT120), .B(n546), .Z(n547) );
  XNOR2_X1 U616 ( .A(G155GAT), .B(n547), .ZN(G1346GAT) );
  NOR2_X1 U617 ( .A1(n549), .A2(n548), .ZN(n551) );
  XNOR2_X1 U618 ( .A(G162GAT), .B(KEYINPUT121), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(G1347GAT) );
  NOR2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(KEYINPUT55), .ZN(n556) );
  NOR2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n566) );
  NAND2_X1 U623 ( .A1(n566), .A2(n557), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n561) );
  NAND2_X1 U626 ( .A1(n566), .A2(n559), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(G176GAT), .B(n562), .ZN(G1349GAT) );
  NAND2_X1 U629 ( .A1(n566), .A2(n563), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U631 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n568) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(G1351GAT) );
  NOR2_X1 U634 ( .A1(n569), .A2(n579), .ZN(n573) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  NOR2_X1 U639 ( .A1(n579), .A2(n574), .ZN(n576) );
  XNOR2_X1 U640 ( .A(KEYINPUT124), .B(KEYINPUT61), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G204GAT), .B(n577), .ZN(G1353GAT) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U644 ( .A(KEYINPUT125), .B(KEYINPUT126), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G211GAT), .B(n582), .ZN(G1354GAT) );
endmodule

