

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590;

  NOR2_X4 U323 ( .A1(n533), .A2(n291), .ZN(n570) );
  XNOR2_X1 U324 ( .A(n479), .B(KEYINPUT65), .ZN(n573) );
  XNOR2_X1 U325 ( .A(n476), .B(KEYINPUT48), .ZN(n546) );
  XNOR2_X1 U326 ( .A(n422), .B(n421), .ZN(n560) );
  XOR2_X1 U327 ( .A(KEYINPUT55), .B(n481), .Z(n291) );
  XNOR2_X1 U328 ( .A(KEYINPUT45), .B(KEYINPUT118), .ZN(n292) );
  NOR2_X1 U329 ( .A1(n576), .A2(n467), .ZN(n468) );
  OR2_X1 U330 ( .A1(n373), .A2(n523), .ZN(n352) );
  INV_X1 U331 ( .A(KEYINPUT98), .ZN(n329) );
  XNOR2_X1 U332 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U333 ( .A(n352), .B(KEYINPUT100), .ZN(n547) );
  XNOR2_X1 U334 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U335 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U336 ( .A(n332), .B(n331), .ZN(n333) );
  NAND2_X1 U337 ( .A1(n570), .A2(n538), .ZN(n564) );
  INV_X1 U338 ( .A(G99GAT), .ZN(n461) );
  XNOR2_X1 U339 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U340 ( .A(n461), .B(KEYINPUT116), .ZN(n462) );
  XNOR2_X1 U341 ( .A(n483), .B(n482), .ZN(G1348GAT) );
  XNOR2_X1 U342 ( .A(n463), .B(n462), .ZN(G1338GAT) );
  XOR2_X1 U343 ( .A(KEYINPUT0), .B(G127GAT), .Z(n340) );
  XOR2_X1 U344 ( .A(G190GAT), .B(G134GAT), .Z(n294) );
  XNOR2_X1 U345 ( .A(G43GAT), .B(G99GAT), .ZN(n293) );
  XNOR2_X1 U346 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U347 ( .A(n340), .B(n295), .Z(n297) );
  NAND2_X1 U348 ( .A1(G227GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U349 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U350 ( .A(KEYINPUT83), .B(KEYINPUT20), .Z(n299) );
  XNOR2_X1 U351 ( .A(G113GAT), .B(KEYINPUT86), .ZN(n298) );
  XNOR2_X1 U352 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U353 ( .A(n301), .B(n300), .Z(n311) );
  XOR2_X1 U354 ( .A(KEYINPUT18), .B(KEYINPUT84), .Z(n303) );
  XNOR2_X1 U355 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U357 ( .A(n304), .B(KEYINPUT85), .Z(n306) );
  XNOR2_X1 U358 ( .A(G169GAT), .B(G183GAT), .ZN(n305) );
  XNOR2_X1 U359 ( .A(n306), .B(n305), .ZN(n334) );
  XOR2_X1 U360 ( .A(G120GAT), .B(G176GAT), .Z(n308) );
  XNOR2_X1 U361 ( .A(G15GAT), .B(G71GAT), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U363 ( .A(n334), .B(n309), .ZN(n310) );
  XNOR2_X1 U364 ( .A(n311), .B(n310), .ZN(n533) );
  INV_X1 U365 ( .A(KEYINPUT103), .ZN(n384) );
  XOR2_X1 U366 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n313) );
  XNOR2_X1 U367 ( .A(G218GAT), .B(KEYINPUT88), .ZN(n312) );
  XNOR2_X1 U368 ( .A(n313), .B(n312), .ZN(n315) );
  INV_X1 U369 ( .A(KEYINPUT21), .ZN(n314) );
  XNOR2_X1 U370 ( .A(n315), .B(n314), .ZN(n317) );
  XNOR2_X1 U371 ( .A(G197GAT), .B(G211GAT), .ZN(n316) );
  XNOR2_X1 U372 ( .A(n317), .B(n316), .ZN(n322) );
  INV_X1 U373 ( .A(n322), .ZN(n365) );
  XOR2_X1 U374 ( .A(KEYINPUT97), .B(G92GAT), .Z(n319) );
  XOR2_X1 U375 ( .A(G36GAT), .B(G190GAT), .Z(n404) );
  XOR2_X1 U376 ( .A(G8GAT), .B(KEYINPUT80), .Z(n391) );
  XNOR2_X1 U377 ( .A(n404), .B(n391), .ZN(n318) );
  XOR2_X1 U378 ( .A(n319), .B(n318), .Z(n321) );
  INV_X1 U379 ( .A(n321), .ZN(n320) );
  NAND2_X1 U380 ( .A1(n365), .A2(n320), .ZN(n324) );
  NAND2_X1 U381 ( .A1(n322), .A2(n321), .ZN(n323) );
  NAND2_X1 U382 ( .A1(n324), .A2(n323), .ZN(n326) );
  NAND2_X1 U383 ( .A1(G226GAT), .A2(G233GAT), .ZN(n325) );
  XNOR2_X1 U384 ( .A(n326), .B(n325), .ZN(n332) );
  XOR2_X1 U385 ( .A(G64GAT), .B(KEYINPUT76), .Z(n328) );
  XNOR2_X1 U386 ( .A(G176GAT), .B(G204GAT), .ZN(n327) );
  XNOR2_X1 U387 ( .A(n328), .B(n327), .ZN(n435) );
  XNOR2_X1 U388 ( .A(KEYINPUT99), .B(n435), .ZN(n330) );
  XOR2_X1 U389 ( .A(n334), .B(n333), .Z(n527) );
  XNOR2_X1 U390 ( .A(n527), .B(KEYINPUT27), .ZN(n373) );
  XOR2_X1 U391 ( .A(KEYINPUT3), .B(G162GAT), .Z(n336) );
  XNOR2_X1 U392 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n335) );
  XNOR2_X1 U393 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U394 ( .A(G141GAT), .B(n337), .ZN(n363) );
  XOR2_X1 U395 ( .A(KEYINPUT6), .B(KEYINPUT94), .Z(n339) );
  XNOR2_X1 U396 ( .A(KEYINPUT95), .B(KEYINPUT5), .ZN(n338) );
  XNOR2_X1 U397 ( .A(n339), .B(n338), .ZN(n350) );
  XOR2_X1 U398 ( .A(G120GAT), .B(G57GAT), .Z(n430) );
  XOR2_X1 U399 ( .A(G85GAT), .B(n430), .Z(n342) );
  XNOR2_X1 U400 ( .A(n340), .B(G148GAT), .ZN(n341) );
  XNOR2_X1 U401 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U402 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n344) );
  NAND2_X1 U403 ( .A1(G225GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U404 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U405 ( .A(n346), .B(n345), .Z(n348) );
  XOR2_X1 U406 ( .A(G113GAT), .B(G1GAT), .Z(n452) );
  XOR2_X1 U407 ( .A(G29GAT), .B(G134GAT), .Z(n410) );
  XNOR2_X1 U408 ( .A(n452), .B(n410), .ZN(n347) );
  XNOR2_X1 U409 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U410 ( .A(n350), .B(n349), .Z(n351) );
  XNOR2_X1 U411 ( .A(n363), .B(n351), .ZN(n379) );
  XNOR2_X1 U412 ( .A(KEYINPUT96), .B(n379), .ZN(n523) );
  XOR2_X1 U413 ( .A(KEYINPUT93), .B(KEYINPUT91), .Z(n354) );
  XNOR2_X1 U414 ( .A(KEYINPUT87), .B(KEYINPUT22), .ZN(n353) );
  XNOR2_X1 U415 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U416 ( .A(KEYINPUT92), .B(KEYINPUT24), .Z(n356) );
  XNOR2_X1 U417 ( .A(G204GAT), .B(KEYINPUT23), .ZN(n355) );
  XNOR2_X1 U418 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U419 ( .A(n358), .B(n357), .ZN(n369) );
  XOR2_X1 U420 ( .A(G78GAT), .B(G148GAT), .Z(n360) );
  XNOR2_X1 U421 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n359) );
  XNOR2_X1 U422 ( .A(n360), .B(n359), .ZN(n436) );
  XOR2_X1 U423 ( .A(G22GAT), .B(n436), .Z(n362) );
  NAND2_X1 U424 ( .A1(G228GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U425 ( .A(n362), .B(n361), .ZN(n364) );
  XNOR2_X1 U426 ( .A(n364), .B(n363), .ZN(n367) );
  XNOR2_X1 U427 ( .A(G50GAT), .B(n322), .ZN(n366) );
  XNOR2_X1 U428 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U429 ( .A(n369), .B(n368), .ZN(n480) );
  XOR2_X1 U430 ( .A(n480), .B(KEYINPUT28), .Z(n495) );
  NOR2_X1 U431 ( .A1(n547), .A2(n495), .ZN(n535) );
  NAND2_X1 U432 ( .A1(n535), .A2(n533), .ZN(n382) );
  INV_X1 U433 ( .A(n533), .ZN(n370) );
  NOR2_X1 U434 ( .A1(n480), .A2(n370), .ZN(n372) );
  XNOR2_X1 U435 ( .A(KEYINPUT101), .B(KEYINPUT26), .ZN(n371) );
  XNOR2_X1 U436 ( .A(n372), .B(n371), .ZN(n575) );
  OR2_X1 U437 ( .A1(n575), .A2(n373), .ZN(n378) );
  OR2_X1 U438 ( .A1(n533), .A2(n527), .ZN(n374) );
  NAND2_X1 U439 ( .A1(n374), .A2(n480), .ZN(n375) );
  XNOR2_X1 U440 ( .A(n375), .B(KEYINPUT25), .ZN(n376) );
  XOR2_X1 U441 ( .A(KEYINPUT102), .B(n376), .Z(n377) );
  NAND2_X1 U442 ( .A1(n378), .A2(n377), .ZN(n380) );
  NAND2_X1 U443 ( .A1(n380), .A2(n379), .ZN(n381) );
  NAND2_X1 U444 ( .A1(n382), .A2(n381), .ZN(n383) );
  XNOR2_X1 U445 ( .A(n384), .B(n383), .ZN(n487) );
  XOR2_X1 U446 ( .A(G78GAT), .B(G127GAT), .Z(n386) );
  XNOR2_X1 U447 ( .A(G1GAT), .B(G183GAT), .ZN(n385) );
  XNOR2_X1 U448 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U449 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n388) );
  XNOR2_X1 U450 ( .A(G57GAT), .B(G64GAT), .ZN(n387) );
  XNOR2_X1 U451 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U452 ( .A(n390), .B(n389), .ZN(n401) );
  XOR2_X1 U453 ( .A(G71GAT), .B(KEYINPUT13), .Z(n429) );
  XNOR2_X1 U454 ( .A(n429), .B(n391), .ZN(n393) );
  XOR2_X1 U455 ( .A(G211GAT), .B(G155GAT), .Z(n392) );
  XNOR2_X1 U456 ( .A(n393), .B(n392), .ZN(n399) );
  XOR2_X1 U457 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n395) );
  NAND2_X1 U458 ( .A1(G231GAT), .A2(G233GAT), .ZN(n394) );
  XOR2_X1 U459 ( .A(n395), .B(n394), .Z(n397) );
  XOR2_X1 U460 ( .A(G22GAT), .B(G15GAT), .Z(n448) );
  XNOR2_X1 U461 ( .A(n448), .B(KEYINPUT12), .ZN(n396) );
  XNOR2_X1 U462 ( .A(n401), .B(n400), .ZN(n584) );
  XOR2_X1 U463 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n403) );
  XNOR2_X1 U464 ( .A(G106GAT), .B(KEYINPUT10), .ZN(n402) );
  XNOR2_X1 U465 ( .A(n403), .B(n402), .ZN(n405) );
  XOR2_X1 U466 ( .A(n405), .B(n404), .Z(n407) );
  XNOR2_X1 U467 ( .A(G218GAT), .B(G162GAT), .ZN(n406) );
  XOR2_X1 U468 ( .A(n407), .B(n406), .Z(n414) );
  XOR2_X1 U469 ( .A(KEYINPUT75), .B(G92GAT), .Z(n409) );
  XNOR2_X1 U470 ( .A(G99GAT), .B(G85GAT), .ZN(n408) );
  XNOR2_X1 U471 ( .A(n409), .B(n408), .ZN(n434) );
  XOR2_X1 U472 ( .A(n434), .B(n410), .Z(n412) );
  NAND2_X1 U473 ( .A1(G232GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U474 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U475 ( .A(n414), .B(n413), .ZN(n422) );
  XOR2_X1 U476 ( .A(KEYINPUT7), .B(KEYINPUT72), .Z(n416) );
  XNOR2_X1 U477 ( .A(G50GAT), .B(G43GAT), .ZN(n415) );
  XNOR2_X1 U478 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U479 ( .A(KEYINPUT8), .B(n417), .ZN(n457) );
  XOR2_X1 U480 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n419) );
  XNOR2_X1 U481 ( .A(KEYINPUT67), .B(KEYINPUT66), .ZN(n418) );
  XNOR2_X1 U482 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U483 ( .A(n457), .B(n420), .Z(n421) );
  XNOR2_X1 U484 ( .A(n560), .B(KEYINPUT36), .ZN(n588) );
  NOR2_X1 U485 ( .A1(n584), .A2(n588), .ZN(n423) );
  NAND2_X1 U486 ( .A1(n487), .A2(n423), .ZN(n424) );
  XOR2_X1 U487 ( .A(KEYINPUT37), .B(n424), .Z(n500) );
  XOR2_X1 U488 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n426) );
  NAND2_X1 U489 ( .A1(G230GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U490 ( .A(n426), .B(n425), .ZN(n428) );
  INV_X1 U491 ( .A(KEYINPUT31), .ZN(n427) );
  XNOR2_X1 U492 ( .A(n428), .B(n427), .ZN(n432) );
  XNOR2_X1 U493 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U494 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U495 ( .A(n434), .B(n433), .Z(n438) );
  XNOR2_X1 U496 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U497 ( .A(n438), .B(n437), .ZN(n581) );
  XNOR2_X1 U498 ( .A(n581), .B(KEYINPUT64), .ZN(n439) );
  XNOR2_X1 U499 ( .A(n439), .B(KEYINPUT41), .ZN(n538) );
  XOR2_X1 U500 ( .A(KEYINPUT71), .B(KEYINPUT73), .Z(n441) );
  XNOR2_X1 U501 ( .A(KEYINPUT69), .B(KEYINPUT70), .ZN(n440) );
  XNOR2_X1 U502 ( .A(n441), .B(n440), .ZN(n456) );
  XOR2_X1 U503 ( .A(G141GAT), .B(G197GAT), .Z(n443) );
  XNOR2_X1 U504 ( .A(G29GAT), .B(G36GAT), .ZN(n442) );
  XNOR2_X1 U505 ( .A(n443), .B(n442), .ZN(n447) );
  XOR2_X1 U506 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n445) );
  XNOR2_X1 U507 ( .A(G169GAT), .B(G8GAT), .ZN(n444) );
  XNOR2_X1 U508 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U509 ( .A(n447), .B(n446), .Z(n454) );
  XOR2_X1 U510 ( .A(n448), .B(KEYINPUT29), .Z(n450) );
  NAND2_X1 U511 ( .A1(G229GAT), .A2(G233GAT), .ZN(n449) );
  XNOR2_X1 U512 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U513 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U514 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U515 ( .A(n456), .B(n455), .ZN(n458) );
  XNOR2_X1 U516 ( .A(n458), .B(n457), .ZN(n576) );
  INV_X1 U517 ( .A(n576), .ZN(n550) );
  NAND2_X1 U518 ( .A1(n538), .A2(n550), .ZN(n459) );
  XNOR2_X1 U519 ( .A(n459), .B(KEYINPUT110), .ZN(n513) );
  NOR2_X1 U520 ( .A1(n500), .A2(n513), .ZN(n460) );
  XNOR2_X1 U521 ( .A(n460), .B(KEYINPUT113), .ZN(n529) );
  NOR2_X1 U522 ( .A1(n533), .A2(n529), .ZN(n463) );
  INV_X1 U523 ( .A(n584), .ZN(n556) );
  NOR2_X1 U524 ( .A1(n588), .A2(n556), .ZN(n464) );
  XNOR2_X1 U525 ( .A(n464), .B(n292), .ZN(n465) );
  NAND2_X1 U526 ( .A1(n465), .A2(n581), .ZN(n466) );
  XOR2_X1 U527 ( .A(KEYINPUT119), .B(n466), .Z(n467) );
  XNOR2_X1 U528 ( .A(n468), .B(KEYINPUT120), .ZN(n475) );
  XOR2_X1 U529 ( .A(KEYINPUT46), .B(KEYINPUT117), .Z(n470) );
  NAND2_X1 U530 ( .A1(n538), .A2(n576), .ZN(n469) );
  XNOR2_X1 U531 ( .A(n470), .B(n469), .ZN(n471) );
  NAND2_X1 U532 ( .A1(n560), .A2(n471), .ZN(n472) );
  NOR2_X1 U533 ( .A1(n584), .A2(n472), .ZN(n473) );
  XOR2_X1 U534 ( .A(KEYINPUT47), .B(n473), .Z(n474) );
  NOR2_X1 U535 ( .A1(n475), .A2(n474), .ZN(n476) );
  NOR2_X1 U536 ( .A1(n527), .A2(n546), .ZN(n477) );
  XNOR2_X1 U537 ( .A(n477), .B(KEYINPUT54), .ZN(n478) );
  NAND2_X1 U538 ( .A1(n478), .A2(n523), .ZN(n479) );
  NAND2_X1 U539 ( .A1(n573), .A2(n480), .ZN(n481) );
  NAND2_X1 U540 ( .A1(n570), .A2(n576), .ZN(n483) );
  XNOR2_X1 U541 ( .A(G169GAT), .B(KEYINPUT124), .ZN(n482) );
  NAND2_X1 U542 ( .A1(n576), .A2(n581), .ZN(n484) );
  XOR2_X1 U543 ( .A(KEYINPUT77), .B(n484), .Z(n499) );
  INV_X1 U544 ( .A(n560), .ZN(n569) );
  NOR2_X1 U545 ( .A1(n556), .A2(n569), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n485), .B(KEYINPUT16), .ZN(n486) );
  NAND2_X1 U547 ( .A1(n487), .A2(n486), .ZN(n512) );
  OR2_X1 U548 ( .A1(n499), .A2(n512), .ZN(n496) );
  NOR2_X1 U549 ( .A1(n523), .A2(n496), .ZN(n489) );
  XNOR2_X1 U550 ( .A(KEYINPUT34), .B(KEYINPUT104), .ZN(n488) );
  XNOR2_X1 U551 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U552 ( .A(G1GAT), .B(n490), .Z(G1324GAT) );
  NOR2_X1 U553 ( .A1(n527), .A2(n496), .ZN(n491) );
  XOR2_X1 U554 ( .A(G8GAT), .B(n491), .Z(G1325GAT) );
  NOR2_X1 U555 ( .A1(n533), .A2(n496), .ZN(n493) );
  XNOR2_X1 U556 ( .A(KEYINPUT105), .B(KEYINPUT35), .ZN(n492) );
  XNOR2_X1 U557 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U558 ( .A(G15GAT), .B(n494), .Z(G1326GAT) );
  INV_X1 U559 ( .A(n495), .ZN(n530) );
  NOR2_X1 U560 ( .A1(n530), .A2(n496), .ZN(n497) );
  XOR2_X1 U561 ( .A(KEYINPUT106), .B(n497), .Z(n498) );
  XNOR2_X1 U562 ( .A(G22GAT), .B(n498), .ZN(G1327GAT) );
  NOR2_X1 U563 ( .A1(n500), .A2(n499), .ZN(n502) );
  XNOR2_X1 U564 ( .A(KEYINPUT38), .B(KEYINPUT107), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n502), .B(n501), .ZN(n510) );
  NOR2_X1 U566 ( .A1(n510), .A2(n523), .ZN(n504) );
  XNOR2_X1 U567 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n504), .B(n503), .ZN(G1328GAT) );
  NOR2_X1 U569 ( .A1(n527), .A2(n510), .ZN(n505) );
  XOR2_X1 U570 ( .A(KEYINPUT108), .B(n505), .Z(n506) );
  XNOR2_X1 U571 ( .A(G36GAT), .B(n506), .ZN(G1329GAT) );
  XNOR2_X1 U572 ( .A(KEYINPUT40), .B(KEYINPUT109), .ZN(n508) );
  NOR2_X1 U573 ( .A1(n533), .A2(n510), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U575 ( .A(G43GAT), .B(n509), .ZN(G1330GAT) );
  NOR2_X1 U576 ( .A1(n510), .A2(n530), .ZN(n511) );
  XOR2_X1 U577 ( .A(G50GAT), .B(n511), .Z(G1331GAT) );
  OR2_X1 U578 ( .A1(n513), .A2(n512), .ZN(n520) );
  NOR2_X1 U579 ( .A1(n523), .A2(n520), .ZN(n515) );
  XNOR2_X1 U580 ( .A(KEYINPUT42), .B(KEYINPUT111), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U582 ( .A(G57GAT), .B(n516), .ZN(G1332GAT) );
  NOR2_X1 U583 ( .A1(n527), .A2(n520), .ZN(n517) );
  XOR2_X1 U584 ( .A(KEYINPUT112), .B(n517), .Z(n518) );
  XNOR2_X1 U585 ( .A(G64GAT), .B(n518), .ZN(G1333GAT) );
  NOR2_X1 U586 ( .A1(n533), .A2(n520), .ZN(n519) );
  XOR2_X1 U587 ( .A(G71GAT), .B(n519), .Z(G1334GAT) );
  NOR2_X1 U588 ( .A1(n530), .A2(n520), .ZN(n522) );
  XNOR2_X1 U589 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n521) );
  XNOR2_X1 U590 ( .A(n522), .B(n521), .ZN(G1335GAT) );
  NOR2_X1 U591 ( .A1(n523), .A2(n529), .ZN(n525) );
  XNOR2_X1 U592 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n524) );
  XNOR2_X1 U593 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U594 ( .A(G85GAT), .B(n526), .ZN(G1336GAT) );
  NOR2_X1 U595 ( .A1(n527), .A2(n529), .ZN(n528) );
  XOR2_X1 U596 ( .A(G92GAT), .B(n528), .Z(G1337GAT) );
  NOR2_X1 U597 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U598 ( .A(KEYINPUT44), .B(n531), .Z(n532) );
  XNOR2_X1 U599 ( .A(G106GAT), .B(n532), .ZN(G1339GAT) );
  NOR2_X1 U600 ( .A1(n546), .A2(n533), .ZN(n534) );
  NAND2_X1 U601 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U602 ( .A(KEYINPUT121), .B(n536), .ZN(n543) );
  NAND2_X1 U603 ( .A1(n543), .A2(n576), .ZN(n537) );
  XNOR2_X1 U604 ( .A(G113GAT), .B(n537), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .Z(n540) );
  INV_X1 U606 ( .A(n538), .ZN(n552) );
  NAND2_X1 U607 ( .A1(n543), .A2(n538), .ZN(n539) );
  XNOR2_X1 U608 ( .A(n540), .B(n539), .ZN(G1341GAT) );
  NAND2_X1 U609 ( .A1(n543), .A2(n584), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n541), .B(KEYINPUT50), .ZN(n542) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n542), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U613 ( .A1(n543), .A2(n569), .ZN(n544) );
  XNOR2_X1 U614 ( .A(n545), .B(n544), .ZN(G1343GAT) );
  INV_X1 U615 ( .A(n546), .ZN(n549) );
  NOR2_X1 U616 ( .A1(n575), .A2(n547), .ZN(n548) );
  NAND2_X1 U617 ( .A1(n549), .A2(n548), .ZN(n559) );
  NOR2_X1 U618 ( .A1(n550), .A2(n559), .ZN(n551) );
  XOR2_X1 U619 ( .A(G141GAT), .B(n551), .Z(G1344GAT) );
  NOR2_X1 U620 ( .A1(n552), .A2(n559), .ZN(n554) );
  XNOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(n555), .ZN(G1345GAT) );
  NOR2_X1 U624 ( .A1(n556), .A2(n559), .ZN(n557) );
  XOR2_X1 U625 ( .A(KEYINPUT122), .B(n557), .Z(n558) );
  XNOR2_X1 U626 ( .A(G155GAT), .B(n558), .ZN(G1346GAT) );
  NOR2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n562) );
  XNOR2_X1 U628 ( .A(G162GAT), .B(KEYINPUT123), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(G1347GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n563) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(n565), .ZN(G1349GAT) );
  NAND2_X1 U632 ( .A1(n570), .A2(n584), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U634 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n567), .B(KEYINPUT125), .ZN(n568) );
  XOR2_X1 U636 ( .A(KEYINPUT126), .B(n568), .Z(n572) );
  NAND2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(G1351GAT) );
  XOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT60), .Z(n578) );
  INV_X1 U640 ( .A(n573), .ZN(n574) );
  NOR2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n585) );
  NAND2_X1 U642 ( .A1(n585), .A2(n576), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n580) );
  XOR2_X1 U644 ( .A(KEYINPUT127), .B(KEYINPUT59), .Z(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .Z(n583) );
  INV_X1 U647 ( .A(n585), .ZN(n587) );
  OR2_X1 U648 ( .A1(n587), .A2(n581), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U653 ( .A(KEYINPUT62), .B(n589), .Z(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

