//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 1 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n819, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n979, new_n980,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1021, new_n1022, new_n1023, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G22gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G211gat), .A2(G218gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT22), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G204gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G197gat), .ZN(new_n211));
  INV_X1    g010(.A(G197gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G204gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n209), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n207), .ZN(new_n215));
  NOR2_X1   g014(.A1(G211gat), .A2(G218gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(G211gat), .B(G218gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(G197gat), .B(G204gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(new_n220), .A3(new_n209), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT29), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT3), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G141gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n225), .A2(KEYINPUT76), .A3(G148gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT76), .ZN(new_n227));
  INV_X1    g026(.A(G148gat), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n227), .B1(G141gat), .B2(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(G141gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n226), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(G155gat), .A2(G162gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT2), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G155gat), .ZN(new_n235));
  INV_X1    g034(.A(G162gat), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n234), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n231), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n225), .A2(G148gat), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n233), .B1(new_n230), .B2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(G155gat), .B(G162gat), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT77), .ZN(new_n245));
  AOI22_X1  g044(.A1(new_n231), .A2(new_n237), .B1(new_n240), .B2(new_n242), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT77), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n224), .B1(new_n245), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT29), .B1(new_n246), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n251), .A2(new_n222), .ZN(new_n252));
  INV_X1    g051(.A(G228gat), .ZN(new_n253));
  INV_X1    g052(.A(G233gat), .ZN(new_n254));
  OAI22_X1  g053(.A1(new_n249), .A2(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n253), .A2(new_n254), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n214), .A2(new_n217), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n219), .B1(new_n209), .B2(new_n220), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n223), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(new_n250), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT82), .B1(new_n260), .B2(new_n244), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT29), .B1(new_n218), .B2(new_n221), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n244), .B(KEYINPUT82), .C1(new_n262), .C2(KEYINPUT3), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n256), .B1(new_n261), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT83), .B1(new_n251), .B2(new_n222), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT83), .ZN(new_n267));
  INV_X1    g066(.A(new_n222), .ZN(new_n268));
  AND2_X1   g067(.A1(G155gat), .A2(G162gat), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n269), .B1(new_n233), .B2(new_n232), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n225), .A2(G148gat), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n271), .B1(new_n239), .B2(new_n227), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n270), .B1(new_n226), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n228), .A2(G141gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n241), .B1(new_n233), .B2(new_n275), .ZN(new_n276));
  NOR3_X1   g075(.A1(new_n273), .A2(KEYINPUT3), .A3(new_n276), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n267), .B(new_n268), .C1(new_n277), .C2(KEYINPUT29), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n266), .A2(new_n278), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n206), .B(new_n255), .C1(new_n265), .C2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT84), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n255), .B1(new_n265), .B2(new_n279), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(G22gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n282), .A2(KEYINPUT84), .A3(G22gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT82), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n287), .B1(new_n224), .B2(new_n246), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(new_n263), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n289), .A2(new_n256), .A3(new_n266), .A4(new_n278), .ZN(new_n290));
  AND3_X1   g089(.A1(new_n290), .A2(new_n206), .A3(new_n255), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n206), .B1(new_n290), .B2(new_n255), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT81), .ZN(new_n293));
  OAI22_X1  g092(.A1(new_n291), .A2(new_n292), .B1(new_n293), .B2(new_n205), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n205), .B1(new_n286), .B2(new_n294), .ZN(new_n295));
  AOI211_X1 g094(.A(new_n293), .B(new_n204), .C1(new_n283), .C2(new_n280), .ZN(new_n296));
  OAI21_X1  g095(.A(KEYINPUT85), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n292), .B1(KEYINPUT84), .B2(new_n280), .ZN(new_n298));
  INV_X1    g097(.A(new_n285), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n294), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(new_n204), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT85), .ZN(new_n302));
  INV_X1    g101(.A(new_n296), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n297), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT34), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT68), .B(G190gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT27), .B(G183gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n309), .A2(KEYINPUT70), .A3(KEYINPUT28), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G183gat), .A2(G190gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT26), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n313), .B(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n312), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT28), .B1(new_n309), .B2(KEYINPUT70), .ZN(new_n319));
  NOR3_X1   g118(.A1(new_n311), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n313), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT23), .ZN(new_n323));
  OAI211_X1 g122(.A(KEYINPUT25), .B(new_n316), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT66), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n325), .B1(new_n313), .B2(KEYINPUT23), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n322), .A2(KEYINPUT66), .A3(new_n323), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n324), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT69), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT67), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT24), .B1(new_n312), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n312), .A2(new_n330), .A3(KEYINPUT24), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G190gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT68), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT68), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(G190gat), .ZN(new_n338));
  INV_X1    g137(.A(G183gat), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n336), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n329), .B1(new_n334), .B2(new_n340), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n312), .A2(new_n330), .A3(KEYINPUT24), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n340), .B(new_n329), .C1(new_n342), .C2(new_n331), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n328), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n327), .A2(new_n326), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT65), .B(G176gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n323), .A2(G169gat), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n317), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n312), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT64), .ZN(new_n352));
  INV_X1    g151(.A(new_n312), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n351), .A2(new_n352), .B1(KEYINPUT24), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT24), .ZN(new_n355));
  NOR3_X1   g154(.A1(new_n312), .A2(new_n355), .A3(KEYINPUT64), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n346), .B(new_n349), .C1(new_n354), .C2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT25), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n345), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(G120gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(G113gat), .ZN(new_n362));
  INV_X1    g161(.A(G113gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(G120gat), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT1), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(G127gat), .B(G134gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  OR2_X1    g167(.A1(KEYINPUT71), .A2(G134gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(KEYINPUT71), .A2(G134gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n369), .A2(G127gat), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(G127gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(G134gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n365), .B1(new_n374), .B2(KEYINPUT72), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT72), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n371), .A2(new_n376), .A3(new_n373), .ZN(new_n377));
  AOI211_X1 g176(.A(KEYINPUT73), .B(new_n368), .C1(new_n375), .C2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT73), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n374), .A2(KEYINPUT72), .ZN(new_n380));
  INV_X1    g179(.A(new_n365), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(new_n377), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n379), .B1(new_n382), .B2(new_n367), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n321), .B(new_n360), .C1(new_n378), .C2(new_n383), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n371), .A2(new_n376), .A3(new_n373), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n376), .B1(new_n371), .B2(new_n373), .ZN(new_n386));
  NOR3_X1   g185(.A1(new_n385), .A2(new_n386), .A3(new_n365), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT73), .B1(new_n387), .B2(new_n368), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n382), .A2(new_n379), .A3(new_n367), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n340), .B1(new_n342), .B2(new_n331), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT69), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(new_n343), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n392), .A2(new_n328), .B1(new_n357), .B2(new_n358), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n388), .B(new_n389), .C1(new_n393), .C2(new_n320), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n384), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(G227gat), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n396), .A2(new_n254), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n306), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  AOI211_X1 g198(.A(KEYINPUT34), .B(new_n397), .C1(new_n384), .C2(new_n394), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n394), .A3(new_n397), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT33), .ZN(new_n403));
  XOR2_X1   g202(.A(G15gat), .B(G43gat), .Z(new_n404));
  XNOR2_X1  g203(.A(G71gat), .B(G99gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n404), .B(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n402), .B(KEYINPUT32), .C1(new_n403), .C2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n402), .A2(new_n403), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n402), .A2(KEYINPUT32), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n410), .A3(new_n406), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n401), .A2(new_n408), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n399), .ZN(new_n413));
  INV_X1    g212(.A(new_n400), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n411), .A2(new_n408), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  XOR2_X1   g215(.A(G1gat), .B(G29gat), .Z(new_n417));
  XNOR2_X1  g216(.A(G57gat), .B(G85gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n420));
  XOR2_X1   g219(.A(new_n419), .B(new_n420), .Z(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT78), .ZN(new_n423));
  NAND2_X1  g222(.A1(G225gat), .A2(G233gat), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n244), .B1(new_n387), .B2(new_n368), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n382), .A2(new_n367), .A3(new_n246), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT5), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n423), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n424), .ZN(new_n430));
  NOR3_X1   g229(.A1(new_n387), .A2(new_n368), .A3(new_n244), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n246), .B1(new_n382), .B2(new_n367), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n433), .A2(KEYINPUT78), .A3(KEYINPUT5), .ZN(new_n434));
  NOR3_X1   g233(.A1(new_n273), .A2(KEYINPUT77), .A3(new_n276), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n247), .B1(new_n238), .B2(new_n243), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n388), .A2(new_n437), .A3(KEYINPUT4), .A4(new_n389), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n250), .B1(new_n238), .B2(new_n243), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n277), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n382), .A2(new_n367), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n430), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT4), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n438), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n429), .A2(new_n434), .A3(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n246), .B(new_n250), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n387), .A2(new_n368), .ZN(new_n448));
  OAI22_X1  g247(.A1(new_n447), .A2(new_n448), .B1(new_n426), .B2(new_n443), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n430), .A2(KEYINPUT5), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n388), .A2(new_n437), .A3(new_n389), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n450), .B(new_n451), .C1(KEYINPUT4), .C2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n422), .B1(new_n446), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n446), .A2(new_n453), .A3(new_n422), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT6), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n456), .A2(KEYINPUT80), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT80), .B1(new_n456), .B2(new_n457), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n455), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n454), .A2(KEYINPUT6), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n223), .B1(new_n393), .B2(new_n320), .ZN(new_n462));
  NAND2_X1  g261(.A1(G226gat), .A2(G233gat), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI211_X1 g263(.A(G226gat), .B(G233gat), .C1(new_n393), .C2(new_n320), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(new_n465), .A3(new_n222), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT75), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n464), .A2(KEYINPUT75), .A3(new_n465), .A4(new_n222), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n464), .A2(new_n465), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n268), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n468), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(G8gat), .B(G36gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(G64gat), .B(G92gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n473), .B(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n222), .B1(new_n464), .B2(new_n465), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n477), .B1(new_n467), .B2(new_n466), .ZN(new_n478));
  INV_X1    g277(.A(new_n475), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(new_n479), .A3(new_n469), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n476), .A2(new_n480), .A3(KEYINPUT30), .ZN(new_n481));
  OR3_X1    g280(.A1(new_n472), .A2(KEYINPUT30), .A3(new_n475), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n460), .A2(new_n461), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n305), .A2(new_n416), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT35), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n456), .A2(new_n457), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(new_n455), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n454), .A2(KEYINPUT88), .A3(KEYINPUT6), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT88), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n461), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n487), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n481), .A2(new_n482), .ZN(new_n492));
  XOR2_X1   g291(.A(KEYINPUT90), .B(KEYINPUT35), .Z(new_n493));
  AND2_X1   g292(.A1(new_n416), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n305), .A2(new_n491), .A3(new_n492), .A4(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT74), .B1(new_n412), .B2(new_n415), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT36), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g297(.A(KEYINPUT74), .B(KEYINPUT36), .C1(new_n412), .C2(new_n415), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n302), .B1(new_n301), .B2(new_n303), .ZN(new_n501));
  AOI211_X1 g300(.A(KEYINPUT85), .B(new_n296), .C1(new_n300), .C2(new_n204), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n460), .A2(new_n461), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n492), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n500), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n452), .A2(KEYINPUT4), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n430), .B1(new_n507), .B2(new_n449), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n431), .A2(new_n432), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n424), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n508), .A2(KEYINPUT39), .A3(new_n510), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n511), .B(new_n422), .C1(KEYINPUT39), .C2(new_n508), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT40), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n454), .B1(new_n512), .B2(new_n513), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n514), .A2(new_n515), .A3(new_n481), .A4(new_n482), .ZN(new_n516));
  XOR2_X1   g315(.A(KEYINPUT87), .B(KEYINPUT38), .Z(new_n517));
  NOR2_X1   g316(.A1(new_n472), .A2(KEYINPUT37), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n479), .B1(new_n472), .B2(KEYINPUT37), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n518), .B1(new_n519), .B2(KEYINPUT89), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT89), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT37), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n522), .B1(new_n478), .B2(new_n469), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n521), .B1(new_n523), .B2(new_n479), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n517), .B1(new_n520), .B2(new_n524), .ZN(new_n525));
  AOI22_X1  g324(.A1(new_n486), .A2(new_n455), .B1(new_n461), .B2(new_n489), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n466), .A2(KEYINPUT86), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT86), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n464), .A2(new_n528), .A3(new_n465), .A4(new_n222), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n527), .A2(new_n471), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT37), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n475), .A2(new_n517), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n531), .B(new_n532), .C1(KEYINPUT37), .C2(new_n472), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n526), .A2(new_n533), .A3(new_n488), .A4(new_n480), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n305), .B(new_n516), .C1(new_n525), .C2(new_n534), .ZN(new_n535));
  AOI22_X1  g334(.A1(new_n485), .A2(new_n495), .B1(new_n506), .B2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G113gat), .B(G141gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(KEYINPUT11), .ZN(new_n538));
  INV_X1    g337(.A(G169gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(G197gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT12), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n540), .B(new_n212), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT12), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT17), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT15), .ZN(new_n549));
  OR2_X1    g348(.A1(G43gat), .A2(G50gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(G43gat), .A2(G50gat), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G29gat), .A2(G36gat), .ZN(new_n554));
  OR3_X1    g353(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n550), .A2(new_n549), .A3(new_n551), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n553), .A2(new_n554), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n556), .A2(KEYINPUT91), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT91), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n561), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n560), .A2(new_n555), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT92), .ZN(new_n564));
  AOI22_X1  g363(.A1(new_n563), .A2(new_n564), .B1(G29gat), .B2(G36gat), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n560), .A2(new_n555), .A3(KEYINPUT92), .A4(new_n562), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n548), .B(new_n559), .C1(new_n567), .C2(new_n553), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n553), .B1(new_n565), .B2(new_n566), .ZN(new_n569));
  INV_X1    g368(.A(new_n559), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT17), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G15gat), .B(G22gat), .ZN(new_n573));
  INV_X1    g372(.A(G1gat), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n573), .A2(KEYINPUT16), .A3(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n575), .B1(new_n574), .B2(new_n573), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(G8gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n572), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G229gat), .A2(G233gat), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n569), .A2(new_n570), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n580), .A2(new_n577), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n578), .A2(KEYINPUT18), .A3(new_n579), .A4(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n579), .B(KEYINPUT13), .Z(new_n584));
  INV_X1    g383(.A(new_n580), .ZN(new_n585));
  INV_X1    g384(.A(new_n577), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n584), .B1(new_n587), .B2(new_n581), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n583), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n581), .B1(new_n572), .B2(new_n577), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT18), .B1(new_n590), .B2(new_n579), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n547), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n578), .A2(new_n579), .A3(new_n582), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT18), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n595), .A2(new_n583), .A3(new_n588), .A4(new_n546), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n592), .A2(KEYINPUT93), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(KEYINPUT93), .B1(new_n592), .B2(new_n596), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n536), .A2(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(G57gat), .A2(G64gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(G57gat), .A2(G64gat), .ZN(new_n602));
  INV_X1    g401(.A(G71gat), .ZN(new_n603));
  INV_X1    g402(.A(G78gat), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n601), .B(new_n602), .C1(new_n605), .C2(KEYINPUT9), .ZN(new_n606));
  XOR2_X1   g405(.A(G71gat), .B(G78gat), .Z(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n586), .B1(KEYINPUT21), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n612));
  INV_X1    g411(.A(KEYINPUT94), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT21), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n613), .B1(new_n608), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n608), .A2(new_n613), .A3(new_n614), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n616), .A2(G231gat), .A3(G233gat), .A4(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619));
  INV_X1    g418(.A(new_n617), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n619), .B1(new_n620), .B2(new_n615), .ZN(new_n621));
  XNOR2_X1  g420(.A(G127gat), .B(G155gat), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n618), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n622), .B1(new_n618), .B2(new_n621), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n612), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n625), .ZN(new_n627));
  INV_X1    g426(.A(new_n612), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n627), .A2(new_n623), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n611), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n626), .A2(new_n629), .A3(new_n611), .ZN(new_n632));
  XOR2_X1   g431(.A(G183gat), .B(G211gat), .Z(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n631), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n632), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n633), .B1(new_n636), .B2(new_n630), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(G134gat), .B(G162gat), .Z(new_n639));
  AND2_X1   g438(.A1(G232gat), .A2(G233gat), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n640), .A2(KEYINPUT41), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n639), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(G99gat), .A2(G106gat), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n643), .A2(KEYINPUT8), .ZN(new_n644));
  NOR2_X1   g443(.A1(G85gat), .A2(G92gat), .ZN(new_n645));
  OAI21_X1  g444(.A(KEYINPUT95), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n645), .B1(KEYINPUT8), .B2(new_n643), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT95), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(G85gat), .A2(G92gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT7), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(G99gat), .B(G106gat), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT96), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  OR2_X1    g455(.A1(G99gat), .A2(G106gat), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n657), .A2(KEYINPUT96), .A3(new_n643), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n653), .A2(new_n660), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n644), .A2(KEYINPUT95), .A3(new_n645), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n647), .A2(new_n648), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n659), .B(new_n652), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n572), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n640), .A2(KEYINPUT41), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n667), .B1(new_n580), .B2(new_n665), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(G190gat), .B(G218gat), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n666), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n642), .B1(new_n672), .B2(KEYINPUT97), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n661), .A2(new_n664), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n674), .B1(new_n568), .B2(new_n571), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n670), .B1(new_n675), .B2(new_n668), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n672), .B(new_n676), .C1(KEYINPUT97), .C2(new_n642), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(G120gat), .B(G148gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(G176gat), .B(G204gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(G230gat), .A2(G233gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT99), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT10), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT98), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n664), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n661), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n653), .A2(new_n688), .A3(new_n660), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n608), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n665), .A2(new_n609), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n687), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n665), .A2(new_n687), .A3(new_n608), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n686), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n659), .B1(new_n650), .B2(new_n652), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n699), .B1(new_n688), .B2(new_n664), .ZN(new_n700));
  INV_X1    g499(.A(new_n691), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n609), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n685), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n674), .A2(new_n608), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n684), .B1(new_n698), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(KEYINPUT100), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n703), .B1(new_n694), .B2(new_n696), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(new_n684), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n705), .ZN(new_n712));
  OAI211_X1 g511(.A(KEYINPUT100), .B(new_n683), .C1(new_n697), .C2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n707), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n638), .A2(new_n680), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(KEYINPUT101), .ZN(new_n717));
  OR2_X1    g516(.A1(new_n716), .A2(KEYINPUT101), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n600), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n719), .A2(new_n504), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(new_n574), .ZN(G1324gat));
  NOR2_X1   g520(.A1(new_n719), .A2(new_n492), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n722), .A2(KEYINPUT102), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n722), .A2(KEYINPUT102), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT42), .ZN(new_n725));
  OAI22_X1  g524(.A1(new_n723), .A2(new_n724), .B1(new_n725), .B2(G8gat), .ZN(new_n726));
  XOR2_X1   g525(.A(KEYINPUT16), .B(G8gat), .Z(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(KEYINPUT42), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n727), .A2(KEYINPUT42), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n728), .B1(new_n722), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n726), .A2(new_n730), .ZN(G1325gat));
  AND2_X1   g530(.A1(new_n498), .A2(new_n499), .ZN(new_n732));
  OAI21_X1  g531(.A(G15gat), .B1(new_n719), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n416), .ZN(new_n734));
  OR2_X1    g533(.A1(new_n734), .A2(G15gat), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n733), .B1(new_n719), .B2(new_n735), .ZN(G1326gat));
  OR3_X1    g535(.A1(new_n719), .A2(KEYINPUT103), .A3(new_n305), .ZN(new_n737));
  OAI21_X1  g536(.A(KEYINPUT103), .B1(new_n719), .B2(new_n305), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT43), .B(G22gat), .Z(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1327gat));
  INV_X1    g540(.A(new_n715), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n638), .A2(new_n680), .A3(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT104), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n600), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n504), .A2(G29gat), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT105), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT105), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n746), .A2(new_n750), .A3(new_n747), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT45), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT106), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n678), .A2(new_n756), .A3(new_n679), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n756), .B1(new_n678), .B2(new_n679), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n755), .B1(new_n536), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n305), .A2(new_n516), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n525), .A2(new_n534), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n732), .B1(new_n305), .B2(new_n483), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT35), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n734), .B1(new_n297), .B2(new_n304), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n766), .B1(new_n767), .B2(new_n483), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n491), .A2(new_n492), .A3(new_n416), .A4(new_n493), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n503), .A2(new_n769), .ZN(new_n770));
  OAI22_X1  g569(.A1(new_n764), .A2(new_n765), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n680), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n771), .A2(KEYINPUT44), .A3(new_n772), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n761), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n592), .A2(new_n596), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n638), .A2(new_n742), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(G29gat), .B1(new_n778), .B2(new_n504), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n749), .A2(KEYINPUT45), .A3(new_n751), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n754), .A2(new_n779), .A3(new_n780), .ZN(G1328gat));
  OAI21_X1  g580(.A(G36gat), .B1(new_n778), .B2(new_n492), .ZN(new_n782));
  INV_X1    g581(.A(G36gat), .ZN(new_n783));
  INV_X1    g582(.A(new_n492), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n746), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n785), .A2(KEYINPUT46), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT107), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n785), .A2(new_n787), .A3(KEYINPUT46), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n787), .B1(new_n785), .B2(KEYINPUT46), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n782), .B(new_n786), .C1(new_n788), .C2(new_n789), .ZN(G1329gat));
  NOR2_X1   g589(.A1(new_n734), .A2(G43gat), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n600), .A2(new_n744), .A3(new_n791), .ZN(new_n792));
  MUX2_X1   g591(.A(KEYINPUT108), .B(new_n792), .S(KEYINPUT47), .Z(new_n793));
  NAND4_X1  g592(.A1(new_n761), .A2(new_n773), .A3(new_n500), .A4(new_n777), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(G43gat), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n795), .A2(KEYINPUT108), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n792), .B(KEYINPUT109), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n796), .B1(new_n799), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g599(.A1(new_n503), .A2(G50gat), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n745), .A2(new_n305), .ZN(new_n802));
  OAI22_X1  g601(.A1(new_n778), .A2(new_n801), .B1(G50gat), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g603(.A(new_n638), .ZN(new_n805));
  NOR4_X1   g604(.A1(new_n805), .A2(new_n775), .A3(new_n772), .A4(new_n715), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n771), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n807), .A2(new_n504), .ZN(new_n808));
  XOR2_X1   g607(.A(new_n808), .B(G57gat), .Z(G1332gat));
  INV_X1    g608(.A(new_n807), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n784), .ZN(new_n811));
  NOR2_X1   g610(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n812));
  AND2_X1   g611(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n812), .B2(new_n811), .ZN(G1333gat));
  NOR3_X1   g614(.A1(new_n807), .A2(new_n603), .A3(new_n732), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n810), .A2(new_n416), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n816), .B1(new_n603), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g617(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n818), .B(new_n819), .ZN(G1334gat));
  NOR2_X1   g619(.A1(new_n807), .A2(new_n305), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(new_n604), .ZN(G1335gat));
  NOR3_X1   g621(.A1(new_n504), .A2(new_n715), .A3(G85gat), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT51), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n771), .A2(KEYINPUT112), .A3(new_n772), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n638), .A2(new_n775), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(KEYINPUT112), .B1(new_n771), .B2(new_n772), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n824), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n826), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n485), .A2(new_n495), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n506), .A2(new_n535), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n680), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n830), .B1(new_n833), .B2(KEYINPUT112), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT112), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n835), .B1(new_n536), .B2(new_n680), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(KEYINPUT51), .A3(new_n836), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n829), .A2(KEYINPUT113), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT113), .B1(new_n829), .B2(new_n837), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n823), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n826), .A2(new_n742), .ZN(new_n841));
  XOR2_X1   g640(.A(new_n841), .B(KEYINPUT111), .Z(new_n842));
  NAND2_X1  g641(.A1(new_n774), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(G85gat), .B1(new_n843), .B2(new_n504), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n840), .A2(new_n844), .ZN(G1336gat));
  NOR2_X1   g644(.A1(KEYINPUT114), .A2(KEYINPUT52), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n715), .A2(new_n492), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(G92gat), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n850), .B1(new_n829), .B2(new_n837), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n761), .A2(new_n773), .A3(new_n784), .A4(new_n842), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(G92gat), .ZN(new_n853));
  NAND2_X1  g652(.A1(KEYINPUT114), .A2(KEYINPUT52), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n846), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n827), .A2(new_n824), .A3(new_n828), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT51), .B1(new_n834), .B2(new_n836), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n849), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n846), .ZN(new_n860));
  AOI22_X1  g659(.A1(new_n852), .A2(G92gat), .B1(KEYINPUT114), .B2(KEYINPUT52), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n856), .A2(new_n862), .ZN(G1337gat));
  NOR3_X1   g662(.A1(new_n734), .A2(new_n715), .A3(G99gat), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n864), .B1(new_n838), .B2(new_n839), .ZN(new_n865));
  OAI21_X1  g664(.A(G99gat), .B1(new_n843), .B2(new_n732), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(G1338gat));
  NOR3_X1   g666(.A1(new_n305), .A2(G106gat), .A3(new_n715), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n869), .B1(new_n829), .B2(new_n837), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n761), .A2(new_n773), .A3(new_n503), .A4(new_n842), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(G106gat), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n871), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n874), .ZN(new_n876));
  OAI21_X1  g675(.A(KEYINPUT53), .B1(new_n870), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n877), .ZN(G1339gat));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n684), .B1(new_n697), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n694), .A2(new_n696), .A3(new_n686), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n702), .A2(new_n704), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n695), .B1(new_n882), .B2(new_n687), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n881), .B(KEYINPUT54), .C1(new_n883), .C2(new_n703), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT55), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n880), .A2(new_n884), .A3(KEYINPUT55), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n887), .A2(new_n775), .A3(new_n711), .A4(new_n888), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n590), .A2(new_n579), .ZN(new_n890));
  OR3_X1    g689(.A1(new_n587), .A2(new_n581), .A3(new_n584), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n543), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n589), .A2(new_n591), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n892), .B1(new_n893), .B2(new_n546), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n894), .B1(new_n707), .B2(new_n714), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n759), .B1(new_n889), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n680), .A2(KEYINPUT106), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n678), .A2(new_n756), .A3(new_n679), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n897), .A2(new_n898), .A3(new_n894), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n710), .B1(new_n885), .B2(new_n886), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n888), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n805), .B1(new_n896), .B2(new_n902), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n638), .A2(new_n776), .A3(new_n680), .A4(new_n715), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n784), .A2(new_n504), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n907), .A2(new_n767), .ZN(new_n908));
  INV_X1    g707(.A(new_n599), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n363), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  XOR2_X1   g709(.A(new_n910), .B(KEYINPUT115), .Z(new_n911));
  NAND3_X1  g710(.A1(new_n908), .A2(new_n363), .A3(new_n775), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1340gat));
  NAND2_X1  g712(.A1(new_n908), .A2(new_n742), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT116), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n914), .A2(new_n915), .A3(new_n361), .ZN(new_n916));
  XOR2_X1   g715(.A(KEYINPUT116), .B(G120gat), .Z(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n914), .B2(new_n917), .ZN(G1341gat));
  NAND2_X1  g717(.A1(new_n908), .A2(new_n638), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g719(.A1(new_n907), .A2(new_n772), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(new_n767), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(G134gat), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT117), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n369), .A2(new_n370), .ZN(new_n926));
  OAI21_X1  g725(.A(KEYINPUT56), .B1(new_n923), .B2(new_n926), .ZN(new_n927));
  OR3_X1    g726(.A1(new_n923), .A2(KEYINPUT56), .A3(new_n926), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n925), .A2(new_n927), .A3(new_n928), .ZN(G1343gat));
  NAND2_X1  g728(.A1(new_n732), .A2(new_n906), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n503), .A2(KEYINPUT57), .ZN(new_n932));
  INV_X1    g731(.A(new_n904), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n900), .B(new_n888), .C1(new_n597), .C2(new_n598), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n772), .B1(new_n934), .B2(new_n895), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n805), .B1(new_n935), .B2(new_n902), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n933), .B1(new_n936), .B2(KEYINPUT118), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT118), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n938), .B(new_n805), .C1(new_n935), .C2(new_n902), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n932), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT57), .B1(new_n905), .B2(new_n503), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n931), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(G141gat), .B1(new_n942), .B2(new_n599), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT58), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n500), .A2(new_n305), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n907), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n909), .A2(new_n225), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n943), .A2(new_n944), .A3(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT119), .ZN(new_n951));
  OAI211_X1 g750(.A(new_n775), .B(new_n931), .C1(new_n940), .C2(new_n941), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(G141gat), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(new_n949), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n951), .B1(new_n954), .B2(KEYINPUT58), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n948), .B1(new_n952), .B2(G141gat), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n956), .A2(KEYINPUT119), .A3(new_n944), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n950), .B1(new_n955), .B2(new_n957), .ZN(G1344gat));
  INV_X1    g757(.A(new_n946), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n959), .A2(new_n228), .A3(new_n742), .ZN(new_n960));
  XNOR2_X1  g759(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n718), .A2(new_n599), .A3(new_n717), .ZN(new_n962));
  AND4_X1   g761(.A1(new_n772), .A2(new_n900), .A3(new_n888), .A4(new_n894), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n805), .B1(new_n935), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT57), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n965), .A2(new_n966), .A3(new_n503), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n905), .A2(new_n503), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(KEYINPUT57), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n967), .A2(new_n742), .A3(new_n969), .ZN(new_n970));
  OR2_X1    g769(.A1(new_n970), .A2(new_n930), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n961), .B1(new_n971), .B2(G148gat), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n942), .A2(new_n715), .ZN(new_n973));
  NOR3_X1   g772(.A1(new_n973), .A2(KEYINPUT59), .A3(new_n228), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n960), .B1(new_n972), .B2(new_n974), .ZN(G1345gat));
  OAI21_X1  g774(.A(G155gat), .B1(new_n942), .B2(new_n805), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n959), .A2(new_n235), .A3(new_n638), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(G1346gat));
  OAI21_X1  g777(.A(G162gat), .B1(new_n942), .B2(new_n760), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n922), .A2(new_n236), .A3(new_n945), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(G1347gat));
  NAND3_X1  g780(.A1(new_n784), .A2(new_n504), .A3(new_n416), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT121), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n305), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n984), .B1(new_n983), .B2(new_n982), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n985), .A2(new_n905), .ZN(new_n986));
  NOR3_X1   g785(.A1(new_n986), .A2(new_n539), .A3(new_n599), .ZN(new_n987));
  AND2_X1   g786(.A1(new_n905), .A2(new_n504), .ZN(new_n988));
  AND3_X1   g787(.A1(new_n988), .A2(new_n784), .A3(new_n767), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n989), .A2(new_n775), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n987), .B1(new_n990), .B2(new_n539), .ZN(G1348gat));
  AOI21_X1  g790(.A(G176gat), .B1(new_n989), .B2(new_n742), .ZN(new_n992));
  OR3_X1    g791(.A1(new_n986), .A2(new_n347), .A3(new_n715), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT122), .ZN(new_n994));
  OR2_X1    g793(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n993), .A2(new_n994), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n992), .B1(new_n995), .B2(new_n996), .ZN(G1349gat));
  NAND3_X1  g796(.A1(new_n989), .A2(new_n308), .A3(new_n638), .ZN(new_n998));
  OAI21_X1  g797(.A(G183gat), .B1(new_n986), .B2(new_n805), .ZN(new_n999));
  NAND2_X1  g798(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  NOR2_X1   g800(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n1002));
  XOR2_X1   g801(.A(new_n1001), .B(new_n1002), .Z(G1350gat));
  NAND3_X1  g802(.A1(new_n989), .A2(new_n307), .A3(new_n759), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n985), .A2(new_n772), .A3(new_n905), .ZN(new_n1005));
  INV_X1    g804(.A(KEYINPUT61), .ZN(new_n1006));
  AND3_X1   g805(.A1(new_n1005), .A2(new_n1006), .A3(G190gat), .ZN(new_n1007));
  AOI21_X1  g806(.A(new_n1006), .B1(new_n1005), .B2(G190gat), .ZN(new_n1008));
  OAI21_X1  g807(.A(new_n1004), .B1(new_n1007), .B2(new_n1008), .ZN(G1351gat));
  AND2_X1   g808(.A1(new_n988), .A2(new_n945), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1010), .A2(new_n784), .ZN(new_n1011));
  XNOR2_X1  g810(.A(KEYINPUT124), .B(G197gat), .ZN(new_n1012));
  OR3_X1    g811(.A1(new_n1011), .A2(new_n776), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n784), .A2(new_n504), .ZN(new_n1014));
  NOR2_X1   g813(.A1(new_n1014), .A2(new_n500), .ZN(new_n1015));
  AND3_X1   g814(.A1(new_n967), .A2(new_n969), .A3(new_n1015), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n1016), .A2(KEYINPUT125), .A3(new_n909), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1017), .A2(new_n1012), .ZN(new_n1018));
  AOI21_X1  g817(.A(KEYINPUT125), .B1(new_n1016), .B2(new_n909), .ZN(new_n1019));
  OAI21_X1  g818(.A(new_n1013), .B1(new_n1018), .B2(new_n1019), .ZN(G1352gat));
  NAND3_X1  g819(.A1(new_n1010), .A2(new_n210), .A3(new_n847), .ZN(new_n1021));
  XOR2_X1   g820(.A(new_n1021), .B(KEYINPUT62), .Z(new_n1022));
  NOR3_X1   g821(.A1(new_n970), .A2(new_n500), .A3(new_n1014), .ZN(new_n1023));
  OAI21_X1  g822(.A(new_n1022), .B1(new_n1023), .B2(new_n210), .ZN(G1353gat));
  INV_X1    g823(.A(G211gat), .ZN(new_n1025));
  AOI21_X1  g824(.A(new_n1025), .B1(new_n1016), .B2(new_n638), .ZN(new_n1026));
  INV_X1    g825(.A(KEYINPUT63), .ZN(new_n1027));
  OR2_X1    g826(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g827(.A1(new_n1010), .A2(new_n1025), .A3(new_n784), .A4(new_n638), .ZN(new_n1029));
  XNOR2_X1  g828(.A(new_n1029), .B(KEYINPUT126), .ZN(new_n1030));
  NAND2_X1  g829(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1031));
  NAND3_X1  g830(.A1(new_n1028), .A2(new_n1030), .A3(new_n1031), .ZN(G1354gat));
  INV_X1    g831(.A(G218gat), .ZN(new_n1033));
  NAND4_X1  g832(.A1(new_n1010), .A2(new_n1033), .A3(new_n784), .A4(new_n759), .ZN(new_n1034));
  AND2_X1   g833(.A1(new_n1016), .A2(new_n772), .ZN(new_n1035));
  OAI211_X1 g834(.A(new_n1034), .B(KEYINPUT127), .C1(new_n1035), .C2(new_n1033), .ZN(new_n1036));
  INV_X1    g835(.A(KEYINPUT127), .ZN(new_n1037));
  AOI21_X1  g836(.A(new_n1033), .B1(new_n1016), .B2(new_n772), .ZN(new_n1038));
  INV_X1    g837(.A(new_n1034), .ZN(new_n1039));
  OAI21_X1  g838(.A(new_n1037), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g839(.A1(new_n1036), .A2(new_n1040), .ZN(G1355gat));
endmodule


