//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1287, new_n1288, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1342, new_n1343, new_n1344;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND3_X1  g0009(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(G58), .A2(G68), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G50), .ZN(new_n213));
  XNOR2_X1  g0013(.A(KEYINPUT64), .B(G68), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G58), .A2(G232), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n206), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n209), .B1(new_n210), .B2(new_n213), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT2), .B(G226), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n228), .B(new_n229), .Z(new_n230));
  XOR2_X1   g0030(.A(G264), .B(G270), .Z(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XOR2_X1   g0034(.A(G50), .B(G58), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT65), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G68), .B(G77), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  INV_X1    g0042(.A(KEYINPUT66), .ZN(new_n243));
  AND2_X1   g0043(.A1(G33), .A2(G41), .ZN(new_n244));
  NAND2_X1  g0044(.A1(G1), .A2(G13), .ZN(new_n245));
  OAI21_X1  g0045(.A(G274), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  OAI21_X1  g0046(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n247));
  OAI21_X1  g0047(.A(new_n243), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  INV_X1    g0049(.A(G41), .ZN(new_n250));
  OAI211_X1 g0050(.A(G1), .B(G13), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G45), .ZN(new_n252));
  AOI21_X1  g0052(.A(G1), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  NAND4_X1  g0053(.A1(new_n251), .A2(KEYINPUT66), .A3(new_n253), .A4(G274), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n248), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT70), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT70), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n248), .A2(new_n257), .A3(new_n254), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n251), .A2(new_n247), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(new_n216), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT67), .B(G1698), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n262), .A2(G226), .B1(G232), .B2(G1698), .ZN(new_n263));
  AND2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G97), .ZN(new_n267));
  OAI22_X1  g0067(.A1(new_n263), .A2(new_n266), .B1(new_n249), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n244), .A2(new_n245), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n261), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT13), .ZN(new_n271));
  AND3_X1   g0071(.A1(new_n259), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n271), .B1(new_n259), .B2(new_n270), .ZN(new_n273));
  OAI21_X1  g0073(.A(G169), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT14), .ZN(new_n275));
  AND3_X1   g0075(.A1(new_n248), .A2(new_n257), .A3(new_n254), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n257), .B1(new_n248), .B2(new_n254), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n249), .A2(new_n267), .ZN(new_n279));
  INV_X1    g0079(.A(G1698), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT67), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT67), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G1698), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G226), .ZN(new_n285));
  OAI22_X1  g0085(.A1(new_n284), .A2(new_n285), .B1(new_n227), .B2(new_n280), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT3), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n249), .ZN(new_n288));
  NAND2_X1  g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n279), .B1(new_n286), .B2(new_n290), .ZN(new_n291));
  OAI22_X1  g0091(.A1(new_n291), .A2(new_n251), .B1(new_n216), .B2(new_n260), .ZN(new_n292));
  OAI21_X1  g0092(.A(KEYINPUT13), .B1(new_n278), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT71), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n259), .A2(new_n270), .A3(new_n271), .ZN(new_n296));
  OAI211_X1 g0096(.A(KEYINPUT71), .B(KEYINPUT13), .C1(new_n278), .C2(new_n292), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n295), .A2(G179), .A3(new_n296), .A4(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n293), .A2(new_n296), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT14), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(new_n300), .A3(G169), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n275), .A2(new_n298), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G13), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(G1), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G20), .ZN(new_n305));
  OAI21_X1  g0105(.A(KEYINPUT12), .B1(new_n305), .B2(new_n214), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n306), .B(KEYINPUT72), .ZN(new_n307));
  OR2_X1    g0107(.A1(KEYINPUT12), .A2(G68), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n307), .B1(new_n305), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n245), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n214), .A2(new_n204), .ZN(new_n312));
  NOR2_X1   g0112(.A1(G20), .A2(G33), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G50), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n204), .A2(G33), .ZN(new_n316));
  INV_X1    g0116(.A(G77), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n314), .A2(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n311), .B1(new_n312), .B2(new_n318), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n319), .B(KEYINPUT11), .ZN(new_n320));
  NOR3_X1   g0120(.A1(new_n303), .A2(new_n204), .A3(G1), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n321), .A2(new_n311), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n203), .A2(G20), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n322), .A2(G68), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n309), .A2(new_n320), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n302), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n325), .B1(new_n299), .B2(G200), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n295), .A2(G190), .A3(new_n296), .A4(new_n297), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT73), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n326), .A2(KEYINPUT73), .A3(new_n329), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT16), .ZN(new_n334));
  INV_X1    g0134(.A(G159), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n314), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n211), .B1(new_n214), .B2(G58), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n337), .B1(new_n338), .B2(new_n204), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n288), .A2(new_n204), .A3(new_n289), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT7), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n288), .A2(KEYINPUT7), .A3(new_n204), .A4(new_n289), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n215), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n334), .B1(new_n339), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT75), .ZN(new_n346));
  AND2_X1   g0146(.A1(KEYINPUT64), .A2(G68), .ZN(new_n347));
  NOR2_X1   g0147(.A1(KEYINPUT64), .A2(G68), .ZN(new_n348));
  OAI21_X1  g0148(.A(G58), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n204), .B1(new_n349), .B2(new_n212), .ZN(new_n350));
  OAI21_X1  g0150(.A(KEYINPUT74), .B1(new_n350), .B2(new_n336), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT74), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n352), .B(new_n337), .C1(new_n338), .C2(new_n204), .ZN(new_n353));
  AOI21_X1  g0153(.A(KEYINPUT7), .B1(new_n266), .B2(new_n204), .ZN(new_n354));
  INV_X1    g0154(.A(new_n343), .ZN(new_n355));
  OAI21_X1  g0155(.A(G68), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n351), .A2(new_n353), .A3(KEYINPUT16), .A4(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT75), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n358), .B(new_n334), .C1(new_n339), .C2(new_n344), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n346), .A2(new_n311), .A3(new_n357), .A4(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n322), .ZN(new_n361));
  XOR2_X1   g0161(.A(KEYINPUT8), .B(G58), .Z(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n323), .ZN(new_n363));
  OAI22_X1  g0163(.A1(new_n361), .A2(new_n363), .B1(new_n305), .B2(new_n362), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n260), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(G232), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n255), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT76), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n248), .A2(new_n254), .B1(new_n367), .B2(G232), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT76), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n290), .A2(G226), .A3(G1698), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G33), .A2(G87), .ZN(new_n375));
  INV_X1    g0175(.A(G223), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n281), .B(new_n283), .C1(new_n264), .C2(new_n265), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n374), .B(new_n375), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(G179), .B1(new_n378), .B2(new_n269), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n370), .A2(new_n373), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT77), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n378), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n371), .B1(new_n383), .B2(new_n251), .ZN(new_n384));
  INV_X1    g0184(.A(G169), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n370), .A2(new_n373), .A3(KEYINPUT77), .A4(new_n379), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n382), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(KEYINPUT18), .B1(new_n366), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G200), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n384), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(G190), .B1(new_n378), .B2(new_n269), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n370), .A2(new_n373), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n366), .A2(KEYINPUT17), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n360), .A2(new_n365), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n387), .A2(new_n386), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT18), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n396), .A2(new_n397), .A3(new_n398), .A4(new_n382), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n394), .A2(new_n360), .A3(new_n365), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT17), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n389), .A2(new_n395), .A3(new_n399), .A4(new_n402), .ZN(new_n403));
  XNOR2_X1  g0203(.A(KEYINPUT8), .B(G58), .ZN(new_n404));
  INV_X1    g0204(.A(G150), .ZN(new_n405));
  OAI22_X1  g0205(.A1(new_n404), .A2(new_n316), .B1(new_n405), .B2(new_n314), .ZN(new_n406));
  NOR2_X1   g0206(.A1(G50), .A2(G58), .ZN(new_n407));
  INV_X1    g0207(.A(G68), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n204), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n311), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n315), .B1(new_n203), .B2(G20), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n322), .A2(new_n411), .B1(new_n315), .B2(new_n321), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT9), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT9), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT10), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n280), .B1(new_n288), .B2(new_n289), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(G223), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(new_n317), .B2(new_n290), .ZN(new_n422));
  INV_X1    g0222(.A(G222), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n377), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n269), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n248), .A2(new_n254), .B1(new_n367), .B2(G226), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(G190), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n426), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(G200), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n418), .A2(new_n419), .A3(new_n427), .A4(new_n429), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n429), .A2(new_n427), .A3(new_n417), .A4(new_n415), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT10), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT69), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n367), .A2(G244), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n255), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT68), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n420), .A2(G238), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n266), .A2(G107), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n438), .B(new_n439), .C1(new_n227), .C2(new_n377), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n436), .A2(new_n437), .B1(new_n269), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n255), .A2(KEYINPUT68), .A3(new_n435), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n390), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n322), .A2(G77), .A3(new_n323), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(G77), .B2(new_n305), .ZN(new_n445));
  INV_X1    g0245(.A(new_n311), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n362), .A2(new_n313), .B1(G20), .B2(G77), .ZN(new_n447));
  XNOR2_X1  g0247(.A(KEYINPUT15), .B(G87), .ZN(new_n448));
  OR2_X1    g0248(.A1(new_n448), .A2(new_n316), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n446), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n434), .B1(new_n443), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n436), .A2(new_n437), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n440), .A2(new_n269), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n454), .A2(new_n442), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G200), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n457), .A2(KEYINPUT69), .A3(new_n451), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n441), .A2(G190), .A3(new_n442), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n453), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n456), .A2(new_n385), .ZN(new_n461));
  INV_X1    g0261(.A(G179), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n441), .A2(new_n462), .A3(new_n442), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n461), .A2(new_n452), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n428), .A2(new_n385), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n465), .B(new_n413), .C1(G179), .C2(new_n428), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n433), .A2(new_n460), .A3(new_n464), .A4(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n403), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n332), .A2(new_n333), .A3(new_n468), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n203), .B(G45), .C1(new_n250), .C2(KEYINPUT5), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT79), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT5), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G41), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n474), .A2(KEYINPUT79), .A3(new_n203), .A4(G45), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n250), .A2(KEYINPUT5), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n472), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n477), .A2(G270), .A3(new_n251), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT81), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n470), .A2(new_n471), .B1(KEYINPUT5), .B2(new_n250), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n480), .A2(G274), .A3(new_n251), .A4(new_n475), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT81), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n477), .A2(new_n482), .A3(G270), .A4(new_n251), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G283), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n485), .B(new_n204), .C1(G33), .C2(new_n267), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT82), .ZN(new_n487));
  AOI21_X1  g0287(.A(G20), .B1(new_n249), .B2(G97), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT82), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(new_n489), .A3(new_n485), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(G116), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n310), .A2(new_n245), .B1(G20), .B2(new_n492), .ZN(new_n493));
  AND3_X1   g0293(.A1(new_n491), .A2(KEYINPUT20), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(KEYINPUT20), .B1(new_n491), .B2(new_n493), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n446), .B(new_n305), .C1(G1), .C2(new_n249), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n496), .A2(G116), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n321), .A2(G116), .ZN(new_n498));
  OAI22_X1  g0298(.A1(new_n494), .A2(new_n495), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n290), .A2(new_n262), .A3(G257), .ZN(new_n500));
  OAI211_X1 g0300(.A(G264), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n288), .A2(G303), .A3(new_n289), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n462), .B1(new_n503), .B2(new_n269), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n484), .A2(new_n499), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n503), .A2(new_n269), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n479), .A2(new_n506), .A3(new_n481), .A4(new_n483), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n507), .A2(new_n499), .A3(KEYINPUT21), .A4(G169), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n499), .B1(new_n507), .B2(G200), .ZN(new_n510));
  INV_X1    g0310(.A(G190), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n510), .B1(new_n511), .B2(new_n507), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n507), .A2(new_n499), .A3(G169), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT21), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n513), .A2(KEYINPUT83), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(KEYINPUT83), .B1(new_n513), .B2(new_n514), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n509), .B(new_n512), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(G107), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n321), .A2(new_n518), .ZN(new_n519));
  XOR2_X1   g0319(.A(KEYINPUT84), .B(KEYINPUT25), .Z(new_n520));
  XNOR2_X1  g0320(.A(new_n519), .B(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n496), .A2(new_n518), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n290), .A2(new_n204), .A3(G87), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT22), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT22), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n290), .A2(new_n527), .A3(new_n204), .A4(G87), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G33), .A2(G116), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n530), .A2(G20), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT23), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(new_n204), .B2(G107), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n518), .A2(KEYINPUT23), .A3(G20), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n529), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(KEYINPUT24), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT24), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n529), .A2(new_n538), .A3(new_n535), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n524), .B1(new_n540), .B2(new_n311), .ZN(new_n541));
  OAI211_X1 g0341(.A(G257), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G294), .ZN(new_n543));
  INV_X1    g0343(.A(G250), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n542), .B(new_n543), .C1(new_n377), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n269), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n477), .A2(G264), .A3(new_n251), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n546), .A2(new_n547), .A3(new_n481), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n548), .A2(KEYINPUT86), .A3(new_n390), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n546), .A2(KEYINPUT85), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT85), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n545), .A2(new_n551), .A3(new_n269), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n550), .A2(new_n481), .A3(new_n552), .A4(new_n547), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n549), .B1(new_n553), .B2(G190), .ZN(new_n554));
  AOI21_X1  g0354(.A(KEYINPUT86), .B1(new_n548), .B2(new_n390), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n541), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n553), .A2(G169), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n269), .B1(new_n480), .B2(new_n475), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n558), .A2(G264), .B1(new_n545), .B2(new_n269), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n559), .A2(G179), .A3(new_n481), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n539), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n538), .B1(new_n529), .B2(new_n535), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n311), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n523), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n556), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(G244), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n530), .B(new_n568), .C1(new_n377), .C2(new_n216), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n269), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n544), .B1(new_n252), .B2(G1), .ZN(new_n571));
  INV_X1    g0371(.A(G274), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n203), .A2(new_n572), .A3(G45), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n251), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT80), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT80), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n570), .A2(new_n577), .A3(new_n574), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n462), .A3(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n448), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n580), .A2(new_n305), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n290), .A2(new_n204), .A3(G68), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n316), .A2(new_n267), .ZN(new_n583));
  AOI21_X1  g0383(.A(G20), .B1(new_n279), .B2(KEYINPUT19), .ZN(new_n584));
  NOR3_X1   g0384(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n585));
  OAI221_X1 g0385(.A(new_n582), .B1(KEYINPUT19), .B2(new_n583), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n581), .B1(new_n586), .B2(new_n311), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(new_n448), .B2(new_n496), .ZN(new_n588));
  INV_X1    g0388(.A(new_n574), .ZN(new_n589));
  AOI211_X1 g0389(.A(KEYINPUT80), .B(new_n589), .C1(new_n569), .C2(new_n269), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n577), .B1(new_n570), .B2(new_n574), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n579), .B(new_n588), .C1(new_n592), .C2(G169), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n576), .A2(G190), .A3(new_n578), .ZN(new_n594));
  OAI21_X1  g0394(.A(G200), .B1(new_n590), .B2(new_n591), .ZN(new_n595));
  INV_X1    g0395(.A(G87), .ZN(new_n596));
  OR2_X1    g0396(.A1(new_n496), .A2(new_n596), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n587), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n594), .A2(new_n595), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n477), .A2(G257), .A3(new_n251), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n600), .A2(new_n481), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT4), .ZN(new_n602));
  INV_X1    g0402(.A(G244), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n602), .B1(new_n377), .B2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n290), .A2(new_n262), .A3(KEYINPUT4), .A4(G244), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n420), .A2(G250), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n604), .A2(new_n485), .A3(new_n605), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n269), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n601), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n385), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n601), .A2(new_n608), .A3(new_n462), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT6), .ZN(new_n612));
  NOR3_X1   g0412(.A1(new_n612), .A2(new_n267), .A3(G107), .ZN(new_n613));
  XNOR2_X1  g0413(.A(G97), .B(G107), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n613), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  OAI22_X1  g0415(.A1(new_n615), .A2(new_n204), .B1(new_n317), .B2(new_n314), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n518), .B1(new_n342), .B2(new_n343), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n311), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(KEYINPUT78), .B1(new_n305), .B2(G97), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT78), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n321), .A2(new_n620), .A3(new_n267), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n618), .B(new_n622), .C1(new_n267), .C2(new_n496), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n610), .A2(new_n611), .A3(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n622), .B1(new_n267), .B2(new_n496), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n614), .A2(new_n612), .ZN(new_n626));
  INV_X1    g0426(.A(new_n613), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n628), .A2(G20), .B1(G77), .B2(new_n313), .ZN(new_n629));
  INV_X1    g0429(.A(new_n617), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n625), .B1(new_n631), .B2(new_n311), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n601), .A2(new_n608), .A3(G190), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n600), .A2(new_n481), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n634), .B1(new_n269), .B2(new_n607), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n632), .B(new_n633), .C1(new_n635), .C2(new_n390), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n593), .A2(new_n599), .A3(new_n624), .A4(new_n636), .ZN(new_n637));
  NOR4_X1   g0437(.A1(new_n469), .A2(new_n517), .A3(new_n567), .A4(new_n637), .ZN(G372));
  XNOR2_X1  g0438(.A(new_n433), .B(KEYINPUT91), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n464), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n329), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n326), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(KEYINPUT90), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n395), .A2(new_n402), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n302), .A2(new_n325), .B1(new_n329), .B2(new_n641), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT90), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n644), .A2(new_n646), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n389), .A2(new_n399), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n640), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n466), .ZN(new_n654));
  OAI21_X1  g0454(.A(KEYINPUT92), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT92), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n645), .B1(new_n643), .B2(KEYINPUT90), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n651), .B1(new_n657), .B2(new_n649), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n656), .B(new_n466), .C1(new_n658), .C2(new_n640), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n469), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n575), .A2(G200), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n594), .A2(new_n598), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n575), .A2(new_n385), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n579), .A2(new_n588), .A3(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT26), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT89), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n624), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n610), .A2(new_n623), .A3(KEYINPUT89), .A4(new_n611), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n666), .A2(new_n667), .A3(new_n669), .A4(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n611), .ZN(new_n672));
  AOI21_X1  g0472(.A(G169), .B1(new_n601), .B2(new_n608), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n672), .A2(new_n673), .A3(new_n632), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n674), .A2(new_n593), .A3(new_n599), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(KEYINPUT26), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n671), .A2(new_n665), .A3(new_n676), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n561), .A2(new_n565), .A3(KEYINPUT88), .ZN(new_n678));
  AOI21_X1  g0478(.A(KEYINPUT88), .B1(new_n561), .B2(new_n565), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n509), .B1(new_n515), .B2(new_n516), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT87), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OAI211_X1 g0483(.A(new_n509), .B(KEYINPUT87), .C1(new_n515), .C2(new_n516), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n680), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n624), .A2(new_n636), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n686), .A2(new_n666), .A3(new_n556), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n677), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n661), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n660), .A2(new_n689), .ZN(G369));
  INV_X1    g0490(.A(new_n517), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n304), .A2(new_n204), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(new_n694), .A3(G213), .ZN(new_n695));
  INV_X1    g0495(.A(G343), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n499), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n691), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n683), .A2(new_n684), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n699), .B1(new_n700), .B2(new_n698), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(G330), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n697), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n556), .B(new_n566), .C1(new_n541), .C2(new_n704), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT93), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n566), .B2(new_n704), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n680), .A2(new_n704), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n681), .A2(new_n704), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n708), .A2(new_n709), .A3(new_n711), .ZN(G399));
  INV_X1    g0512(.A(new_n207), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G41), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n585), .A2(new_n492), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(G1), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(new_n213), .B2(new_n715), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT94), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT28), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT29), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n688), .A2(new_n721), .A3(new_n704), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n674), .A2(new_n593), .A3(new_n599), .A4(new_n667), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n723), .A2(new_n665), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n669), .A2(new_n665), .A3(new_n663), .A4(new_n670), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(KEYINPUT26), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n566), .B(new_n509), .C1(new_n515), .C2(new_n516), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OAI211_X1 g0528(.A(new_n724), .B(new_n726), .C1(new_n728), .C2(new_n687), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n704), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT29), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n722), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n504), .A2(new_n546), .A3(new_n547), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n592), .A2(new_n484), .A3(new_n635), .A4(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT30), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AND4_X1   g0537(.A1(new_n504), .A2(new_n601), .A3(new_n559), .A4(new_n608), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n738), .A2(KEYINPUT30), .A3(new_n484), .A4(new_n592), .ZN(new_n739));
  AOI21_X1  g0539(.A(G179), .B1(new_n570), .B2(new_n574), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n609), .A2(new_n507), .A3(new_n548), .A4(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n737), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(new_n697), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT31), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n742), .A2(KEYINPUT31), .A3(new_n697), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR4_X1   g0547(.A1(new_n517), .A2(new_n567), .A3(new_n637), .A4(new_n697), .ZN(new_n748));
  OAI21_X1  g0548(.A(G330), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n733), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n720), .B1(new_n751), .B2(G1), .ZN(G364));
  NOR2_X1   g0552(.A1(new_n303), .A2(G20), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n203), .B1(new_n753), .B2(G45), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n714), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G13), .A2(G33), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n701), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n207), .A2(new_n290), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(KEYINPUT95), .B2(G355), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n764), .B1(KEYINPUT95), .B2(G355), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n238), .A2(new_n252), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n713), .A2(new_n290), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(G45), .B2(new_n213), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n765), .B1(G116), .B2(new_n207), .C1(new_n766), .C2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n245), .B1(G20), .B2(new_n385), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n760), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT96), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n204), .A2(new_n462), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n773), .A2(G190), .A3(new_n390), .ZN(new_n774));
  INV_X1    g0574(.A(G322), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G190), .A2(G200), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G311), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n266), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n204), .A2(G179), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n777), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n776), .B(new_n780), .C1(G329), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n773), .A2(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n511), .ZN(new_n786));
  XNOR2_X1  g0586(.A(KEYINPUT98), .B(G326), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n785), .A2(G190), .ZN(new_n789));
  XNOR2_X1  g0589(.A(KEYINPUT33), .B(G317), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n781), .A2(G190), .A3(G200), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n789), .A2(new_n790), .B1(new_n792), .B2(G303), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n781), .A2(new_n511), .A3(G200), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n462), .A2(new_n390), .A3(G190), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G20), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n795), .A2(G283), .B1(new_n797), .B2(G294), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n784), .A2(new_n788), .A3(new_n793), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n792), .A2(G87), .ZN(new_n800));
  XOR2_X1   g0600(.A(KEYINPUT97), .B(G159), .Z(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(new_n783), .ZN(new_n803));
  INV_X1    g0603(.A(new_n789), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n800), .B1(new_n803), .B2(KEYINPUT32), .C1(new_n408), .C2(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n290), .B1(new_n778), .B2(new_n317), .ZN(new_n806));
  INV_X1    g0606(.A(new_n774), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n806), .B1(G58), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n795), .A2(G107), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n803), .A2(KEYINPUT32), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n786), .A2(G50), .B1(G97), .B2(new_n797), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n799), .B1(new_n805), .B2(new_n812), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n769), .A2(new_n772), .B1(new_n770), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n757), .B1(new_n762), .B2(new_n814), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n701), .A2(G330), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n756), .B1(new_n816), .B2(new_n702), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT99), .ZN(G396));
  NAND2_X1  g0619(.A1(new_n464), .A2(KEYINPUT101), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT101), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n461), .A2(new_n821), .A3(new_n452), .A4(new_n463), .ZN(new_n822));
  AND3_X1   g0622(.A1(new_n460), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n823), .A2(new_n704), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n688), .A2(new_n824), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n688), .A2(new_n704), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n452), .A2(new_n697), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n460), .A2(new_n827), .A3(new_n820), .A4(new_n822), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n641), .A2(new_n697), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n825), .B1(new_n826), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n757), .B1(new_n832), .B2(new_n749), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT102), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n832), .B2(new_n749), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n832), .A2(new_n834), .A3(new_n749), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n830), .A2(new_n758), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n770), .A2(new_n758), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n756), .B1(G77), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n794), .A2(new_n596), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n791), .A2(new_n518), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n843), .B(new_n844), .C1(G303), .C2(new_n786), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n290), .B1(new_n807), .B2(G294), .ZN(new_n846));
  INV_X1    g0646(.A(new_n778), .ZN(new_n847));
  AOI22_X1  g0647(.A1(G116), .A2(new_n847), .B1(new_n783), .B2(G311), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n789), .A2(G283), .B1(G97), .B2(new_n797), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n845), .A2(new_n846), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n791), .A2(new_n315), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n795), .A2(G68), .ZN(new_n852));
  INV_X1    g0652(.A(G132), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n852), .B(new_n290), .C1(new_n853), .C2(new_n782), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n851), .B(new_n854), .C1(G58), .C2(new_n797), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT100), .ZN(new_n856));
  AOI22_X1  g0656(.A1(G143), .A2(new_n807), .B1(new_n802), .B2(new_n847), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(new_n405), .B2(new_n804), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(G137), .B2(new_n786), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT34), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n850), .B1(new_n856), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n842), .B1(new_n861), .B2(new_n770), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n839), .A2(new_n862), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n838), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(G384));
  NAND2_X1  g0665(.A1(new_n628), .A2(KEYINPUT35), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n210), .A2(new_n492), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n628), .B2(KEYINPUT35), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT103), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n866), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n869), .B2(new_n868), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(KEYINPUT36), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n349), .A2(G50), .A3(G77), .A4(new_n212), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n315), .A2(G68), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n203), .B(G13), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n742), .A2(KEYINPUT31), .A3(new_n697), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT31), .B1(new_n742), .B2(new_n697), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n567), .A2(new_n637), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n880), .A2(new_n691), .A3(new_n704), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n661), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT107), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n396), .A2(new_n397), .A3(new_n382), .ZN(new_n885));
  INV_X1    g0685(.A(new_n695), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT105), .B1(new_n396), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT105), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n888), .B(new_n695), .C1(new_n360), .C2(new_n365), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n885), .B(new_n400), .C1(new_n887), .C2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n396), .A2(new_n886), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n888), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n396), .A2(KEYINPUT105), .A3(new_n886), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n400), .B1(new_n366), .B2(new_n388), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT37), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n895), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n891), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n895), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n403), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT38), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n357), .A2(new_n311), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n351), .A2(new_n353), .A3(new_n356), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n334), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n364), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n400), .B1(new_n388), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n907), .A2(new_n695), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT37), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n890), .B2(KEYINPUT37), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n403), .A2(new_n909), .ZN(new_n912));
  AND3_X1   g0712(.A1(new_n911), .A2(KEYINPUT38), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT106), .B1(new_n903), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n830), .B1(new_n879), .B2(new_n881), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n325), .A2(new_n697), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n327), .A2(new_n328), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n916), .B1(new_n917), .B2(new_n302), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT104), .ZN(new_n919));
  INV_X1    g0719(.A(new_n916), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n326), .A2(new_n329), .A3(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT104), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n922), .B(new_n916), .C1(new_n917), .C2(new_n302), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n919), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n915), .A2(new_n924), .A3(KEYINPUT40), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n911), .A2(KEYINPUT38), .A3(new_n912), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT106), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n891), .A2(new_n899), .B1(new_n403), .B2(new_n901), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n926), .B(new_n927), .C1(new_n928), .C2(KEYINPUT38), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n914), .A2(new_n925), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT38), .B1(new_n911), .B2(new_n912), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n924), .B(new_n915), .C1(new_n913), .C2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT40), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(G330), .B1(new_n884), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(new_n935), .B2(new_n884), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n469), .B1(new_n722), .B2(new_n731), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n660), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT39), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n903), .B2(new_n913), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n326), .A2(new_n697), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n911), .A2(new_n912), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT38), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n946), .A2(KEYINPUT39), .A3(new_n926), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n942), .A2(new_n943), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n697), .B1(new_n820), .B2(new_n822), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n825), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n946), .A2(new_n926), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n951), .A2(new_n952), .A3(new_n924), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n651), .A2(new_n695), .ZN(new_n954));
  AND3_X1   g0754(.A1(new_n948), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n940), .B(new_n955), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n937), .A2(new_n956), .B1(new_n203), .B2(new_n753), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n937), .A2(new_n956), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n876), .B1(new_n957), .B2(new_n958), .ZN(G367));
  OAI21_X1  g0759(.A(new_n686), .B1(new_n632), .B2(new_n704), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n674), .A2(new_n697), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n711), .A2(new_n963), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n964), .A2(KEYINPUT42), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n960), .A2(new_n566), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n697), .B1(new_n966), .B2(new_n624), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(new_n964), .B2(KEYINPUT42), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n666), .B1(new_n598), .B2(new_n704), .ZN(new_n969));
  OR3_X1    g0769(.A1(new_n665), .A2(new_n598), .A3(new_n704), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n965), .A2(new_n968), .B1(KEYINPUT43), .B2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n971), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT43), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n708), .A2(new_n963), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n965), .A2(new_n968), .A3(new_n974), .A4(new_n973), .ZN(new_n978));
  AND3_X1   g0778(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n977), .B1(new_n976), .B2(new_n978), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n714), .B(KEYINPUT41), .Z(new_n982));
  NAND3_X1  g0782(.A1(new_n711), .A2(new_n709), .A3(new_n962), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT45), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n983), .B(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n711), .A2(new_n709), .ZN(new_n986));
  AOI21_X1  g0786(.A(KEYINPUT44), .B1(new_n986), .B2(new_n963), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n963), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT44), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n985), .B1(new_n987), .B2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n708), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n710), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n711), .B1(new_n707), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(new_n703), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n751), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n985), .B(new_n708), .C1(new_n987), .C2(new_n990), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n993), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n982), .B1(new_n1000), .B2(new_n751), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n981), .B1(new_n1001), .B2(new_n755), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(KEYINPUT108), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT108), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n981), .B(new_n1004), .C1(new_n1001), .C2(new_n755), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n772), .B1(new_n207), .B2(new_n448), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n767), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1008), .A2(new_n233), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n756), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT109), .Z(new_n1011));
  INV_X1    g0811(.A(new_n770), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n786), .A2(G311), .B1(G107), .B2(new_n797), .ZN(new_n1013));
  INV_X1    g0813(.A(G294), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1013), .B1(new_n267), .B2(new_n794), .C1(new_n1014), .C2(new_n804), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n807), .A2(G303), .B1(new_n783), .B2(G317), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT46), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n791), .B2(new_n492), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n792), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n290), .B1(new_n847), .B2(G283), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1016), .A2(new_n1018), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n795), .A2(G77), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n797), .A2(G68), .ZN(new_n1023));
  INV_X1    g0823(.A(G58), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1022), .B(new_n1023), .C1(new_n1024), .C2(new_n791), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n802), .A2(new_n789), .B1(new_n786), .B2(G143), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n266), .B1(new_n807), .B2(G150), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G50), .A2(new_n847), .B1(new_n783), .B2(G137), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n1015), .A2(new_n1021), .B1(new_n1025), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT47), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1012), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n1031), .B2(new_n1030), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1011), .A2(new_n1033), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT110), .Z(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n761), .B2(new_n971), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1006), .A2(new_n1036), .ZN(G387));
  NAND2_X1  g0837(.A1(new_n996), .A2(new_n755), .ZN(new_n1038));
  AND2_X1   g0838(.A1(new_n1038), .A2(KEYINPUT111), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1038), .A2(KEYINPUT111), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n996), .A2(new_n751), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1042), .A2(new_n714), .A3(new_n997), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n807), .A2(G317), .B1(new_n847), .B2(G303), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n786), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1044), .B1(new_n804), .B2(new_n779), .C1(new_n775), .C2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT48), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n792), .A2(G294), .B1(new_n797), .B2(G283), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1052), .A2(KEYINPUT49), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(KEYINPUT49), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n794), .A2(new_n492), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n290), .B(new_n1055), .C1(new_n783), .C2(new_n787), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1053), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n778), .A2(new_n408), .B1(new_n782), .B2(new_n405), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n266), .B(new_n1058), .C1(G50), .C2(new_n807), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n792), .A2(G77), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n789), .A2(new_n362), .B1(new_n580), .B2(new_n797), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n786), .A2(G159), .B1(new_n795), .B2(G97), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1012), .B1(new_n1057), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n230), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT112), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n362), .A2(new_n315), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT50), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n716), .B(new_n252), .C1(new_n408), .C2(new_n317), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n767), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n1065), .A2(G45), .B1(new_n1066), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n1066), .B2(new_n1070), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(G107), .B2(new_n207), .C1(new_n716), .C2(new_n763), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n757), .B(new_n1064), .C1(new_n772), .C2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n707), .B2(new_n761), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1041), .A2(new_n1043), .A3(new_n1075), .ZN(G393));
  NAND2_X1  g0876(.A1(new_n1000), .A2(new_n714), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n999), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n988), .B(new_n989), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n708), .B1(new_n1079), .B2(new_n985), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(KEYINPUT115), .B1(new_n1081), .B2(new_n998), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT115), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n997), .B(new_n1083), .C1(new_n1078), .C2(new_n1080), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1077), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1081), .A2(new_n755), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n772), .B1(new_n267), .B2(new_n207), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1008), .A2(new_n241), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n756), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n789), .A2(G50), .B1(new_n847), .B2(new_n362), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n1090), .A2(KEYINPUT113), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(KEYINPUT113), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n266), .B(new_n843), .C1(G143), .C2(new_n783), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n792), .A2(new_n214), .B1(new_n797), .B2(G77), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(G150), .A2(new_n786), .B1(new_n807), .B2(G159), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT51), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(G317), .A2(new_n786), .B1(new_n807), .B2(G311), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT52), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n266), .B1(new_n782), .B2(new_n775), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(G294), .B2(new_n847), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n789), .A2(G303), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n792), .A2(G283), .B1(new_n797), .B2(G116), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1101), .A2(new_n809), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n1095), .A2(new_n1097), .B1(new_n1099), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1089), .B1(new_n1105), .B2(new_n770), .ZN(new_n1106));
  XOR2_X1   g0906(.A(new_n1106), .B(KEYINPUT114), .Z(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n962), .B2(new_n761), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1086), .A2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1085), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(G390));
  NAND2_X1  g0911(.A1(new_n942), .A2(new_n947), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n943), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n949), .B1(new_n688), .B2(new_n824), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n924), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1112), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n915), .A2(new_n924), .A3(G330), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n729), .A2(new_n704), .A3(new_n823), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n950), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n943), .B1(new_n1120), .B2(new_n924), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1121), .A2(new_n914), .A3(new_n929), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n1117), .A2(new_n1118), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1118), .B1(new_n1117), .B2(new_n1122), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1112), .A2(new_n758), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n841), .A2(new_n362), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n266), .B1(new_n783), .B2(G125), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n853), .B2(new_n774), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(KEYINPUT54), .B(G143), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT118), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1129), .B1(new_n1132), .B2(new_n847), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n791), .A2(new_n405), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT53), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n789), .A2(G137), .B1(G159), .B2(new_n797), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n786), .A2(G128), .B1(new_n795), .B2(G50), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1133), .A2(new_n1135), .A3(new_n1136), .A4(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT119), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n786), .A2(G283), .B1(G77), .B2(new_n797), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1140), .A2(new_n800), .A3(new_n852), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n266), .B1(new_n782), .B2(new_n1014), .C1(new_n774), .C2(new_n492), .ZN(new_n1142));
  OR2_X1    g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n789), .A2(G107), .B1(new_n847), .B2(G97), .ZN(new_n1144));
  XOR2_X1   g0944(.A(new_n1144), .B(KEYINPUT120), .Z(new_n1145));
  OAI21_X1  g0945(.A(new_n1139), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1146), .A2(KEYINPUT121), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1012), .B1(new_n1146), .B2(KEYINPUT121), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n757), .B(new_n1127), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n1125), .A2(new_n755), .B1(new_n1126), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1117), .A2(new_n1122), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1118), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1117), .A2(new_n1118), .A3(new_n1122), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n469), .A2(new_n749), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1157), .B(new_n938), .C1(new_n655), .C2(new_n659), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1153), .A2(new_n1120), .ZN(new_n1159));
  INV_X1    g0959(.A(G330), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n879), .B2(new_n881), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT116), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n831), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n749), .A2(KEYINPUT116), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1115), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1159), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n882), .A2(G330), .A3(new_n831), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n1115), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n1118), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n951), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1166), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT117), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1158), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1157), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n643), .A2(KEYINPUT90), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n652), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n639), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n656), .B1(new_n1178), .B2(new_n466), .ZN(new_n1179));
  AOI211_X1 g0979(.A(KEYINPUT92), .B(new_n654), .C1(new_n1177), .C2(new_n639), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n939), .B(new_n1174), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1159), .A2(new_n1165), .B1(new_n1169), .B2(new_n951), .ZN(new_n1182));
  OAI21_X1  g0982(.A(KEYINPUT117), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n1156), .A2(new_n1173), .A3(new_n1183), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1154), .A2(new_n1155), .A3(new_n1158), .A4(new_n1171), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n714), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1151), .B1(new_n1184), .B2(new_n1186), .ZN(G378));
  XNOR2_X1  g0987(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n639), .A2(new_n466), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n414), .A2(new_n695), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1189), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  OR2_X1    g0995(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1196), .A2(new_n1192), .A3(new_n1188), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n758), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n756), .B1(G50), .B2(new_n841), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1023), .B1(new_n1045), .B2(new_n492), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT123), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n794), .A2(new_n1024), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT122), .Z(new_n1204));
  NAND2_X1  g1004(.A1(new_n266), .A2(new_n250), .ZN(new_n1205));
  INV_X1    g1005(.A(G283), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n778), .A2(new_n448), .B1(new_n782), .B2(new_n1206), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1205), .B(new_n1207), .C1(G107), .C2(new_n807), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n789), .A2(G97), .B1(new_n792), .B2(G77), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1202), .A2(new_n1204), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT58), .ZN(new_n1211));
  AOI21_X1  g1011(.A(G50), .B1(new_n249), .B2(new_n250), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1210), .A2(new_n1211), .B1(new_n1205), .B2(new_n1212), .ZN(new_n1213));
  AOI211_X1 g1013(.A(G33), .B(G41), .C1(new_n783), .C2(G124), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n786), .A2(G125), .B1(new_n847), .B2(G137), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n789), .A2(G132), .B1(G150), .B2(new_n797), .ZN(new_n1216));
  INV_X1    g1016(.A(G128), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n1131), .A2(new_n791), .B1(new_n1217), .B2(new_n774), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT124), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1215), .B(new_n1216), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT125), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT59), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1214), .B1(new_n801), .B2(new_n794), .C1(new_n1223), .C2(new_n1224), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1213), .B1(new_n1211), .B2(new_n1210), .C1(new_n1225), .C2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1200), .B1(new_n1227), .B2(new_n770), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1199), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT126), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1199), .A2(KEYINPUT126), .A3(new_n1228), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n948), .A2(new_n953), .A3(new_n954), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1160), .B1(new_n932), .B2(new_n933), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1236));
  AND3_X1   g1036(.A1(new_n1235), .A2(new_n1236), .A3(new_n930), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1236), .B1(new_n1235), .B2(new_n930), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1234), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1235), .A2(new_n930), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n1198), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1235), .A2(new_n1236), .A3(new_n930), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1241), .A2(new_n955), .A3(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1239), .A2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1233), .B1(new_n1244), .B2(new_n755), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(new_n1237), .A2(new_n1238), .A3(new_n1234), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n955), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1247));
  OAI21_X1  g1047(.A(KEYINPUT57), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1181), .B1(new_n1125), .B2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n714), .B1(new_n1248), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1185), .A2(new_n1158), .ZN(new_n1252));
  AOI21_X1  g1052(.A(KEYINPUT57), .B1(new_n1252), .B2(new_n1244), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1245), .B1(new_n1251), .B2(new_n1253), .ZN(G375));
  INV_X1    g1054(.A(new_n982), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1173), .A2(new_n1183), .A3(new_n1255), .A4(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1115), .A2(new_n758), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n756), .B1(G68), .B2(new_n841), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n804), .A2(new_n492), .B1(new_n1045), .B2(new_n1014), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(G97), .B2(new_n792), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n580), .A2(new_n797), .ZN(new_n1262));
  INV_X1    g1062(.A(G303), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n778), .A2(new_n518), .B1(new_n782), .B2(new_n1263), .ZN(new_n1264));
  AOI211_X1 g1064(.A(new_n290), .B(new_n1264), .C1(G283), .C2(new_n807), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1261), .A2(new_n1022), .A3(new_n1262), .A4(new_n1265), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n1045), .A2(new_n853), .B1(new_n791), .B2(new_n335), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(G50), .B2(new_n797), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n778), .A2(new_n405), .B1(new_n782), .B2(new_n1217), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n266), .B(new_n1269), .C1(G137), .C2(new_n807), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1268), .B(new_n1270), .C1(new_n804), .C2(new_n1131), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1204), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1266), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1259), .B1(new_n1273), .B2(new_n770), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n1171), .A2(new_n755), .B1(new_n1258), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1257), .A2(new_n1275), .ZN(G381));
  INV_X1    g1076(.A(G396), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1041), .A2(new_n1277), .A3(new_n1043), .A4(new_n1075), .ZN(new_n1278));
  NOR4_X1   g1078(.A1(G390), .A2(G384), .A3(G381), .A4(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1126), .A2(new_n1150), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n1156), .B2(new_n754), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1156), .A2(new_n1173), .A3(new_n1183), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n715), .B1(new_n1125), .B2(new_n1249), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1281), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1279), .A2(new_n1006), .A3(new_n1036), .A4(new_n1284), .ZN(new_n1285));
  OR2_X1    g1085(.A1(new_n1285), .A2(G375), .ZN(G407));
  NAND2_X1  g1086(.A1(new_n696), .A2(G213), .ZN(new_n1287));
  OR3_X1    g1087(.A1(G375), .A2(G378), .A3(new_n1287), .ZN(new_n1288));
  OAI211_X1 g1088(.A(G213), .B(new_n1288), .C1(new_n1285), .C2(G375), .ZN(G409));
  OAI21_X1  g1089(.A(new_n1075), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1043), .ZN(new_n1291));
  OAI21_X1  g1091(.A(G396), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1278), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1109), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1293), .B(new_n1294), .C1(new_n1295), .C2(new_n1077), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n1278), .B(new_n1292), .C1(new_n1085), .C2(new_n1109), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(G387), .A2(new_n1298), .ZN(new_n1299));
  AOI22_X1  g1099(.A1(new_n1006), .A2(new_n1036), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  OAI211_X1 g1101(.A(G378), .B(new_n1245), .C1(new_n1251), .C2(new_n1253), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1252), .A2(new_n1255), .A3(new_n1244), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1245), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1284), .ZN(new_n1305));
  AOI22_X1  g1105(.A1(new_n1302), .A2(new_n1305), .B1(G213), .B2(new_n696), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1181), .A2(KEYINPUT60), .A3(new_n1182), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n714), .ZN(new_n1308));
  OAI21_X1  g1108(.A(KEYINPUT60), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1308), .B1(new_n1256), .B2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1275), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n864), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1308), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1309), .A2(new_n1256), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1315), .A2(G384), .A3(new_n1275), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1312), .A2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1306), .A2(KEYINPUT63), .A3(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1302), .A2(new_n1305), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1320), .A2(new_n1287), .A3(new_n1318), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT63), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1320), .A2(new_n1287), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n696), .A2(G213), .A3(G2897), .ZN(new_n1325));
  AND3_X1   g1125(.A1(new_n1312), .A2(new_n1316), .A3(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1325), .B1(new_n1312), .B2(new_n1316), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(KEYINPUT61), .B1(new_n1324), .B2(new_n1328), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1301), .A2(new_n1319), .A3(new_n1323), .A4(new_n1329), .ZN(new_n1330));
  AND4_X1   g1130(.A1(KEYINPUT62), .A2(new_n1320), .A3(new_n1287), .A4(new_n1318), .ZN(new_n1331));
  AOI21_X1  g1131(.A(KEYINPUT62), .B1(new_n1306), .B2(new_n1318), .ZN(new_n1332));
  OAI211_X1 g1132(.A(new_n1329), .B(KEYINPUT127), .C1(new_n1331), .C2(new_n1332), .ZN(new_n1333));
  XNOR2_X1  g1133(.A(G387), .B(new_n1298), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT62), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1321), .A2(new_n1336), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1306), .A2(KEYINPUT62), .A3(new_n1318), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(KEYINPUT127), .B1(new_n1339), .B2(new_n1329), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1330), .B1(new_n1335), .B2(new_n1340), .ZN(G405));
  NAND2_X1  g1141(.A1(G375), .A2(new_n1284), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(new_n1302), .ZN(new_n1343));
  XNOR2_X1  g1143(.A(new_n1343), .B(new_n1317), .ZN(new_n1344));
  XNOR2_X1  g1144(.A(new_n1301), .B(new_n1344), .ZN(G402));
endmodule


