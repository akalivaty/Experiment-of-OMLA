//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 0 0 1 0 0 0 1 1 0 0 1 0 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1280, new_n1281, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(KEYINPUT64), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n208), .B(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n211));
  INV_X1    g0011(.A(G50), .ZN(new_n212));
  INV_X1    g0012(.A(G226), .ZN(new_n213));
  INV_X1    g0013(.A(G97), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n217), .B1(new_n202), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n210), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  OR2_X1    g0023(.A1(new_n203), .A2(KEYINPUT65), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n203), .A2(KEYINPUT65), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n224), .A2(G50), .A3(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n228), .A2(new_n207), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n210), .A2(G13), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(G264), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n220), .B(new_n232), .C1(new_n215), .C2(new_n233), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n230), .B1(new_n234), .B2(KEYINPUT0), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n223), .B(new_n235), .C1(KEYINPUT0), .C2(new_n234), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G250), .B(G257), .Z(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  NOR2_X1   g0051(.A1(new_n207), .A2(G1), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(KEYINPUT66), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n254), .A2(new_n228), .A3(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G50), .ZN(new_n260));
  OAI21_X1  g0060(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n261));
  INV_X1    g0061(.A(G150), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G20), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT8), .B(G58), .ZN(new_n268));
  OAI221_X1 g0068(.A(new_n261), .B1(new_n262), .B2(new_n264), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n255), .A2(new_n228), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n254), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n212), .ZN(new_n273));
  AND3_X1   g0073(.A1(new_n260), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT9), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n260), .A2(new_n271), .A3(new_n273), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT9), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AND2_X1   g0078(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT67), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(KEYINPUT10), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT3), .B(G33), .ZN(new_n283));
  INV_X1    g0083(.A(G1698), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(G222), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G77), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n283), .A2(G1698), .ZN(new_n287));
  INV_X1    g0087(.A(G223), .ZN(new_n288));
  OAI221_X1 g0088(.A(new_n285), .B1(new_n286), .B2(new_n283), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G41), .ZN(new_n290));
  OAI211_X1 g0090(.A(G1), .B(G13), .C1(new_n265), .C2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n294));
  INV_X1    g0094(.A(G274), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n291), .A2(new_n294), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n297), .B1(new_n299), .B2(G226), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n293), .A2(new_n300), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n301), .A2(G200), .B1(new_n280), .B2(KEYINPUT10), .ZN(new_n302));
  INV_X1    g0102(.A(new_n301), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G190), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n279), .A2(new_n282), .A3(new_n302), .A4(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT10), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n275), .A2(new_n304), .A3(new_n278), .ZN(new_n307));
  INV_X1    g0107(.A(G200), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  OAI211_X1 g0109(.A(KEYINPUT67), .B(new_n306), .C1(new_n307), .C2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G169), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n274), .B1(new_n311), .B2(new_n301), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(G179), .B2(new_n301), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n305), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n296), .B1(new_n298), .B2(new_n218), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT68), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n316), .B(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT13), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n283), .A2(G232), .A3(G1698), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n283), .A2(G226), .A3(new_n284), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G33), .A2(G97), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n292), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n318), .A2(new_n319), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n319), .B1(new_n318), .B2(new_n324), .ZN(new_n326));
  OAI21_X1  g0126(.A(G200), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n318), .A2(new_n324), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT13), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n318), .A2(new_n319), .A3(new_n324), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n329), .A2(G190), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n270), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n266), .A2(G77), .B1(G20), .B2(new_n202), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n263), .A2(G50), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  XOR2_X1   g0135(.A(new_n335), .B(KEYINPUT11), .Z(new_n336));
  NAND2_X1  g0136(.A1(new_n272), .A2(new_n202), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n337), .B(KEYINPUT12), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n259), .A2(G68), .ZN(new_n339));
  AND3_X1   g0139(.A1(new_n336), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  AND3_X1   g0140(.A1(new_n327), .A2(new_n331), .A3(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(G169), .B1(new_n325), .B2(new_n326), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT14), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT14), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n344), .B(G169), .C1(new_n325), .C2(new_n326), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n325), .A2(new_n326), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G179), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n343), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n340), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n341), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n272), .A2(new_n286), .ZN(new_n351));
  INV_X1    g0151(.A(new_n268), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n352), .A2(new_n263), .B1(G20), .B2(G77), .ZN(new_n353));
  XNOR2_X1  g0153(.A(KEYINPUT15), .B(G87), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n266), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  OAI221_X1 g0157(.A(new_n351), .B1(new_n286), .B2(new_n258), .C1(new_n357), .C2(new_n332), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n299), .A2(G244), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n283), .A2(G232), .A3(new_n284), .ZN(new_n360));
  INV_X1    g0160(.A(G107), .ZN(new_n361));
  OAI221_X1 g0161(.A(new_n360), .B1(new_n361), .B2(new_n283), .C1(new_n287), .C2(new_n218), .ZN(new_n362));
  AOI211_X1 g0162(.A(new_n297), .B(new_n359), .C1(new_n292), .C2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n358), .B1(G190), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n308), .B2(new_n363), .ZN(new_n365));
  INV_X1    g0165(.A(G179), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n358), .B1(new_n363), .B2(G169), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n315), .A2(new_n350), .A3(new_n365), .A4(new_n370), .ZN(new_n371));
  AND2_X1   g0171(.A1(KEYINPUT70), .A2(KEYINPUT3), .ZN(new_n372));
  NOR2_X1   g0172(.A1(KEYINPUT70), .A2(KEYINPUT3), .ZN(new_n373));
  OAI21_X1  g0173(.A(G33), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  XNOR2_X1  g0174(.A(KEYINPUT69), .B(G33), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT3), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n233), .A2(G1698), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(G257), .B2(G1698), .ZN(new_n379));
  INV_X1    g0179(.A(G303), .ZN(new_n380));
  OAI22_X1  g0180(.A1(new_n377), .A2(new_n379), .B1(new_n380), .B2(new_n283), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT82), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT82), .ZN(new_n383));
  OAI221_X1 g0183(.A(new_n383), .B1(new_n380), .B2(new_n283), .C1(new_n377), .C2(new_n379), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n382), .A2(new_n384), .A3(new_n292), .ZN(new_n385));
  INV_X1    g0185(.A(G45), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n386), .A2(G1), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n290), .A2(KEYINPUT5), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT5), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G41), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n387), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n391), .A2(new_n295), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n391), .A2(new_n291), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n392), .B1(new_n393), .B2(G270), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n385), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT76), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n265), .B2(G1), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n206), .A2(KEYINPUT76), .A3(G33), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n256), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(G116), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT78), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT78), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(G116), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n400), .A2(G116), .B1(new_n405), .B2(new_n272), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT83), .ZN(new_n407));
  XNOR2_X1  g0207(.A(KEYINPUT78), .B(G116), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n270), .B1(new_n408), .B2(new_n207), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G33), .A2(G283), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n207), .ZN(new_n411));
  XNOR2_X1  g0211(.A(KEYINPUT75), .B(G97), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n411), .B1(new_n412), .B2(new_n265), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n407), .B1(new_n414), .B2(KEYINPUT20), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n214), .A2(KEYINPUT75), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT75), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(G97), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n207), .B(new_n410), .C1(new_n419), .C2(G33), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n405), .A2(G20), .B1(new_n228), .B2(new_n255), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n420), .A2(new_n421), .A3(new_n407), .A4(KEYINPUT20), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT20), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(new_n409), .B2(new_n413), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n406), .B1(new_n415), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n395), .A2(G169), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT21), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n395), .A2(KEYINPUT21), .A3(new_n426), .A4(G169), .ZN(new_n430));
  INV_X1    g0230(.A(new_n426), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n385), .A2(G190), .A3(new_n394), .ZN(new_n432));
  INV_X1    g0232(.A(new_n394), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n291), .B1(new_n381), .B2(KEYINPUT82), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n433), .B1(new_n434), .B2(new_n384), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n431), .B(new_n432), .C1(new_n308), .C2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(new_n426), .A3(G179), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n429), .A2(new_n430), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n375), .A2(G294), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n220), .A2(new_n284), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n215), .A2(G1698), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n440), .B1(new_n377), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n391), .A2(G264), .A3(new_n291), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT88), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n391), .A2(KEYINPUT88), .A3(G264), .A4(new_n291), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n444), .A2(new_n292), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n392), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(G169), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n449), .A2(G179), .A3(new_n450), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n452), .A2(KEYINPUT89), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT89), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n444), .A2(new_n292), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n447), .A2(new_n448), .ZN(new_n457));
  AND4_X1   g0257(.A1(G179), .A2(new_n456), .A3(new_n450), .A4(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n311), .B1(new_n449), .B2(new_n450), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n455), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n454), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT69), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(G33), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n265), .A2(KEYINPUT69), .ZN(new_n464));
  OAI21_X1  g0264(.A(KEYINPUT3), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n219), .A2(G20), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n465), .A2(new_n374), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT84), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT84), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n465), .A2(new_n469), .A3(new_n374), .A4(new_n466), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n468), .A2(KEYINPUT22), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT22), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n283), .A2(new_n472), .A3(new_n466), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT86), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n265), .A2(KEYINPUT69), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n462), .A2(G33), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n402), .A2(new_n404), .A3(new_n476), .A4(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n475), .B1(new_n478), .B2(G20), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n408), .A2(new_n375), .A3(KEYINPUT86), .A4(new_n207), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT87), .B1(new_n361), .B2(G20), .ZN(new_n482));
  XOR2_X1   g0282(.A(new_n482), .B(KEYINPUT23), .Z(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  XNOR2_X1  g0285(.A(KEYINPUT85), .B(KEYINPUT24), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n474), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n473), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n472), .B1(new_n467), .B2(KEYINPUT84), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n489), .B1(new_n490), .B2(new_n470), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n486), .B1(new_n491), .B2(new_n484), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n488), .A2(new_n492), .A3(new_n270), .ZN(new_n493));
  INV_X1    g0293(.A(new_n400), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n494), .A2(new_n361), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n272), .A2(new_n361), .ZN(new_n496));
  XNOR2_X1  g0296(.A(new_n496), .B(KEYINPUT25), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n461), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n449), .A2(G190), .A3(new_n450), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n451), .A2(G200), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n493), .A2(new_n498), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n478), .ZN(new_n504));
  OR2_X1    g0304(.A1(KEYINPUT70), .A2(KEYINPUT3), .ZN(new_n505));
  NAND2_X1  g0305(.A1(KEYINPUT70), .A2(KEYINPUT3), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n265), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n376), .B1(new_n476), .B2(new_n477), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n218), .A2(G1698), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n504), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n465), .A2(G244), .A3(G1698), .A4(new_n374), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n291), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n291), .B(G250), .C1(G1), .C2(new_n386), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n387), .A2(G274), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(G200), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n355), .A2(new_n254), .ZN(new_n518));
  NOR3_X1   g0318(.A1(new_n256), .A2(new_n399), .A3(new_n219), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n219), .A2(KEYINPUT80), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT80), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G87), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n419), .A2(new_n523), .A3(new_n361), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT19), .ZN(new_n525));
  OAI211_X1 g0325(.A(KEYINPUT79), .B(new_n207), .C1(new_n322), .C2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n207), .B1(new_n322), .B2(new_n525), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT79), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n524), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n202), .A2(G20), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n374), .B(new_n531), .C1(new_n376), .C2(new_n375), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n525), .B1(new_n419), .B2(new_n267), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n530), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AOI211_X1 g0334(.A(new_n518), .B(new_n519), .C1(new_n534), .C2(new_n270), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n465), .A2(new_n374), .A3(new_n510), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n512), .A2(new_n478), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n516), .B1(new_n537), .B2(new_n292), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G190), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n517), .A2(new_n535), .A3(new_n539), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n524), .A2(new_n526), .A3(new_n529), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n532), .A2(new_n533), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n270), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(KEYINPUT81), .B1(new_n400), .B2(new_n355), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT81), .ZN(new_n545));
  NOR4_X1   g0345(.A1(new_n256), .A2(new_n399), .A3(new_n545), .A4(new_n354), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n518), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n543), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n537), .A2(new_n292), .ZN(new_n550));
  INV_X1    g0350(.A(new_n516), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n550), .A2(new_n366), .A3(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n549), .B(new_n552), .C1(G169), .C2(new_n538), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n540), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT7), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n555), .A2(G20), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n505), .A2(new_n265), .A3(new_n506), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n476), .A2(new_n477), .A3(new_n376), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AND2_X1   g0360(.A1(KEYINPUT3), .A2(G33), .ZN(new_n561));
  NOR2_X1   g0361(.A1(KEYINPUT3), .A2(G33), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(KEYINPUT7), .B1(new_n563), .B2(new_n207), .ZN(new_n564));
  OAI21_X1  g0364(.A(G107), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT6), .ZN(new_n566));
  AND2_X1   g0366(.A1(G97), .A2(G107), .ZN(new_n567));
  NOR2_X1   g0367(.A1(G97), .A2(G107), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n361), .A2(KEYINPUT6), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n569), .B1(new_n419), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n571), .A2(G20), .B1(G77), .B2(new_n263), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n565), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n270), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n254), .A2(G97), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n575), .B1(new_n400), .B2(G97), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(KEYINPUT77), .A3(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT77), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n332), .B1(new_n565), .B2(new_n572), .ZN(new_n579));
  INV_X1    g0379(.A(new_n576), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n392), .B1(new_n393), .B2(G257), .ZN(new_n582));
  AND2_X1   g0382(.A1(KEYINPUT4), .A2(G244), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n284), .B(new_n583), .C1(new_n561), .C2(new_n562), .ZN(new_n584));
  OAI211_X1 g0384(.A(G250), .B(G1698), .C1(new_n561), .C2(new_n562), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n584), .A2(new_n585), .A3(new_n410), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n465), .A2(G244), .A3(new_n284), .A4(new_n374), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT4), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n582), .B1(new_n589), .B2(new_n291), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G169), .ZN(new_n591));
  OAI211_X1 g0391(.A(G179), .B(new_n582), .C1(new_n589), .C2(new_n291), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n577), .A2(new_n581), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n590), .A2(G200), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n580), .B1(new_n573), .B2(new_n270), .ZN(new_n595));
  OAI211_X1 g0395(.A(G190), .B(new_n582), .C1(new_n589), .C2(new_n291), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n554), .A2(new_n593), .A3(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n439), .A2(new_n500), .A3(new_n503), .A4(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(G159), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n264), .A2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(G58), .A2(G68), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n207), .B1(new_n203), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT71), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n602), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(KEYINPUT71), .B1(new_n601), .B2(new_n604), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(G20), .B1(new_n465), .B2(new_n374), .ZN(new_n610));
  OAI21_X1  g0410(.A(G68), .B1(new_n610), .B2(new_n555), .ZN(new_n611));
  AOI211_X1 g0411(.A(KEYINPUT7), .B(G20), .C1(new_n465), .C2(new_n374), .ZN(new_n612));
  OAI211_X1 g0412(.A(KEYINPUT16), .B(new_n609), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT16), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n476), .A2(new_n477), .A3(new_n376), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n372), .A2(new_n373), .A3(G33), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n556), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n555), .B1(new_n283), .B2(G20), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n202), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n602), .A2(new_n605), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n614), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n613), .A2(new_n270), .A3(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(G223), .A2(G1698), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n623), .B1(new_n213), .B2(G1698), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n624), .B(new_n374), .C1(new_n376), .C2(new_n375), .ZN(new_n625));
  NAND2_X1  g0425(.A1(G33), .A2(G87), .ZN(new_n626));
  XNOR2_X1  g0426(.A(new_n626), .B(KEYINPUT72), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n292), .ZN(new_n629));
  INV_X1    g0429(.A(G232), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n296), .B1(new_n298), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n308), .B1(new_n629), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n291), .B1(new_n625), .B2(new_n627), .ZN(new_n634));
  INV_X1    g0434(.A(G190), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n634), .A2(new_n635), .A3(new_n631), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n268), .A2(new_n254), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(new_n259), .B2(new_n268), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n622), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(KEYINPUT74), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT74), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n622), .A2(new_n637), .A3(new_n642), .A4(new_n639), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n641), .A2(KEYINPUT17), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n622), .A2(new_n639), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT73), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n629), .A2(new_n366), .A3(new_n632), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n311), .B1(new_n634), .B2(new_n631), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n647), .A2(new_n646), .A3(new_n648), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n645), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(KEYINPUT18), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT18), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n645), .A2(new_n654), .A3(new_n650), .A4(new_n651), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT17), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n640), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n644), .A2(new_n653), .A3(new_n655), .A4(new_n657), .ZN(new_n658));
  NOR3_X1   g0458(.A1(new_n371), .A2(new_n599), .A3(new_n658), .ZN(G372));
  NAND2_X1  g0459(.A1(new_n653), .A2(new_n655), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n342), .A2(KEYINPUT14), .B1(new_n346), .B2(G179), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n340), .B1(new_n661), .B2(new_n345), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n341), .B1(new_n663), .B2(new_n370), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n644), .A2(new_n657), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n660), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n305), .A2(new_n310), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n313), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n595), .B1(new_n591), .B2(new_n592), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT26), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n671), .A2(new_n540), .A3(new_n553), .A4(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n577), .A2(new_n581), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n591), .A2(new_n592), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n554), .A2(new_n676), .ZN(new_n677));
  OAI211_X1 g0477(.A(new_n553), .B(new_n673), .C1(new_n677), .C2(new_n672), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n593), .A2(new_n597), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n540), .A2(new_n553), .ZN(new_n680));
  AND3_X1   g0480(.A1(new_n679), .A2(new_n503), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT90), .ZN(new_n682));
  INV_X1    g0482(.A(new_n498), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n484), .B1(new_n471), .B2(new_n473), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n332), .B1(new_n684), .B2(new_n487), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n683), .B1(new_n685), .B2(new_n492), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n458), .A2(new_n459), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n682), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n687), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n499), .A2(KEYINPUT90), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n430), .A2(new_n437), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n311), .B1(new_n385), .B2(new_n394), .ZN(new_n692));
  AOI21_X1  g0492(.A(KEYINPUT21), .B1(new_n692), .B2(new_n426), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n688), .A2(new_n690), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n678), .B1(new_n681), .B2(new_n695), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n371), .A2(new_n696), .A3(new_n658), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n670), .A2(new_n697), .ZN(G369));
  NAND3_X1  g0498(.A1(new_n429), .A2(new_n430), .A3(new_n437), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n207), .A2(G13), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n206), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n701), .A2(KEYINPUT27), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(KEYINPUT27), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G213), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(G343), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n431), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n699), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n438), .B2(new_n708), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(G330), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n499), .B1(new_n461), .B2(new_n706), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n454), .A2(new_n460), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(new_n686), .ZN(new_n716));
  AOI22_X1  g0516(.A1(new_n714), .A2(new_n503), .B1(new_n716), .B2(new_n706), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n699), .A2(new_n707), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n713), .A2(new_n719), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n688), .A2(new_n690), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n706), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n714), .A2(new_n503), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n718), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n720), .A2(new_n723), .A3(new_n726), .ZN(G399));
  NOR2_X1   g0527(.A1(new_n232), .A2(G41), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G1), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n524), .A2(G116), .ZN(new_n731));
  OAI22_X1  g0531(.A1(new_n730), .A2(new_n731), .B1(new_n226), .B2(new_n729), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(KEYINPUT28), .ZN(new_n733));
  OAI211_X1 g0533(.A(new_n598), .B(new_n503), .C1(new_n716), .C2(new_n699), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n671), .A2(new_n540), .A3(new_n553), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(KEYINPUT26), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n593), .A2(new_n672), .A3(new_n553), .A4(new_n540), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n736), .A2(new_n553), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n706), .B1(new_n734), .B2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT29), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT91), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT30), .ZN(new_n743));
  OR2_X1    g0543(.A1(new_n589), .A2(new_n291), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n744), .A2(new_n449), .A3(new_n538), .A4(new_n582), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n385), .A2(G179), .A3(new_n394), .ZN(new_n746));
  OAI211_X1 g0546(.A(new_n742), .B(new_n743), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n538), .A2(G179), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n395), .A2(new_n748), .A3(new_n451), .A4(new_n590), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n538), .A2(new_n449), .ZN(new_n751));
  INV_X1    g0551(.A(new_n590), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n751), .A2(new_n435), .A3(G179), .A4(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n743), .B1(new_n753), .B2(new_n742), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n706), .B1(new_n750), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT31), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI211_X1 g0557(.A(KEYINPUT31), .B(new_n706), .C1(new_n750), .C2(new_n754), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n757), .B(new_n758), .C1(new_n599), .C2(new_n706), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G330), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n695), .A2(new_n681), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n673), .A2(new_n553), .ZN(new_n762));
  INV_X1    g0562(.A(new_n677), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n762), .B1(new_n763), .B2(KEYINPUT26), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n706), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(new_n740), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n741), .A2(new_n760), .A3(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n733), .B1(new_n768), .B2(G1), .ZN(G364));
  AOI21_X1  g0569(.A(new_n206), .B1(new_n700), .B2(G45), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n728), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n713), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n773), .B1(G330), .B2(new_n710), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n772), .B(KEYINPUT92), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n231), .A2(G355), .A3(new_n283), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(G116), .B2(new_n231), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n232), .A2(new_n509), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n780), .B1(new_n386), .B2(new_n227), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n247), .A2(new_n386), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n778), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G13), .A2(G33), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G20), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n228), .B1(G20), .B2(new_n311), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n776), .B1(new_n783), .B2(new_n789), .ZN(new_n790));
  XOR2_X1   g0590(.A(KEYINPUT33), .B(G317), .Z(new_n791));
  NOR2_X1   g0591(.A1(new_n366), .A2(new_n308), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n207), .A2(G190), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n207), .A2(new_n635), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n308), .A2(G179), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n791), .A2(new_n794), .B1(new_n797), .B2(new_n380), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n793), .A2(new_n796), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n283), .B(new_n798), .C1(G283), .C2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n795), .A2(new_n792), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(G179), .A2(G200), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n793), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n803), .A2(G326), .B1(new_n806), .B2(G329), .ZN(new_n807));
  INV_X1    g0607(.A(new_n795), .ZN(new_n808));
  NOR3_X1   g0608(.A1(new_n808), .A2(new_n366), .A3(G200), .ZN(new_n809));
  INV_X1    g0609(.A(new_n793), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n810), .A2(new_n366), .A3(G200), .ZN(new_n811));
  AOI22_X1  g0611(.A1(G322), .A2(new_n809), .B1(new_n811), .B2(G311), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n207), .B1(new_n804), .B2(G190), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G294), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n801), .A2(new_n807), .A3(new_n812), .A4(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n809), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n817), .A2(new_n201), .B1(new_n802), .B2(new_n212), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(G77), .B2(new_n811), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT93), .Z(new_n820));
  NAND2_X1  g0620(.A1(new_n806), .A2(G159), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n821), .A2(KEYINPUT32), .B1(new_n214), .B2(new_n813), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(KEYINPUT32), .B2(new_n821), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n799), .A2(new_n361), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n283), .B1(new_n797), .B2(new_n523), .ZN(new_n825));
  INV_X1    g0625(.A(new_n794), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n824), .B(new_n825), .C1(G68), .C2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n816), .B1(new_n820), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n790), .B1(new_n829), .B2(new_n787), .ZN(new_n830));
  INV_X1    g0630(.A(new_n786), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n830), .B1(new_n710), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n774), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(G396));
  NAND2_X1  g0634(.A1(new_n358), .A2(new_n706), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n369), .B1(new_n365), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n369), .A2(new_n707), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n765), .B(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n772), .B1(new_n840), .B2(new_n760), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n760), .B2(new_n840), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n809), .A2(G143), .B1(G150), .B2(new_n826), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n811), .A2(G159), .B1(new_n803), .B2(G137), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OR2_X1    g0645(.A1(new_n845), .A2(KEYINPUT34), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n799), .A2(new_n202), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n797), .A2(new_n212), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n847), .B(new_n848), .C1(G132), .C2(new_n806), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n377), .B1(G58), .B2(new_n814), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n846), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(KEYINPUT34), .B2(new_n845), .ZN(new_n852));
  AOI22_X1  g0652(.A1(G87), .A2(new_n800), .B1(new_n806), .B2(G311), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(KEYINPUT95), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n802), .A2(new_n380), .B1(new_n797), .B2(new_n361), .ZN(new_n855));
  INV_X1    g0655(.A(G294), .ZN(new_n856));
  INV_X1    g0656(.A(new_n811), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n817), .A2(new_n856), .B1(new_n857), .B2(new_n405), .ZN(new_n858));
  INV_X1    g0658(.A(G283), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n563), .B1(new_n813), .B2(new_n214), .C1(new_n859), .C2(new_n794), .ZN(new_n860));
  NOR4_X1   g0660(.A1(new_n854), .A2(new_n855), .A3(new_n858), .A4(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n787), .B1(new_n852), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n787), .A2(new_n784), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT94), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n775), .B1(new_n286), .B2(new_n865), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n862), .B(new_n866), .C1(new_n839), .C2(new_n785), .ZN(new_n867));
  XOR2_X1   g0667(.A(new_n867), .B(KEYINPUT96), .Z(new_n868));
  NAND2_X1  g0668(.A1(new_n842), .A2(new_n868), .ZN(G384));
  OAI211_X1 g0669(.A(G116), .B(new_n229), .C1(new_n571), .C2(KEYINPUT35), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(KEYINPUT35), .B2(new_n571), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(KEYINPUT36), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n227), .A2(G77), .A3(new_n603), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n212), .A2(G68), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n206), .B(G13), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT98), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n609), .B1(new_n611), .B2(new_n612), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n878), .A2(new_n614), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n613), .A2(new_n270), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n639), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n704), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n658), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n651), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n704), .B1(new_n885), .B2(new_n649), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n641), .A2(new_n643), .B1(new_n886), .B2(new_n881), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n641), .A2(new_n643), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n645), .A2(new_n882), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n652), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  OAI22_X1  g0691(.A1(new_n887), .A2(new_n888), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n884), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n884), .A2(KEYINPUT38), .A3(new_n892), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n895), .A2(KEYINPUT97), .A3(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT97), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n884), .A2(new_n892), .A3(new_n898), .A4(KEYINPUT38), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n897), .A2(KEYINPUT39), .A3(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT39), .ZN(new_n901));
  INV_X1    g0701(.A(new_n890), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n641), .A2(new_n643), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n903), .A2(new_n888), .A3(new_n652), .A4(new_n890), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n652), .A2(new_n640), .A3(new_n890), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT37), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n658), .A2(new_n902), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n896), .B(new_n901), .C1(KEYINPUT38), .C2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n900), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n662), .A2(new_n707), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n660), .A2(new_n704), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n897), .A2(new_n899), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n349), .A2(new_n706), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n350), .A2(new_n916), .B1(new_n662), .B2(new_n706), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n839), .ZN(new_n919));
  NOR3_X1   g0719(.A1(new_n696), .A2(new_n706), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n918), .B1(new_n920), .B2(new_n838), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n914), .B1(new_n915), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n877), .B1(new_n912), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n910), .B1(new_n900), .B2(new_n908), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n897), .A2(new_n899), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n913), .B1(new_n926), .B2(new_n921), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n925), .A2(new_n927), .A3(KEYINPUT98), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n924), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n679), .A2(new_n503), .A3(new_n680), .ZN(new_n930));
  NOR3_X1   g0730(.A1(new_n930), .A2(new_n716), .A3(new_n438), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n931), .A2(new_n707), .B1(new_n756), .B2(new_n755), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n750), .A2(new_n754), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n933), .A2(KEYINPUT99), .A3(KEYINPUT31), .A4(new_n706), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT99), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n758), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  AOI211_X1 g0737(.A(new_n919), .B(new_n917), .C1(new_n932), .C2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT40), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n938), .A2(new_n939), .A3(new_n899), .A4(new_n897), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n919), .B1(new_n932), .B2(new_n937), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n896), .B1(new_n907), .B2(KEYINPUT38), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n941), .A2(new_n942), .A3(new_n918), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(KEYINPUT40), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(G330), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n932), .A2(new_n937), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n371), .A2(new_n658), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n947), .A2(new_n948), .A3(G330), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n947), .A2(new_n948), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n946), .A2(new_n949), .B1(new_n945), .B2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n929), .B(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n741), .A2(new_n766), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n670), .B1(new_n953), .B2(new_n948), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n206), .B2(new_n700), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n952), .A2(new_n954), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n876), .B1(new_n956), .B2(new_n957), .ZN(G367));
  XNOR2_X1  g0758(.A(new_n728), .B(KEYINPUT41), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n706), .B1(new_n579), .B2(new_n580), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n679), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n671), .A2(new_n706), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n725), .B2(new_n722), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT44), .Z(new_n966));
  NOR3_X1   g0766(.A1(new_n725), .A2(new_n722), .A3(new_n964), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT45), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n966), .A2(new_n968), .A3(new_n720), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n720), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n971), .A2(new_n725), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n713), .A2(new_n719), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n768), .ZN(new_n976));
  OAI21_X1  g0776(.A(KEYINPUT102), .B1(new_n970), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n974), .A2(new_n767), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT102), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n978), .A2(new_n969), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n959), .B1(new_n982), .B2(new_n767), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n770), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n725), .A2(new_n679), .A3(new_n960), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n985), .A2(KEYINPUT42), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n676), .B1(new_n964), .B2(new_n500), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n985), .A2(KEYINPUT42), .B1(new_n707), .B2(new_n987), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n535), .A2(new_n707), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n680), .A2(new_n989), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n989), .A2(new_n553), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n986), .A2(new_n988), .B1(KEYINPUT43), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n993), .B(new_n994), .Z(new_n995));
  INV_X1    g0795(.A(KEYINPUT101), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n720), .A2(new_n964), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT100), .ZN(new_n998));
  OR3_X1    g0798(.A1(new_n995), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n995), .A2(new_n998), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n996), .B1(new_n995), .B2(new_n998), .ZN(new_n1001));
  AND3_X1   g0801(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n984), .A2(new_n1002), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n788), .B1(new_n231), .B2(new_n354), .C1(new_n780), .C2(new_n243), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n776), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(G143), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n802), .A2(new_n1006), .B1(new_n799), .B2(new_n286), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n797), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n563), .B(new_n1007), .C1(G58), .C2(new_n1008), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(G159), .A2(new_n826), .B1(new_n806), .B2(G137), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(G150), .A2(new_n809), .B1(new_n811), .B2(G50), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n814), .A2(G68), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(KEYINPUT103), .B(KEYINPUT46), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n797), .B2(new_n405), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1015), .B(new_n377), .C1(new_n361), .C2(new_n813), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n809), .A2(G303), .B1(new_n803), .B2(G311), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n811), .A2(G283), .B1(new_n826), .B2(G294), .ZN(new_n1018));
  AND2_X1   g0818(.A1(KEYINPUT46), .A2(G116), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n1008), .A2(new_n1019), .B1(new_n800), .B2(new_n412), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n806), .A2(G317), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1017), .A2(new_n1018), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1013), .B1(new_n1016), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT47), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n787), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1005), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n990), .A2(new_n786), .A3(new_n991), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1003), .A2(new_n1030), .ZN(G387));
  NAND2_X1  g0831(.A1(new_n717), .A2(new_n786), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(G317), .A2(new_n809), .B1(new_n811), .B2(G303), .ZN(new_n1033));
  XOR2_X1   g0833(.A(KEYINPUT106), .B(G322), .Z(new_n1034));
  AOI22_X1  g0834(.A1(new_n803), .A2(new_n1034), .B1(new_n826), .B2(G311), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT48), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n859), .B2(new_n813), .C1(new_n856), .C2(new_n797), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT49), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n408), .A2(new_n800), .B1(new_n806), .B2(G326), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1040), .A2(new_n377), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n799), .A2(new_n214), .B1(new_n805), .B2(new_n262), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n377), .B(new_n1044), .C1(G77), .C2(new_n1008), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT104), .Z(new_n1046));
  AOI22_X1  g0846(.A1(G159), .A2(new_n803), .B1(new_n826), .B2(new_n352), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n202), .B2(new_n857), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT105), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n809), .A2(G50), .B1(new_n355), .B2(new_n814), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1048), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1046), .B(new_n1051), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1026), .B1(new_n1043), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n779), .B1(new_n240), .B2(new_n386), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n731), .A2(new_n231), .A3(new_n283), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n352), .A2(new_n212), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n386), .B1(new_n202), .B2(new_n286), .C1(new_n1057), .C2(KEYINPUT50), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n731), .B(new_n1058), .C1(KEYINPUT50), .C2(new_n1057), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n1056), .A2(new_n1059), .B1(G107), .B2(new_n231), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n775), .B(new_n1053), .C1(new_n788), .C2(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n975), .A2(new_n771), .B1(new_n1032), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT107), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n974), .A2(new_n1063), .A3(new_n767), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n976), .A2(new_n728), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1063), .B1(new_n974), .B2(new_n767), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1062), .B1(new_n1065), .B2(new_n1066), .ZN(G393));
  OAI221_X1 g0867(.A(new_n788), .B1(new_n231), .B2(new_n419), .C1(new_n780), .C2(new_n250), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n776), .A2(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT109), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n809), .A2(G311), .B1(new_n803), .B2(G317), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT52), .Z(new_n1072));
  AOI22_X1  g0872(.A1(new_n811), .A2(G294), .B1(new_n1008), .B2(G283), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G303), .A2(new_n826), .B1(new_n806), .B2(new_n1034), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n283), .B(new_n824), .C1(new_n408), .C2(new_n814), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT112), .Z(new_n1077));
  AOI22_X1  g0877(.A1(new_n809), .A2(G159), .B1(new_n803), .B2(G150), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT110), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1079), .A2(KEYINPUT51), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(KEYINPUT51), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G50), .A2(new_n826), .B1(new_n800), .B2(G87), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n268), .B2(new_n857), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n813), .A2(new_n286), .ZN(new_n1084));
  NOR3_X1   g0884(.A1(new_n1083), .A2(new_n377), .A3(new_n1084), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n797), .A2(new_n202), .B1(new_n805), .B2(new_n1006), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT111), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1081), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1077), .B1(new_n1080), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1070), .B1(new_n787), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n964), .A2(KEYINPUT108), .A3(new_n786), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT108), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n963), .B2(new_n831), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1090), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n720), .B1(new_n966), .B2(new_n968), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n969), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1094), .B1(new_n1097), .B2(new_n770), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n729), .B1(new_n1097), .B2(new_n976), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT113), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1100), .A2(new_n981), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1101), .B1(new_n1100), .B2(new_n981), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1099), .B1(new_n1103), .B2(new_n1104), .ZN(G390));
  INV_X1    g0905(.A(KEYINPUT116), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n836), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n838), .B1(new_n739), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n918), .B1(new_n941), .B2(G330), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1108), .B1(new_n1109), .B2(KEYINPUT115), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT115), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n758), .B(KEYINPUT99), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n757), .B1(new_n599), .B2(new_n706), .ZN(new_n1113));
  OAI211_X1 g0913(.A(G330), .B(new_n839), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n917), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n918), .A2(new_n759), .A3(G330), .A4(new_n839), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1111), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1106), .B1(new_n1110), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1116), .ZN(new_n1119));
  OAI21_X1  g0919(.A(KEYINPUT115), .B1(new_n1109), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n734), .A2(new_n738), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1121), .A2(new_n707), .A3(new_n1107), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n837), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n1115), .B2(new_n1111), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1120), .A2(new_n1124), .A3(KEYINPUT116), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1118), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n838), .B1(new_n765), .B2(new_n839), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n947), .A2(new_n839), .A3(new_n918), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1128), .A2(new_n712), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n917), .B1(new_n760), .B2(new_n919), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1127), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1126), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n954), .A2(new_n949), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n910), .B1(new_n1127), .B2(new_n917), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n900), .A2(new_n1138), .A3(new_n908), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n911), .B1(new_n1123), .B2(new_n918), .ZN(new_n1140));
  AOI21_X1  g0940(.A(KEYINPUT114), .B1(new_n1140), .B2(new_n942), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n706), .B(new_n836), .C1(new_n734), .C2(new_n738), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n918), .B1(new_n1142), .B2(new_n838), .ZN(new_n1143));
  AND4_X1   g0943(.A1(KEYINPUT114), .A2(new_n1143), .A3(new_n910), .A4(new_n942), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1139), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n1129), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1143), .A2(new_n910), .A3(new_n942), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT114), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1140), .A2(KEYINPUT114), .A3(new_n942), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1151), .A2(new_n1116), .A3(new_n1139), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1146), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1137), .A2(new_n1153), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1146), .A2(new_n1152), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1155), .A2(new_n1136), .A3(new_n1134), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1154), .A2(new_n728), .A3(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n900), .A2(new_n784), .A3(new_n908), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n776), .B1(new_n352), .B2(new_n864), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n817), .A2(new_n401), .B1(new_n802), .B2(new_n859), .ZN(new_n1160));
  NOR4_X1   g0960(.A1(new_n1160), .A2(new_n283), .A3(new_n847), .A4(new_n1084), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(G107), .A2(new_n826), .B1(new_n806), .B2(G294), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n811), .A2(new_n412), .B1(new_n1008), .B2(G87), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n563), .B1(new_n806), .B2(G125), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n212), .B2(new_n799), .ZN(new_n1166));
  XOR2_X1   g0966(.A(new_n1166), .B(KEYINPUT117), .Z(new_n1167));
  NAND2_X1  g0967(.A1(new_n1008), .A2(G150), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1168), .A2(KEYINPUT53), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n1168), .A2(KEYINPUT53), .B1(new_n814), .B2(G159), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n809), .A2(G132), .B1(new_n803), .B2(G128), .ZN(new_n1171));
  XOR2_X1   g0971(.A(KEYINPUT54), .B(G143), .Z(new_n1172));
  AOI22_X1  g0972(.A1(new_n811), .A2(new_n1172), .B1(new_n826), .B2(G137), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .A4(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1164), .B1(new_n1167), .B2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1159), .B1(new_n787), .B2(new_n1175), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1155), .A2(new_n771), .B1(new_n1158), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1157), .A2(new_n1177), .ZN(G378));
  AOI21_X1  g0978(.A(new_n1132), .B1(new_n1118), .B2(new_n1125), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1136), .B1(new_n1153), .B2(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT55), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n314), .A2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n274), .A2(new_n704), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n305), .A2(new_n310), .A3(KEYINPUT55), .A4(new_n313), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n1184), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1186), .B1(new_n1184), .B2(new_n1187), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1182), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1184), .A2(new_n1187), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n1185), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1184), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1192), .A2(new_n1181), .A3(new_n1193), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1190), .A2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1128), .A2(KEYINPUT40), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n1196), .A2(new_n915), .B1(KEYINPUT40), .B2(new_n943), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1195), .B1(new_n1197), .B2(new_n712), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1195), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n945), .A2(G330), .A3(new_n1199), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1198), .B(new_n1200), .C1(new_n924), .C2(new_n928), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n912), .A2(new_n923), .A3(new_n877), .ZN(new_n1202));
  OAI21_X1  g1002(.A(KEYINPUT98), .B1(new_n925), .B2(new_n927), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1199), .B1(new_n945), .B2(G330), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n712), .B(new_n1195), .C1(new_n940), .C2(new_n944), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1202), .B(new_n1203), .C1(new_n1204), .C2(new_n1205), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1180), .A2(KEYINPUT57), .A3(new_n1201), .A4(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT121), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1201), .A2(new_n1206), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1210), .A2(KEYINPUT121), .A3(KEYINPUT57), .A4(new_n1180), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT57), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1135), .B1(new_n1155), .B2(new_n1134), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1201), .A2(new_n1206), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1212), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1209), .A2(new_n1211), .A3(new_n728), .A4(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n799), .A2(new_n201), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G116), .B2(new_n803), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1218), .B1(new_n214), .B2(new_n794), .C1(new_n354), .C2(new_n857), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1012), .B1(new_n859), .B2(new_n805), .C1(new_n817), .C2(new_n361), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n377), .B(new_n290), .C1(new_n286), .C2(new_n797), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT118), .ZN(new_n1223));
  AND2_X1   g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1221), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT58), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n377), .A2(new_n290), .ZN(new_n1228));
  AOI21_X1  g1028(.A(G50), .B1(new_n265), .B2(new_n290), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1226), .A2(new_n1227), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n811), .A2(G137), .B1(new_n1008), .B2(new_n1172), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n809), .A2(G128), .B1(G132), .B2(new_n826), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n803), .A2(G125), .B1(new_n814), .B2(G150), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT119), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1231), .B(new_n1232), .C1(new_n1235), .C2(new_n1236), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1237), .A2(KEYINPUT59), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(KEYINPUT59), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n265), .B(new_n290), .C1(new_n799), .C2(new_n600), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(G124), .B2(new_n806), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n1230), .B1(new_n1227), .B2(new_n1226), .C1(new_n1238), .C2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n787), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n771), .B(new_n728), .C1(new_n212), .C2(new_n865), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1244), .B(new_n1245), .C1(new_n1195), .C2(new_n785), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n1210), .B2(new_n771), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1216), .A2(new_n1248), .ZN(G375));
  NAND2_X1  g1049(.A1(new_n1179), .A2(new_n1135), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1137), .A2(new_n959), .A3(new_n1250), .ZN(new_n1251));
  XOR2_X1   g1051(.A(new_n770), .B(KEYINPUT122), .Z(new_n1252));
  NAND2_X1  g1052(.A1(new_n917), .A2(new_n784), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n776), .B1(G68), .B2(new_n864), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n811), .A2(G107), .B1(new_n1008), .B2(G97), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n283), .B1(new_n800), .B2(G77), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1255), .B(new_n1256), .C1(new_n354), .C2(new_n813), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n817), .A2(new_n859), .B1(new_n805), .B2(new_n380), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n802), .A2(new_n856), .B1(new_n794), .B2(new_n405), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  OR2_X1    g1061(.A1(new_n1261), .A2(KEYINPUT123), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n857), .A2(new_n262), .B1(new_n600), .B2(new_n797), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(new_n826), .B2(new_n1172), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1217), .B1(G132), .B2(new_n803), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n809), .A2(G137), .B1(G128), .B2(new_n806), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n377), .B1(G50), .B2(new_n814), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1264), .A2(new_n1265), .A3(new_n1266), .A4(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1261), .A2(KEYINPUT123), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1262), .A2(new_n1268), .A3(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1254), .B1(new_n1270), .B2(new_n787), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n1134), .A2(new_n1252), .B1(new_n1253), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1251), .A2(new_n1272), .ZN(G381));
  OAI211_X1 g1073(.A(new_n833), .B(new_n1062), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1274));
  OR2_X1    g1074(.A1(new_n1274), .A2(G384), .ZN(new_n1275));
  NOR4_X1   g1075(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(G378), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1216), .A2(new_n1277), .A3(new_n1248), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1276), .A2(new_n1278), .ZN(G407));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n705), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(G407), .A2(G213), .A3(new_n1280), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1281), .B(KEYINPUT124), .ZN(G409));
  NAND2_X1  g1082(.A1(G393), .A2(G396), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1274), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(KEYINPUT126), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT126), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1283), .A2(new_n1286), .A3(new_n1274), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1104), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1098), .B1(new_n1289), .B2(new_n1102), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(G390), .A2(new_n1287), .A3(new_n1285), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(G387), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1291), .A2(new_n1292), .A3(new_n1030), .A4(new_n1003), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1277), .B1(new_n1216), .B2(new_n1248), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n842), .A2(KEYINPUT125), .A3(new_n868), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1272), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT60), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1250), .A2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1179), .A2(KEYINPUT60), .A3(new_n1135), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1302), .A2(new_n728), .A3(new_n1137), .A4(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT125), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(G384), .A2(new_n1305), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n1300), .A2(new_n1304), .A3(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1306), .B1(new_n1300), .B2(new_n1304), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1157), .A2(new_n1177), .A3(new_n1246), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1252), .B1(new_n1180), .B2(new_n959), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1311), .A2(new_n1214), .ZN(new_n1312));
  INV_X1    g1112(.A(G213), .ZN(new_n1313));
  OAI22_X1  g1113(.A1(new_n1310), .A2(new_n1312), .B1(new_n1313), .B2(G343), .ZN(new_n1314));
  NOR3_X1   g1114(.A1(new_n1297), .A2(new_n1309), .A3(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1296), .B1(KEYINPUT63), .B2(new_n1315), .ZN(new_n1316));
  OR2_X1    g1116(.A1(new_n1315), .A2(KEYINPUT63), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT61), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1308), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1300), .A2(new_n1304), .A3(new_n1306), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1313), .A2(G343), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(G2897), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1319), .A2(new_n1320), .A3(new_n1323), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1322), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1325));
  OAI211_X1 g1125(.A(new_n1324), .B(new_n1325), .C1(new_n1297), .C2(new_n1314), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1316), .A2(new_n1317), .A3(new_n1318), .A4(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT62), .ZN(new_n1328));
  OAI211_X1 g1128(.A(new_n1326), .B(new_n1318), .C1(new_n1315), .C2(new_n1328), .ZN(new_n1329));
  AND2_X1   g1129(.A1(new_n1315), .A2(new_n1328), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1296), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1327), .A2(new_n1331), .ZN(G405));
  INV_X1    g1132(.A(KEYINPUT127), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1333), .B1(new_n1278), .B2(new_n1297), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(G375), .A2(G378), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1216), .A2(new_n1277), .A3(new_n1248), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1335), .A2(KEYINPUT127), .A3(new_n1336), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1334), .A2(new_n1337), .A3(new_n1309), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1296), .ZN(new_n1339));
  OAI221_X1 g1139(.A(new_n1333), .B1(new_n1308), .B2(new_n1307), .C1(new_n1278), .C2(new_n1297), .ZN(new_n1340));
  AND3_X1   g1140(.A1(new_n1338), .A2(new_n1339), .A3(new_n1340), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1339), .B1(new_n1338), .B2(new_n1340), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1341), .A2(new_n1342), .ZN(G402));
endmodule


