//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 1 0 0 0 1 1 0 1 0 1 1 0 0 0 1 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 1 0 0 0 1 1 1 0 0 0 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n520, new_n521,
    new_n522, new_n523, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n537, new_n538,
    new_n539, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n610, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177, new_n1178,
    new_n1179;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  XNOR2_X1  g032(.A(KEYINPUT3), .B(G2104), .ZN(new_n458));
  AOI22_X1  g033(.A1(new_n458), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  AND3_X1   g039(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(KEYINPUT3), .B1(KEYINPUT66), .B2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n464), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n461), .A2(new_n469), .ZN(G160));
  OAI21_X1  g045(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(G112), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n471), .B1(new_n472), .B2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(new_n467), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n474), .A2(G136), .ZN(new_n475));
  OAI21_X1  g050(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT67), .ZN(new_n477));
  AOI211_X1 g052(.A(new_n473), .B(new_n475), .C1(G124), .C2(new_n477), .ZN(G162));
  INV_X1    g053(.A(G138), .ZN(new_n479));
  OAI21_X1  g054(.A(KEYINPUT4), .B1(new_n467), .B2(new_n479), .ZN(new_n480));
  NOR3_X1   g055(.A1(new_n479), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n458), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G114), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n476), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(G126), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n483), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G164));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT6), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(G651), .ZN(new_n493));
  INV_X1    g068(.A(G651), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n494), .A2(KEYINPUT68), .A3(KEYINPUT6), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n493), .A2(new_n495), .B1(new_n492), .B2(G651), .ZN(new_n496));
  XNOR2_X1  g071(.A(KEYINPUT5), .B(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G88), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n493), .A2(new_n495), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n492), .A2(G651), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n501), .A2(G543), .A3(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G50), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n497), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  OR2_X1    g081(.A1(new_n506), .A2(new_n494), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n500), .A2(new_n505), .A3(new_n507), .ZN(G303));
  INV_X1    g083(.A(G303), .ZN(G166));
  NAND3_X1  g084(.A1(new_n496), .A2(G89), .A3(new_n497), .ZN(new_n510));
  XOR2_X1   g085(.A(KEYINPUT69), .B(G51), .Z(new_n511));
  NAND3_X1  g086(.A1(new_n496), .A2(G543), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n513), .A2(KEYINPUT7), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(KEYINPUT7), .ZN(new_n515));
  AND2_X1   g090(.A1(G63), .A2(G651), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n514), .A2(new_n515), .B1(new_n497), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n510), .A2(new_n512), .A3(new_n517), .ZN(G286));
  INV_X1    g093(.A(G286), .ZN(G168));
  AOI22_X1  g094(.A1(new_n497), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n520), .A2(new_n494), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n496), .A2(G90), .A3(new_n497), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n496), .A2(G52), .A3(G543), .ZN(new_n523));
  AND3_X1   g098(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(G171));
  NAND3_X1  g099(.A1(new_n496), .A2(G81), .A3(new_n497), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n496), .A2(G43), .A3(G543), .ZN(new_n526));
  INV_X1    g101(.A(G56), .ZN(new_n527));
  OR2_X1    g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(KEYINPUT5), .A2(G543), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AND2_X1   g105(.A1(G68), .A2(G543), .ZN(new_n531));
  OAI21_X1  g106(.A(G651), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n525), .A2(new_n526), .A3(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G860), .ZN(G153));
  NAND4_X1  g110(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g111(.A1(G1), .A2(G3), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT70), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT8), .ZN(new_n539));
  NAND4_X1  g114(.A1(G319), .A2(G483), .A3(G661), .A4(new_n539), .ZN(G188));
  NAND4_X1  g115(.A1(new_n501), .A2(G53), .A3(G543), .A4(new_n502), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(KEYINPUT9), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT9), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n496), .A2(new_n543), .A3(G53), .A4(G543), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  AND2_X1   g120(.A1(KEYINPUT5), .A2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(KEYINPUT5), .A2(G543), .ZN(new_n547));
  OAI21_X1  g122(.A(G65), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(G78), .A2(G543), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n548), .A2(KEYINPUT71), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G651), .ZN(new_n551));
  AOI21_X1  g126(.A(KEYINPUT71), .B1(new_n548), .B2(new_n549), .ZN(new_n552));
  INV_X1    g127(.A(G91), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n551), .A2(new_n552), .B1(new_n553), .B2(new_n498), .ZN(new_n554));
  OAI21_X1  g129(.A(KEYINPUT72), .B1(new_n545), .B2(new_n554), .ZN(new_n555));
  AND4_X1   g130(.A1(G91), .A2(new_n501), .A3(new_n502), .A4(new_n497), .ZN(new_n556));
  INV_X1    g131(.A(new_n549), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n557), .B1(new_n497), .B2(G65), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n494), .B1(new_n558), .B2(KEYINPUT71), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n548), .A2(new_n549), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT71), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n556), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT72), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n542), .A2(new_n544), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n555), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G299));
  NAND3_X1  g143(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(G301));
  OAI21_X1  g144(.A(G651), .B1(new_n497), .B2(G74), .ZN(new_n570));
  INV_X1    g145(.A(G49), .ZN(new_n571));
  INV_X1    g146(.A(G87), .ZN(new_n572));
  OAI221_X1 g147(.A(new_n570), .B1(new_n503), .B2(new_n571), .C1(new_n498), .C2(new_n572), .ZN(G288));
  NAND2_X1  g148(.A1(new_n499), .A2(G86), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n504), .A2(G48), .ZN(new_n575));
  AND2_X1   g150(.A1(new_n497), .A2(G61), .ZN(new_n576));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT73), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n574), .A2(new_n575), .A3(new_n579), .ZN(G305));
  NAND2_X1  g155(.A1(new_n499), .A2(G85), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n504), .A2(G47), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n497), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n583), .A2(new_n494), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n581), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT74), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n585), .A2(new_n586), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(G290));
  INV_X1    g164(.A(G868), .ZN(new_n590));
  NOR2_X1   g165(.A1(G301), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(G54), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n497), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n593));
  OAI22_X1  g168(.A1(new_n503), .A2(new_n592), .B1(new_n593), .B2(new_n494), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n501), .A2(G92), .A3(new_n502), .A4(new_n497), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n596), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n594), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AND2_X1   g174(.A1(new_n599), .A2(KEYINPUT75), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n599), .A2(KEYINPUT75), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n591), .B1(new_n603), .B2(new_n590), .ZN(G284));
  AOI21_X1  g179(.A(new_n591), .B1(new_n603), .B2(new_n590), .ZN(G321));
  NOR2_X1   g180(.A1(G286), .A2(new_n590), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n567), .B(KEYINPUT76), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(new_n590), .ZN(G297));
  AOI21_X1  g183(.A(new_n606), .B1(new_n607), .B2(new_n590), .ZN(G280));
  NOR2_X1   g184(.A1(new_n602), .A2(G559), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(G860), .B2(new_n603), .ZN(G148));
  NAND2_X1  g186(.A1(new_n533), .A2(new_n590), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(new_n610), .B2(new_n590), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g189(.A1(new_n458), .A2(new_n463), .ZN(new_n615));
  XNOR2_X1  g190(.A(KEYINPUT77), .B(KEYINPUT12), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT13), .ZN(new_n619));
  INV_X1    g194(.A(G2100), .ZN(new_n620));
  OAI22_X1  g195(.A1(new_n618), .A2(new_n619), .B1(KEYINPUT78), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(new_n619), .B2(new_n618), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(KEYINPUT78), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n477), .A2(G123), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n474), .A2(G135), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n460), .A2(G111), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n625), .B(new_n626), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2096), .Z(new_n630));
  NAND2_X1  g205(.A1(new_n624), .A2(new_n630), .ZN(G156));
  XOR2_X1   g206(.A(KEYINPUT15), .B(G2435), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2427), .B(G2430), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT79), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n633), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(KEYINPUT14), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n638), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(new_n646), .A3(G14), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT80), .Z(G401));
  XNOR2_X1  g223(.A(G2072), .B(G2078), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT17), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  NOR3_X1   g228(.A1(new_n650), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT81), .Z(new_n655));
  NAND2_X1  g230(.A1(new_n650), .A2(new_n651), .ZN(new_n656));
  OAI211_X1 g231(.A(new_n656), .B(new_n653), .C1(new_n649), .C2(new_n651), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n652), .A2(new_n649), .A3(new_n651), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT18), .Z(new_n659));
  NAND3_X1  g234(.A1(new_n655), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2096), .B(G2100), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(G227));
  XOR2_X1   g237(.A(G1971), .B(G1976), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  XOR2_X1   g239(.A(G1956), .B(G2474), .Z(new_n665));
  XOR2_X1   g240(.A(G1961), .B(G1966), .Z(new_n666));
  AND2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT20), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n665), .A2(new_n666), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n664), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n671), .B1(new_n664), .B2(new_n670), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n673), .B(new_n674), .Z(new_n675));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1981), .B(G1986), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(G229));
  INV_X1    g255(.A(G29), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n681), .B1(KEYINPUT24), .B2(G34), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(KEYINPUT24), .B2(G34), .ZN(new_n683));
  INV_X1    g258(.A(G160), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n683), .B1(new_n684), .B2(G29), .ZN(new_n685));
  INV_X1    g260(.A(G2084), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT92), .Z(new_n688));
  NAND3_X1  g263(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT26), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n463), .A2(G105), .ZN(new_n691));
  AOI211_X1 g266(.A(new_n690), .B(new_n691), .C1(G141), .C2(new_n474), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n477), .A2(G129), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n695), .A2(new_n681), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n681), .B2(G32), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT27), .B(G1996), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n688), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n681), .A2(G33), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n458), .A2(G127), .ZN(new_n701));
  INV_X1    g276(.A(G115), .ZN(new_n702));
  INV_X1    g277(.A(G2104), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT90), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n460), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(new_n705), .B2(new_n704), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT91), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT25), .Z(new_n711));
  INV_X1    g286(.A(G139), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n467), .B2(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT89), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n700), .B1(new_n716), .B2(new_n681), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n699), .B1(G2072), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G2072), .B2(new_n717), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT93), .Z(new_n720));
  NOR2_X1   g295(.A1(G4), .A2(G16), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT84), .ZN(new_n722));
  INV_X1    g297(.A(G16), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n602), .B2(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G1348), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n681), .A2(G26), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT28), .Z(new_n727));
  NAND2_X1  g302(.A1(new_n477), .A2(G128), .ZN(new_n728));
  NOR2_X1   g303(.A1(G104), .A2(G2105), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT86), .Z(new_n730));
  INV_X1    g305(.A(G116), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n703), .B1(new_n731), .B2(G2105), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n730), .A2(new_n732), .B1(new_n474), .B2(G140), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n728), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n727), .B1(new_n734), .B2(G29), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT87), .ZN(new_n736));
  INV_X1    g311(.A(G2067), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(G16), .A2(G19), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n534), .B2(G16), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT85), .B(G1341), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n725), .A2(new_n738), .A3(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT88), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n723), .A2(G22), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G166), .B2(new_n723), .ZN(new_n746));
  INV_X1    g321(.A(G1971), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(G6), .A2(G16), .ZN(new_n749));
  INV_X1    g324(.A(G305), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n749), .B1(new_n750), .B2(G16), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT32), .B(G1981), .Z(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n723), .A2(G23), .ZN(new_n754));
  INV_X1    g329(.A(G288), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n754), .B1(new_n755), .B2(new_n723), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT33), .B(G1976), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  AND3_X1   g333(.A1(new_n748), .A2(new_n753), .A3(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n760), .A2(KEYINPUT34), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n760), .A2(KEYINPUT34), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n681), .A2(G25), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n474), .A2(G131), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT82), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n477), .A2(G119), .ZN(new_n766));
  OR2_X1    g341(.A1(G95), .A2(G2105), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n767), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n765), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n763), .B1(new_n770), .B2(new_n681), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT35), .B(G1991), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n723), .A2(G24), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G290), .B2(G16), .ZN(new_n775));
  INV_X1    g350(.A(G1986), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n773), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  NOR3_X1   g355(.A1(new_n761), .A2(new_n762), .A3(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT36), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n782), .A2(KEYINPUT83), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n744), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n782), .A2(KEYINPUT83), .ZN(new_n785));
  OR3_X1    g360(.A1(new_n781), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n685), .A2(new_n686), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n723), .A2(G5), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G171), .B2(new_n723), .ZN(new_n789));
  OAI221_X1 g364(.A(new_n787), .B1(new_n789), .B2(G1961), .C1(new_n697), .C2(new_n698), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT95), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n681), .A2(G35), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G162), .B2(new_n681), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT29), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G2090), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n723), .A2(G20), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT23), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n567), .B2(new_n723), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G1956), .ZN(new_n799));
  NAND2_X1  g374(.A1(G168), .A2(G16), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n800), .B(KEYINPUT94), .C1(G16), .C2(G21), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(KEYINPUT94), .B2(new_n800), .ZN(new_n802));
  INV_X1    g377(.A(G1966), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT31), .B(G11), .Z(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT30), .B(G28), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n805), .B1(new_n681), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n629), .B2(new_n681), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(G1961), .B2(new_n789), .ZN(new_n809));
  NOR2_X1   g384(.A1(G27), .A2(G29), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G164), .B2(G29), .ZN(new_n811));
  INV_X1    g386(.A(G2078), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n804), .A2(new_n809), .A3(new_n813), .ZN(new_n814));
  NOR4_X1   g389(.A1(new_n791), .A2(new_n795), .A3(new_n799), .A4(new_n814), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n720), .A2(new_n784), .A3(new_n786), .A4(new_n815), .ZN(G150));
  INV_X1    g391(.A(G150), .ZN(G311));
  NAND3_X1  g392(.A1(new_n496), .A2(G93), .A3(new_n497), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n496), .A2(G55), .A3(G543), .ZN(new_n819));
  INV_X1    g394(.A(G67), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(new_n528), .B2(new_n529), .ZN(new_n821));
  AND2_X1   g396(.A1(G80), .A2(G543), .ZN(new_n822));
  OAI21_X1  g397(.A(G651), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n818), .A2(new_n819), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(G860), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT98), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT37), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n603), .A2(G559), .ZN(new_n828));
  XOR2_X1   g403(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT97), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n824), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n818), .A2(new_n819), .A3(KEYINPUT97), .A4(new_n823), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n832), .A2(new_n534), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n533), .A2(new_n824), .A3(new_n831), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n830), .B(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n838), .A2(KEYINPUT39), .ZN(new_n839));
  INV_X1    g414(.A(G860), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n838), .B2(KEYINPUT39), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n827), .B1(new_n839), .B2(new_n841), .ZN(G145));
  INV_X1    g417(.A(KEYINPUT99), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n715), .B(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n734), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(G164), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n734), .A2(new_n489), .ZN(new_n847));
  AND3_X1   g422(.A1(new_n846), .A2(new_n694), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n694), .B1(new_n846), .B2(new_n847), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n844), .A2(new_n850), .ZN(new_n851));
  OAI22_X1  g426(.A1(new_n716), .A2(KEYINPUT99), .B1(new_n848), .B2(new_n849), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n477), .A2(G130), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n474), .A2(G142), .ZN(new_n855));
  OAI21_X1  g430(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n856), .A2(KEYINPUT100), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(KEYINPUT100), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(G118), .B2(new_n460), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n854), .B(new_n855), .C1(new_n857), .C2(new_n859), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n860), .A2(new_n617), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n860), .A2(new_n617), .ZN(new_n862));
  OR3_X1    g437(.A1(new_n861), .A2(new_n862), .A3(new_n769), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n769), .B1(new_n861), .B2(new_n862), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n863), .A2(KEYINPUT101), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n864), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT101), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n853), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n865), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n870), .A2(new_n851), .A3(new_n852), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n629), .B(new_n684), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(G162), .Z(new_n874));
  AOI21_X1  g449(.A(G37), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT102), .ZN(new_n876));
  INV_X1    g451(.A(new_n874), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n871), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n866), .B1(new_n851), .B2(new_n852), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n876), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  AND4_X1   g456(.A1(new_n876), .A2(new_n880), .A3(new_n871), .A4(new_n877), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n875), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g459(.A(new_n610), .B(new_n836), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n555), .A2(new_n566), .A3(new_n599), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n599), .B1(new_n555), .B2(new_n566), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT41), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n597), .A2(new_n598), .ZN(new_n892));
  INV_X1    g467(.A(new_n594), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(KEYINPUT103), .B1(new_n567), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT103), .ZN(new_n896));
  AOI211_X1 g471(.A(new_n896), .B(new_n599), .C1(new_n555), .C2(new_n566), .ZN(new_n897));
  NOR3_X1   g472(.A1(new_n895), .A2(new_n897), .A3(new_n887), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n891), .B1(new_n898), .B2(KEYINPUT41), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n885), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n900), .A2(KEYINPUT104), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT42), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n885), .A2(new_n899), .ZN(new_n904));
  INV_X1    g479(.A(new_n556), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n562), .A2(G651), .A3(new_n550), .ZN(new_n906));
  AND4_X1   g481(.A1(new_n564), .A2(new_n565), .A3(new_n905), .A4(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n564), .B1(new_n563), .B2(new_n565), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n894), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n886), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT104), .B1(new_n885), .B2(new_n911), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n902), .B(new_n903), .C1(new_n904), .C2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n914));
  XNOR2_X1  g489(.A(G288), .B(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n750), .ZN(new_n916));
  XNOR2_X1  g491(.A(G288), .B(KEYINPUT105), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(G305), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(G303), .B1(new_n587), .B2(new_n588), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n587), .A2(new_n588), .A3(G303), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n919), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n920), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n924), .A2(new_n921), .A3(new_n916), .A4(new_n918), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT106), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n904), .A2(new_n912), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT42), .B1(new_n929), .B2(new_n901), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n913), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n928), .B1(new_n913), .B2(new_n930), .ZN(new_n932));
  OAI21_X1  g507(.A(G868), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n824), .A2(new_n590), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(G295));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n934), .ZN(G331));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n923), .A2(new_n925), .ZN(new_n938));
  NAND2_X1  g513(.A1(G171), .A2(G168), .ZN(new_n939));
  NAND2_X1  g514(.A1(G301), .A2(G286), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n836), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n939), .A2(new_n834), .A3(new_n940), .A4(new_n835), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n910), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n938), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT107), .B1(new_n942), .B2(new_n943), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n950), .B1(new_n941), .B2(new_n836), .ZN(new_n951));
  OR2_X1    g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n948), .B1(new_n899), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n909), .A2(new_n896), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n567), .A2(KEYINPUT103), .A3(new_n894), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n954), .A2(new_n886), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n890), .B1(new_n956), .B2(new_n889), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n949), .A2(new_n951), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n957), .A2(KEYINPUT108), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n947), .B1(new_n953), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n895), .A2(new_n897), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n887), .A2(new_n889), .ZN(new_n962));
  AOI22_X1  g537(.A1(new_n961), .A2(new_n962), .B1(new_n910), .B2(new_n889), .ZN(new_n963));
  OAI22_X1  g538(.A1(new_n963), .A2(new_n944), .B1(new_n952), .B2(new_n911), .ZN(new_n964));
  AOI21_X1  g539(.A(G37), .B1(new_n964), .B2(new_n926), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n960), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT109), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n899), .A2(new_n948), .A3(new_n952), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT108), .B1(new_n957), .B2(new_n958), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n946), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(new_n973), .A3(new_n965), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n968), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n945), .B1(new_n953), .B2(new_n959), .ZN(new_n976));
  AOI21_X1  g551(.A(G37), .B1(new_n976), .B2(new_n926), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n966), .B1(new_n977), .B2(new_n960), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n937), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n937), .B1(new_n977), .B2(new_n972), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n962), .A2(new_n954), .A3(new_n955), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n910), .A2(new_n889), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n944), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n949), .A2(new_n911), .A3(new_n951), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n926), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G37), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT110), .B1(new_n971), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n960), .A2(new_n965), .A3(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n988), .A2(new_n990), .A3(KEYINPUT43), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n980), .A2(KEYINPUT111), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT111), .B1(new_n980), .B2(new_n991), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n979), .B1(new_n992), .B2(new_n993), .ZN(G397));
  INV_X1    g569(.A(G1384), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n489), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(G160), .A2(G40), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n1000), .A2(G1996), .A3(new_n694), .ZN(new_n1001));
  XOR2_X1   g576(.A(new_n1001), .B(KEYINPUT112), .Z(new_n1002));
  XNOR2_X1  g577(.A(new_n734), .B(new_n737), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1003), .B1(G1996), .B2(new_n694), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1002), .B1(new_n1000), .B2(new_n1004), .ZN(new_n1005));
  AND2_X1   g580(.A1(new_n770), .A2(new_n772), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n770), .A2(new_n772), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1000), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(G290), .B(G1986), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1009), .B1(new_n1000), .B2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n563), .A2(KEYINPUT57), .A3(new_n565), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n1012), .B(KEYINPUT122), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT57), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n545), .B1(KEYINPUT121), .B2(new_n563), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1015), .B1(KEYINPUT121), .B2(new_n563), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1013), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n996), .A2(KEYINPUT50), .ZN(new_n1018));
  INV_X1    g593(.A(new_n999), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT50), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n489), .A2(new_n1020), .A3(new_n995), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1018), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g597(.A(KEYINPUT120), .B(G1956), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n999), .B1(new_n996), .B2(new_n997), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n489), .A2(KEYINPUT45), .A3(new_n995), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  XOR2_X1   g602(.A(KEYINPUT56), .B(G2072), .Z(new_n1028));
  OAI21_X1  g603(.A(new_n1024), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OR2_X1    g604(.A1(new_n1017), .A2(new_n1029), .ZN(new_n1030));
  OR3_X1    g605(.A1(new_n996), .A2(new_n999), .A3(KEYINPUT123), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT123), .B1(new_n996), .B2(new_n999), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n737), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1018), .A2(KEYINPUT113), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT113), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n996), .A2(new_n1037), .A3(KEYINPUT50), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1035), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1034), .B1(new_n1039), .B2(G1348), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1040), .A2(new_n603), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1017), .A2(new_n1029), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1030), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT60), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1040), .A2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1034), .B(KEYINPUT60), .C1(new_n1039), .C2(G1348), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1046), .A2(new_n603), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT124), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1049), .B1(new_n1017), .B2(new_n1029), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1043), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT61), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(new_n1042), .B2(new_n1049), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1048), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g629(.A(KEYINPUT58), .B(G1341), .ZN(new_n1055));
  OAI22_X1  g630(.A1(new_n1033), .A2(new_n1055), .B1(G1996), .B2(new_n1027), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n534), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT59), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT59), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1056), .A2(new_n1059), .A3(new_n534), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1030), .A2(KEYINPUT61), .A3(new_n1042), .ZN(new_n1062));
  OR2_X1    g637(.A1(new_n1047), .A2(new_n603), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1044), .B1(new_n1054), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT125), .ZN(new_n1066));
  INV_X1    g641(.A(new_n998), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT118), .B1(new_n1067), .B2(new_n999), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1025), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n1026), .B(KEYINPUT119), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n1073), .A2(new_n803), .B1(new_n686), .B2(new_n1039), .ZN(new_n1074));
  INV_X1    g649(.A(G8), .ZN(new_n1075));
  NOR2_X1   g650(.A1(G168), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1066), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1072), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1079), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1039), .ZN(new_n1081));
  OAI22_X1  g656(.A1(new_n1080), .A2(G1966), .B1(G2084), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1082), .A2(KEYINPUT125), .A3(new_n1076), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1078), .A2(new_n1083), .ZN(new_n1084));
  OAI211_X1 g659(.A(KEYINPUT51), .B(new_n1077), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT51), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1086), .B(G8), .C1(new_n1082), .C2(G286), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1084), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n996), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1075), .B1(new_n1089), .B2(new_n1019), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n755), .A2(G1976), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT52), .ZN(new_n1093));
  INV_X1    g668(.A(G1976), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT52), .B1(G288), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1090), .A2(new_n1091), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g672(.A(G305), .B(G1981), .ZN(new_n1098));
  XNOR2_X1  g673(.A(KEYINPUT115), .B(KEYINPUT49), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n1100), .B(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT49), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1090), .B1(new_n1098), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1097), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1027), .A2(new_n747), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(G2090), .B2(new_n1022), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(G8), .ZN(new_n1109));
  NAND2_X1  g684(.A1(G303), .A2(G8), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT55), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  OR2_X1    g687(.A1(new_n1112), .A2(KEYINPUT114), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(KEYINPUT114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1109), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1107), .B1(new_n1081), .B2(G2090), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1119), .A2(G8), .A3(new_n1116), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1106), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1027), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT53), .B1(new_n1122), .B2(new_n812), .ZN(new_n1123));
  INV_X1    g698(.A(G1961), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1123), .B1(new_n1124), .B2(new_n1081), .ZN(new_n1125));
  XNOR2_X1  g700(.A(G301), .B(KEYINPUT54), .ZN(new_n1126));
  OAI21_X1  g701(.A(G2105), .B1(new_n459), .B2(KEYINPUT126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1127), .B1(KEYINPUT126), .B2(new_n459), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n812), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1129));
  NOR4_X1   g704(.A1(new_n1067), .A2(new_n469), .A3(new_n1128), .A4(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1126), .B1(new_n1130), .B2(new_n1026), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1125), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1126), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1080), .A2(KEYINPUT53), .A3(new_n812), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1134), .B1(new_n1125), .B2(new_n1135), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1121), .A2(new_n1133), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1065), .A2(new_n1088), .A3(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(G305), .A2(G1981), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1140));
  NOR2_X1   g715(.A1(G288), .A2(G1976), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1139), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1090), .B(KEYINPUT117), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1106), .ZN(new_n1144));
  OAI22_X1  g719(.A1(new_n1142), .A2(new_n1143), .B1(new_n1144), .B2(new_n1120), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n1106), .A2(new_n1120), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1082), .A2(G8), .A3(G168), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT63), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1119), .A2(G8), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1149), .B1(new_n1150), .B2(new_n1117), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1146), .A2(new_n1148), .A3(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1149), .B1(new_n1121), .B2(new_n1147), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1145), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1138), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(G301), .B1(new_n1135), .B2(new_n1125), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1146), .A2(new_n1118), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT62), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1088), .A2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1084), .A2(KEYINPUT62), .A3(new_n1085), .A4(new_n1087), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1157), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1011), .B1(new_n1155), .B2(new_n1161), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n998), .A2(G1996), .A3(new_n999), .ZN(new_n1163));
  XOR2_X1   g738(.A(new_n1163), .B(KEYINPUT46), .Z(new_n1164));
  INV_X1    g739(.A(new_n1003), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1000), .B1(new_n1165), .B2(new_n694), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT47), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1000), .A2(new_n776), .A3(new_n588), .A4(new_n587), .ZN(new_n1169));
  XOR2_X1   g744(.A(new_n1169), .B(KEYINPUT48), .Z(new_n1170));
  OAI21_X1  g745(.A(new_n1168), .B1(new_n1009), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1172), .B1(G2067), .B2(new_n734), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1171), .B1(new_n1000), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1162), .A2(new_n1174), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g750(.A(G319), .ZN(new_n1177));
  NOR3_X1   g751(.A1(G401), .A2(new_n1177), .A3(G227), .ZN(new_n1178));
  AND2_X1   g752(.A1(new_n1178), .A2(new_n679), .ZN(new_n1179));
  OAI211_X1 g753(.A(new_n883), .B(new_n1179), .C1(new_n975), .C2(new_n978), .ZN(G225));
  INV_X1    g754(.A(G225), .ZN(G308));
endmodule


