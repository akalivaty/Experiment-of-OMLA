//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 1 1 0 0 1 1 1 1 1 1 1 1 0 0 1 1 1 1 1 1 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 0 0 1 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT9), .B(G234), .Z(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n187), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  NOR3_X1   g005(.A1(new_n191), .A2(KEYINPUT3), .A3(G107), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G104), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G101), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n193), .A2(G104), .ZN(new_n197));
  AOI21_X1  g011(.A(KEYINPUT73), .B1(new_n197), .B2(KEYINPUT3), .ZN(new_n198));
  OAI211_X1 g012(.A(KEYINPUT73), .B(KEYINPUT3), .C1(new_n191), .C2(G107), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n195), .B(new_n196), .C1(new_n198), .C2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT75), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT3), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(new_n193), .A3(G104), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n191), .A2(G107), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT3), .B1(new_n191), .B2(G107), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT73), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n206), .B1(new_n209), .B2(new_n199), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT75), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(new_n211), .A3(new_n196), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n202), .A2(new_n212), .A3(KEYINPUT4), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT74), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT4), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n215), .B1(new_n210), .B2(new_n196), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n195), .B1(new_n198), .B2(new_n200), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n217), .A2(new_n214), .A3(KEYINPUT4), .A4(G101), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n213), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(G143), .B(G146), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT0), .ZN(new_n223));
  INV_X1    g037(.A(G128), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NOR3_X1   g039(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n221), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n220), .B1(new_n223), .B2(new_n224), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n219), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT11), .ZN(new_n231));
  INV_X1    g045(.A(G134), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(G137), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(G137), .ZN(new_n234));
  INV_X1    g048(.A(G137), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(KEYINPUT11), .A3(G134), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n233), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G131), .ZN(new_n238));
  INV_X1    g052(.A(G131), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n233), .A2(new_n236), .A3(new_n239), .A4(new_n234), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n196), .B1(new_n197), .B2(new_n205), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G143), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT1), .B1(new_n245), .B2(G146), .ZN(new_n246));
  INV_X1    g060(.A(G146), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G143), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n245), .A2(G146), .ZN(new_n249));
  AOI22_X1  g063(.A1(new_n246), .A2(G128), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT1), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n248), .A2(new_n249), .A3(new_n251), .A4(G128), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT66), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n220), .A2(KEYINPUT66), .A3(new_n251), .A4(G128), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n250), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n201), .A2(KEYINPUT75), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n211), .B1(new_n210), .B2(new_n196), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n244), .B(new_n257), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT10), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n243), .B1(new_n202), .B2(new_n212), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n264), .B(KEYINPUT1), .C1(new_n245), .C2(G146), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G128), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n264), .B1(new_n248), .B2(KEYINPUT1), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n221), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT68), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n254), .A2(new_n255), .ZN(new_n271));
  OAI211_X1 g085(.A(KEYINPUT68), .B(new_n221), .C1(new_n266), .C2(new_n267), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n263), .A2(KEYINPUT10), .A3(new_n273), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n230), .A2(new_n242), .A3(new_n262), .A4(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(G110), .B(G140), .ZN(new_n276));
  INV_X1    g090(.A(G227), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n277), .A2(G953), .ZN(new_n278));
  XOR2_X1   g092(.A(new_n276), .B(new_n278), .Z(new_n279));
  INV_X1    g093(.A(KEYINPUT76), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT12), .B1(new_n241), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n244), .B1(new_n258), .B2(new_n259), .ZN(new_n282));
  INV_X1    g096(.A(new_n273), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI211_X1 g098(.A(new_n242), .B(new_n281), .C1(new_n284), .C2(new_n260), .ZN(new_n285));
  INV_X1    g099(.A(new_n281), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n260), .B1(new_n273), .B2(new_n263), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n286), .B1(new_n287), .B2(new_n241), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n275), .B(new_n279), .C1(new_n285), .C2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT77), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n263), .A2(new_n273), .ZN(new_n292));
  AOI211_X1 g106(.A(new_n243), .B(new_n256), .C1(new_n202), .C2(new_n212), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n241), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n281), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n287), .A2(new_n241), .A3(new_n286), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n297), .A2(KEYINPUT77), .A3(new_n275), .A4(new_n279), .ZN(new_n298));
  INV_X1    g112(.A(new_n279), .ZN(new_n299));
  INV_X1    g113(.A(new_n275), .ZN(new_n300));
  AOI22_X1  g114(.A1(new_n219), .A2(new_n229), .B1(new_n260), .B2(new_n261), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n242), .B1(new_n301), .B2(new_n274), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n299), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n291), .A2(new_n298), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G469), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n305), .A3(new_n189), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT78), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT78), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n304), .A2(new_n308), .A3(new_n305), .A4(new_n189), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n297), .A2(new_n275), .A3(new_n299), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n279), .B1(new_n300), .B2(new_n302), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n312), .A3(new_n189), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G469), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n190), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G119), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G116), .ZN(new_n317));
  INV_X1    g131(.A(G116), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G119), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  XOR2_X1   g134(.A(KEYINPUT2), .B(G113), .Z(new_n321));
  XNOR2_X1  g135(.A(new_n320), .B(new_n321), .ZN(new_n322));
  AOI22_X1  g136(.A1(new_n227), .A2(new_n228), .B1(new_n238), .B2(new_n240), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT65), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n324), .B1(new_n232), .B2(G137), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n235), .A2(KEYINPUT65), .A3(G134), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(new_n234), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G131), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n328), .A2(new_n240), .ZN(new_n329));
  AOI211_X1 g143(.A(new_n322), .B(new_n323), .C1(new_n273), .C2(new_n329), .ZN(new_n330));
  OR2_X1    g144(.A1(new_n330), .A2(KEYINPUT28), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT26), .B(G101), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n332), .B(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G237), .ZN(new_n335));
  INV_X1    g149(.A(G953), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n335), .A2(new_n336), .A3(G210), .ZN(new_n337));
  XOR2_X1   g151(.A(new_n334), .B(new_n337), .Z(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT29), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n322), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n273), .A2(new_n329), .ZN(new_n343));
  INV_X1    g157(.A(new_n323), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(KEYINPUT28), .B1(new_n345), .B2(new_n330), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n346), .A2(KEYINPUT70), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT70), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n348), .B(KEYINPUT28), .C1(new_n345), .C2(new_n330), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n331), .B(new_n341), .C1(new_n347), .C2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT30), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n352), .B1(new_n343), .B2(new_n344), .ZN(new_n353));
  AOI211_X1 g167(.A(KEYINPUT30), .B(new_n323), .C1(new_n273), .C2(new_n329), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n322), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n330), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n339), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n331), .A2(new_n346), .A3(new_n338), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n340), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n351), .A2(new_n360), .A3(new_n189), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G472), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n355), .A2(new_n356), .A3(new_n338), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT31), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n355), .A2(KEYINPUT31), .A3(new_n356), .A4(new_n338), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n331), .A2(new_n346), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n339), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(G472), .A2(G902), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(KEYINPUT32), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT32), .ZN(new_n373));
  AOI22_X1  g187(.A1(new_n365), .A2(new_n366), .B1(new_n368), .B2(new_n339), .ZN(new_n374));
  INV_X1    g188(.A(new_n371), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n362), .A2(new_n372), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n224), .A2(G119), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT23), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n316), .A2(G128), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n224), .A2(KEYINPUT23), .A3(G119), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G110), .ZN(new_n384));
  OR2_X1    g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n381), .A2(new_n378), .ZN(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT24), .B(G110), .ZN(new_n387));
  OR2_X1    g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G140), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G125), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT16), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(KEYINPUT71), .A2(G125), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n394), .B(G140), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n393), .B1(new_n395), .B2(KEYINPUT16), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(new_n247), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n394), .B(new_n389), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n392), .B1(new_n398), .B2(new_n391), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(G146), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n385), .B(new_n388), .C1(new_n397), .C2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT72), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n402), .B1(new_n396), .B2(new_n247), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n383), .A2(new_n384), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n386), .A2(new_n387), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n399), .A2(KEYINPUT72), .A3(G146), .ZN(new_n407));
  INV_X1    g221(.A(G125), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G140), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n390), .A2(new_n409), .A3(new_n247), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n403), .A2(new_n406), .A3(new_n407), .A4(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n401), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(KEYINPUT22), .B(G137), .ZN(new_n413));
  INV_X1    g227(.A(G234), .ZN(new_n414));
  NOR3_X1   g228(.A1(new_n187), .A2(new_n414), .A3(G953), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n413), .B(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n416), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n401), .A2(new_n411), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(new_n189), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT25), .ZN(new_n421));
  INV_X1    g235(.A(G217), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n422), .B1(G234), .B2(new_n189), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT25), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n417), .A2(new_n424), .A3(new_n189), .A4(new_n419), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n421), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  OR2_X1    g240(.A1(new_n420), .A2(new_n423), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n377), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(G113), .B(G122), .ZN(new_n432));
  XNOR2_X1  g246(.A(KEYINPUT85), .B(G104), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n432), .B(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n335), .A2(new_n336), .A3(G214), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(new_n245), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(G131), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n435), .B(G143), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n239), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n395), .A2(KEYINPUT19), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n390), .A2(new_n409), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n441), .B(new_n247), .C1(KEYINPUT19), .C2(new_n442), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n440), .A2(new_n403), .A3(new_n407), .A4(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT18), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n438), .B1(new_n445), .B2(new_n239), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n410), .B1(new_n398), .B2(new_n247), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n446), .B(new_n447), .C1(new_n445), .C2(new_n437), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n444), .A2(KEYINPUT84), .A3(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(KEYINPUT84), .B1(new_n444), .B2(new_n448), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n434), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n397), .A2(new_n400), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n436), .A2(KEYINPUT17), .A3(G131), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n453), .B(new_n454), .C1(KEYINPUT17), .C2(new_n440), .ZN(new_n455));
  INV_X1    g269(.A(new_n434), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(new_n456), .A3(new_n448), .ZN(new_n457));
  AOI21_X1  g271(.A(G475), .B1(new_n452), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT20), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n459), .A3(new_n189), .ZN(new_n460));
  INV_X1    g274(.A(G475), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n444), .A2(new_n448), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT84), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n456), .B1(new_n464), .B2(new_n449), .ZN(new_n465));
  INV_X1    g279(.A(new_n457), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n461), .B(new_n189), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT20), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n460), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n455), .A2(new_n448), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n434), .A2(KEYINPUT87), .ZN(new_n471));
  OR2_X1    g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n471), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n189), .A3(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT86), .B(G475), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n469), .A2(new_n476), .ZN(new_n477));
  OR2_X1    g291(.A1(KEYINPUT92), .A2(G952), .ZN(new_n478));
  NAND2_X1  g292(.A1(KEYINPUT92), .A2(G952), .ZN(new_n479));
  AOI21_X1  g293(.A(G953), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n480), .B1(new_n414), .B2(new_n335), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  XOR2_X1   g296(.A(KEYINPUT21), .B(G898), .Z(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  AOI211_X1 g298(.A(new_n189), .B(new_n336), .C1(G234), .C2(G237), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G478), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n487), .A2(KEYINPUT15), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT14), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(new_n318), .A3(G122), .ZN(new_n490));
  XOR2_X1   g304(.A(new_n490), .B(KEYINPUT90), .Z(new_n491));
  NAND2_X1  g305(.A1(new_n318), .A2(G122), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT14), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT89), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(G122), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(G116), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n492), .A2(KEYINPUT89), .A3(KEYINPUT14), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n495), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(G107), .B1(new_n491), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n497), .A2(new_n492), .A3(new_n193), .ZN(new_n501));
  XOR2_X1   g315(.A(G128), .B(G143), .Z(new_n502));
  OR2_X1    g316(.A1(new_n502), .A2(G134), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(G134), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n500), .A2(new_n501), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT13), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(new_n245), .A3(G128), .ZN(new_n508));
  OAI211_X1 g322(.A(G134), .B(new_n508), .C1(new_n502), .C2(new_n507), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n497), .A2(new_n492), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(G107), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n501), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(new_n503), .A3(new_n512), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n513), .A2(KEYINPUT88), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n513), .A2(KEYINPUT88), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n506), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n188), .ZN(new_n517));
  NOR3_X1   g331(.A1(new_n517), .A2(new_n422), .A3(G953), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n506), .B(new_n518), .C1(new_n514), .C2(new_n515), .ZN(new_n521));
  AOI21_X1  g335(.A(G902), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT91), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI211_X1 g338(.A(KEYINPUT91), .B(G902), .C1(new_n520), .C2(new_n521), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n488), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI22_X1  g340(.A1(new_n522), .A2(new_n523), .B1(KEYINPUT15), .B2(new_n487), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NOR3_X1   g342(.A1(new_n477), .A2(new_n486), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(G214), .B1(G237), .B2(G902), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT6), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n202), .A2(new_n212), .A3(KEYINPUT4), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n218), .A2(new_n216), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n322), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n317), .A2(new_n319), .A3(KEYINPUT5), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n536), .B(G113), .C1(KEYINPUT5), .C2(new_n317), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n320), .A2(new_n321), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI211_X1 g353(.A(new_n243), .B(new_n539), .C1(new_n202), .C2(new_n212), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n535), .A2(new_n541), .ZN(new_n542));
  XOR2_X1   g356(.A(G110), .B(G122), .Z(new_n543));
  AOI21_X1  g357(.A(new_n532), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT79), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n540), .B1(new_n322), .B2(new_n219), .ZN(new_n546));
  INV_X1    g360(.A(new_n543), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AND2_X1   g362(.A1(new_n218), .A2(new_n216), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n342), .B1(new_n549), .B2(new_n213), .ZN(new_n550));
  NOR4_X1   g364(.A1(new_n550), .A2(new_n540), .A3(KEYINPUT79), .A4(new_n543), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n544), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT80), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n283), .A2(new_n408), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n227), .A2(G125), .A3(new_n228), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n336), .A2(G224), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n557), .B(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n542), .A2(new_n532), .A3(new_n543), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n544), .B(KEYINPUT80), .C1(new_n548), .C2(new_n551), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n554), .A2(new_n559), .A3(new_n560), .A4(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n551), .ZN(new_n563));
  OAI21_X1  g377(.A(KEYINPUT79), .B1(new_n542), .B2(new_n543), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n263), .A2(KEYINPUT82), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(new_n539), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n543), .B(KEYINPUT81), .ZN(new_n567));
  XOR2_X1   g381(.A(new_n567), .B(KEYINPUT8), .Z(new_n568));
  AOI22_X1  g382(.A1(new_n563), .A2(new_n564), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n558), .A2(KEYINPUT7), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT83), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n556), .B1(new_n555), .B2(KEYINPUT83), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n557), .A2(new_n572), .B1(new_n573), .B2(new_n570), .ZN(new_n574));
  AOI21_X1  g388(.A(G902), .B1(new_n569), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n562), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(G210), .B1(G237), .B2(G902), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n562), .A2(new_n577), .A3(new_n575), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n531), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n315), .A2(new_n431), .A3(new_n529), .A4(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT93), .B(G101), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(G3));
  INV_X1    g398(.A(new_n315), .ZN(new_n585));
  NAND2_X1  g399(.A1(KEYINPUT94), .A2(G472), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n370), .A2(new_n189), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n586), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n588), .B1(new_n374), .B2(G902), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n585), .A2(new_n428), .A3(new_n590), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n562), .A2(new_n577), .A3(new_n575), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n577), .B1(new_n562), .B2(new_n575), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n530), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n520), .A2(new_n521), .ZN(new_n595));
  OR2_X1    g409(.A1(new_n595), .A2(KEYINPUT33), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(KEYINPUT33), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(G478), .A3(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n487), .A2(new_n189), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n522), .A2(new_n487), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n598), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n477), .A2(new_n603), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n594), .A2(new_n486), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n591), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(new_n191), .ZN(new_n607));
  XNOR2_X1  g421(.A(KEYINPUT95), .B(KEYINPUT34), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G6));
  XNOR2_X1  g423(.A(new_n486), .B(KEYINPUT96), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n530), .B(new_n610), .C1(new_n592), .C2(new_n593), .ZN(new_n611));
  AOI22_X1  g425(.A1(new_n460), .A2(new_n468), .B1(new_n474), .B2(new_n475), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n528), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n591), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT35), .B(G107), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G9));
  NOR2_X1   g431(.A1(new_n416), .A2(KEYINPUT36), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n412), .B(new_n618), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n619), .B(new_n189), .C1(new_n422), .C2(G234), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n426), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT97), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n426), .A2(KEYINPUT97), .A3(new_n620), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n625), .A2(new_n587), .A3(new_n589), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT98), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n627), .A2(new_n529), .A3(new_n315), .A4(new_n581), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT37), .B(G110), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G12));
  INV_X1    g444(.A(new_n314), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n631), .B1(new_n307), .B2(new_n309), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n362), .A2(new_n372), .A3(new_n376), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n632), .A2(new_n633), .A3(new_n190), .ZN(new_n634));
  INV_X1    g448(.A(new_n485), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n481), .B1(new_n635), .B2(G900), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(KEYINPUT99), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  AND4_X1   g452(.A1(new_n469), .A2(new_n528), .A3(new_n476), .A4(new_n638), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n639), .B(new_n530), .C1(new_n592), .C2(new_n593), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT100), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n579), .A2(new_n580), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT100), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n642), .A2(new_n643), .A3(new_n530), .A4(new_n639), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n634), .A2(new_n625), .A3(new_n641), .A4(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G128), .ZN(G30));
  NAND3_X1  g460(.A1(new_n477), .A2(new_n528), .A3(new_n530), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n637), .B(KEYINPUT39), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n315), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT101), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n647), .B1(new_n652), .B2(KEYINPUT40), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n642), .B(KEYINPUT38), .ZN(new_n654));
  INV_X1    g468(.A(new_n357), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n339), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n345), .A2(new_n330), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n189), .B1(new_n657), .B2(new_n338), .ZN(new_n658));
  OAI21_X1  g472(.A(G472), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n372), .A2(new_n376), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n661), .A2(new_n621), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n650), .B(KEYINPUT101), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT40), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n653), .A2(new_n654), .A3(new_n662), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G143), .ZN(G45));
  OAI211_X1 g481(.A(new_n530), .B(new_n625), .C1(new_n592), .C2(new_n593), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n477), .A2(new_n603), .A3(new_n638), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n634), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G146), .ZN(G48));
  AOI21_X1  g487(.A(new_n305), .B1(new_n304), .B2(new_n189), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(new_n307), .B2(new_n309), .ZN(new_n675));
  INV_X1    g489(.A(new_n190), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n675), .A2(new_n377), .A3(new_n429), .A4(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n605), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT102), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT41), .B(G113), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G15));
  INV_X1    g496(.A(KEYINPUT103), .ZN(new_n683));
  AOI211_X1 g497(.A(new_n190), .B(new_n674), .C1(new_n307), .C2(new_n309), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n614), .A2(new_n683), .A3(new_n431), .A4(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n613), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n642), .A2(new_n530), .A3(new_n686), .A4(new_n610), .ZN(new_n687));
  OAI21_X1  g501(.A(KEYINPUT103), .B1(new_n677), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G116), .ZN(G18));
  INV_X1    g504(.A(new_n529), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n668), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT104), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n692), .A2(new_n693), .A3(new_n377), .A4(new_n684), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n642), .A2(new_n529), .A3(new_n530), .A4(new_n625), .ZN(new_n695));
  INV_X1    g509(.A(new_n674), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n310), .A2(new_n377), .A3(new_n676), .A4(new_n696), .ZN(new_n697));
  OAI21_X1  g511(.A(KEYINPUT104), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G119), .ZN(G21));
  AND3_X1   g514(.A1(new_n675), .A2(new_n676), .A3(new_n610), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n592), .A2(new_n593), .ZN(new_n702));
  OR2_X1    g516(.A1(new_n347), .A2(new_n350), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n338), .B1(new_n703), .B2(new_n331), .ZN(new_n704));
  INV_X1    g518(.A(new_n367), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n371), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n428), .B(KEYINPUT105), .ZN(new_n707));
  OAI21_X1  g521(.A(G472), .B1(new_n374), .B2(G902), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n702), .A2(new_n709), .A3(new_n647), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n701), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G122), .ZN(G24));
  NAND2_X1  g526(.A1(new_n706), .A2(new_n708), .ZN(new_n713));
  INV_X1    g527(.A(new_n621), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n713), .A2(new_n714), .A3(new_n670), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n715), .A2(new_n684), .A3(new_n581), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G125), .ZN(G27));
  NOR3_X1   g531(.A1(new_n642), .A2(new_n531), .A3(new_n670), .ZN(new_n718));
  INV_X1    g532(.A(new_n707), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n633), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n718), .A2(KEYINPUT42), .A3(new_n315), .A4(new_n720), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n592), .A2(new_n593), .A3(new_n531), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n315), .A2(new_n431), .A3(new_n671), .A4(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT42), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n723), .A2(KEYINPUT106), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(KEYINPUT106), .B1(new_n723), .B2(new_n724), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n721), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G131), .ZN(G33));
  NAND4_X1  g542(.A1(new_n315), .A2(new_n431), .A3(new_n639), .A4(new_n722), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G134), .ZN(G36));
  NOR3_X1   g544(.A1(new_n477), .A2(KEYINPUT43), .A3(new_n602), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n612), .B(KEYINPUT107), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n603), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n731), .B1(new_n733), .B2(KEYINPUT43), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n590), .A2(new_n621), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n735), .A2(KEYINPUT108), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(KEYINPUT108), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n734), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT44), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n311), .A2(new_n312), .ZN(new_n741));
  XOR2_X1   g555(.A(new_n741), .B(KEYINPUT45), .Z(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(G469), .ZN(new_n743));
  NAND2_X1  g557(.A1(G469), .A2(G902), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(KEYINPUT46), .A3(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT46), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n746), .B(G469), .C1(new_n742), .C2(G902), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n745), .A2(new_n310), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n676), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n749), .A2(new_n648), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n734), .B(KEYINPUT44), .C1(new_n736), .C2(new_n737), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n740), .A2(new_n750), .A3(new_n722), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G137), .ZN(G39));
  INV_X1    g567(.A(KEYINPUT47), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n748), .A2(KEYINPUT47), .A3(new_n676), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n757), .A2(new_n633), .A3(new_n428), .A4(new_n718), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(KEYINPUT109), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G140), .ZN(G42));
  INV_X1    g574(.A(new_n722), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n675), .A2(new_n676), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n428), .A2(new_n481), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n763), .A2(new_n661), .A3(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n480), .B1(new_n766), .B2(new_n604), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n734), .A2(new_n482), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n768), .A2(new_n762), .A3(new_n761), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n720), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT48), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT115), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT114), .ZN(new_n773));
  OR3_X1    g587(.A1(new_n770), .A2(new_n773), .A3(KEYINPUT48), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n773), .B1(new_n770), .B2(KEYINPUT48), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n767), .B1(new_n772), .B2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n684), .A2(new_n531), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n654), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(KEYINPUT112), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT112), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n654), .A2(new_n779), .A3(new_n782), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n768), .A2(new_n709), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT50), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(KEYINPUT113), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n786), .A2(KEYINPUT113), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n784), .A2(new_n785), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n785), .B1(new_n781), .B2(new_n783), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n787), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n675), .A2(new_n190), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n722), .B(new_n785), .C1(new_n757), .C2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n765), .A2(new_n612), .A3(new_n602), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n790), .A2(new_n792), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n713), .A2(new_n714), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n769), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n778), .B1(new_n796), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n777), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n678), .A2(new_n605), .B1(new_n701), .B2(new_n710), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n689), .A2(new_n699), .A3(new_n803), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n604), .A2(new_n613), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n611), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n590), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n806), .A2(new_n429), .A3(new_n315), .A4(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n628), .A2(new_n808), .A3(new_n582), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n477), .A2(new_n528), .A3(new_n637), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n810), .A2(new_n377), .A3(new_n625), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n315), .B(new_n722), .C1(new_n715), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n729), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n804), .A2(new_n727), .A3(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n702), .A2(new_n647), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n816), .A2(new_n315), .A3(new_n662), .A4(new_n638), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n645), .A2(new_n672), .A3(new_n716), .A4(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT52), .ZN(new_n819));
  NOR4_X1   g633(.A1(new_n632), .A2(new_n633), .A3(new_n190), .A4(new_n670), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n581), .A2(new_n676), .A3(new_n675), .ZN(new_n821));
  AOI22_X1  g635(.A1(new_n669), .A2(new_n820), .B1(new_n821), .B2(new_n715), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n822), .A2(new_n823), .A3(new_n645), .A4(new_n817), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n819), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n802), .B1(new_n815), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n819), .A2(new_n824), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n689), .A2(new_n699), .A3(new_n803), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n594), .A2(new_n632), .A3(new_n190), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n830), .B(new_n529), .C1(new_n431), .C2(new_n627), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n729), .A3(new_n812), .A4(new_n808), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n827), .A2(new_n828), .A3(new_n727), .A4(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT54), .B1(new_n826), .B2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n833), .A2(new_n727), .A3(new_n819), .A4(new_n824), .ZN(new_n836));
  INV_X1    g650(.A(new_n802), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT111), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n828), .ZN(new_n839));
  INV_X1    g653(.A(new_n721), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n723), .A2(new_n724), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT106), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n723), .A2(KEYINPUT106), .A3(new_n724), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n840), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n845), .A2(new_n832), .A3(new_n829), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT111), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n846), .A2(new_n847), .A3(new_n827), .A4(new_n802), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n838), .A2(new_n839), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n835), .B1(new_n849), .B2(KEYINPUT54), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n785), .A2(new_n821), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n792), .A2(new_n794), .A3(new_n795), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n852), .A2(KEYINPUT51), .A3(new_n798), .A4(new_n790), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n801), .A2(new_n850), .A3(new_n851), .A4(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n854), .B1(G952), .B2(G953), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n654), .A2(new_n719), .A3(new_n733), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n660), .A2(new_n190), .A3(new_n531), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n675), .B(KEYINPUT49), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n855), .A2(new_n859), .ZN(G75));
  AOI21_X1  g674(.A(new_n837), .B1(new_n846), .B2(new_n827), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n815), .A2(KEYINPUT53), .A3(new_n825), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n861), .A2(new_n862), .A3(new_n189), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(G210), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT56), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n554), .A2(new_n560), .A3(new_n561), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(new_n559), .ZN(new_n867));
  XNOR2_X1  g681(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n867), .B(new_n868), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n864), .A2(new_n865), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n869), .B1(new_n864), .B2(new_n865), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n336), .A2(G952), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(G51));
  XOR2_X1   g687(.A(new_n744), .B(KEYINPUT57), .Z(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT54), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n876), .B1(new_n861), .B2(new_n862), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n826), .A2(new_n834), .A3(KEYINPUT54), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n304), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT117), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n826), .A2(new_n834), .A3(KEYINPUT54), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n874), .B1(new_n882), .B2(new_n835), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT117), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n883), .A2(new_n884), .A3(new_n304), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT118), .ZN(new_n886));
  INV_X1    g700(.A(new_n743), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n863), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n863), .A2(new_n887), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT118), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n881), .A2(new_n885), .A3(new_n888), .A4(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n872), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n891), .A2(new_n892), .ZN(G54));
  NAND3_X1  g707(.A1(new_n863), .A2(KEYINPUT58), .A3(G475), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n894), .A2(new_n452), .A3(new_n457), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n894), .B1(new_n452), .B2(new_n457), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n895), .A2(new_n896), .A3(new_n872), .ZN(G60));
  AND2_X1   g711(.A1(new_n596), .A2(new_n597), .ZN(new_n898));
  XNOR2_X1  g712(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(new_n599), .ZN(new_n900));
  AOI211_X1 g714(.A(new_n898), .B(new_n900), .C1(new_n877), .C2(new_n878), .ZN(new_n901));
  OR2_X1    g715(.A1(new_n901), .A2(new_n872), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n898), .B1(new_n850), .B2(new_n900), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT120), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI211_X1 g719(.A(KEYINPUT120), .B(new_n898), .C1(new_n850), .C2(new_n900), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n902), .B1(new_n905), .B2(new_n906), .ZN(G63));
  NAND2_X1  g721(.A1(G217), .A2(G902), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT60), .Z(new_n909));
  NAND3_X1  g723(.A1(new_n826), .A2(new_n834), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n417), .A2(new_n419), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n619), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n912), .B(new_n892), .C1(new_n913), .C2(new_n910), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(KEYINPUT121), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT61), .ZN(G66));
  AOI21_X1  g730(.A(new_n336), .B1(new_n483), .B2(G224), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n829), .A2(new_n809), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n917), .B1(new_n919), .B2(new_n336), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n866), .B1(G898), .B2(new_n336), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n920), .B(new_n921), .Z(G69));
  NOR2_X1   g736(.A1(new_n353), .A2(new_n354), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n441), .B1(KEYINPUT19), .B2(new_n442), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n923), .B(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(G900), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n926), .A2(KEYINPUT126), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(KEYINPUT126), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n927), .A2(G953), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n727), .A2(new_n729), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT125), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n822), .A2(new_n645), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n750), .A2(new_n816), .A3(new_n720), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n752), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n931), .A2(new_n759), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n929), .B1(new_n935), .B2(G953), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n277), .A2(new_n926), .A3(new_n336), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n925), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n666), .A2(new_n932), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT62), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n315), .A2(new_n431), .A3(new_n649), .A4(new_n722), .ZN(new_n942));
  OR3_X1    g756(.A1(new_n942), .A2(KEYINPUT122), .A3(new_n805), .ZN(new_n943));
  OAI21_X1  g757(.A(KEYINPUT122), .B1(new_n942), .B2(new_n805), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n752), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT123), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n752), .A2(new_n943), .A3(KEYINPUT123), .A4(new_n944), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n941), .A2(KEYINPUT124), .A3(new_n759), .A4(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n939), .A2(new_n940), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT62), .B1(new_n666), .B2(new_n932), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n949), .B(new_n759), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT124), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n950), .A2(new_n955), .A3(new_n336), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n925), .A2(new_n937), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n938), .B1(new_n956), .B2(new_n957), .ZN(G72));
  NAND2_X1  g772(.A1(G472), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT63), .Z(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(new_n935), .B2(new_n919), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n961), .A2(new_n339), .A3(new_n655), .ZN(new_n962));
  INV_X1    g776(.A(new_n363), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n358), .B(KEYINPUT127), .Z(new_n964));
  OAI211_X1 g778(.A(new_n849), .B(new_n960), .C1(new_n963), .C2(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n962), .A2(new_n892), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n950), .A2(new_n955), .A3(new_n918), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n960), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n966), .B1(new_n968), .B2(new_n656), .ZN(G57));
endmodule


