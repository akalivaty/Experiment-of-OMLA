//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1303, new_n1304, new_n1305, new_n1306,
    new_n1307, new_n1308, new_n1309, new_n1310, new_n1311, new_n1312,
    new_n1313, new_n1314, new_n1315, new_n1316, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1328, new_n1329, new_n1330, new_n1331,
    new_n1332, new_n1333, new_n1334, new_n1335, new_n1336, new_n1337,
    new_n1338, new_n1339, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1346, new_n1347, new_n1348, new_n1349, new_n1350, new_n1351,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1411, new_n1412, new_n1413,
    new_n1414, new_n1415, new_n1416, new_n1417, new_n1418, new_n1419,
    new_n1420, new_n1421, new_n1422;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n202), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT65), .B(G244), .ZN(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT64), .B(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  OAI22_X1  g0020(.A1(new_n217), .A2(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n208), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT66), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XOR2_X1   g0038(.A(G107), .B(G116), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT67), .ZN(new_n243));
  XOR2_X1   g0043(.A(G58), .B(G77), .Z(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G169), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  AND2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  OAI211_X1 g0050(.A(G257), .B(new_n248), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  OAI211_X1 g0051(.A(G264), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n252));
  INV_X1    g0052(.A(G303), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT3), .B(G33), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n251), .B(new_n252), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G1), .A3(G13), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT5), .B(G41), .ZN(new_n260));
  INV_X1    g0060(.A(G45), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(G1), .ZN(new_n262));
  AND2_X1   g0062(.A1(G1), .A2(G13), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n260), .A2(new_n262), .B1(new_n263), .B2(new_n256), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n205), .A2(G45), .ZN(new_n265));
  OR2_X1    g0065(.A1(KEYINPUT5), .A2(G41), .ZN(new_n266));
  NAND2_X1  g0066(.A1(KEYINPUT5), .A2(G41), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G274), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n269), .B1(new_n263), .B2(new_n256), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n264), .A2(G270), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n247), .B1(new_n259), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n214), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G13), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(G1), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G20), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT72), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n275), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NOR3_X1   g0080(.A1(new_n276), .A2(new_n206), .A3(G1), .ZN(new_n281));
  OAI21_X1  g0081(.A(KEYINPUT72), .B1(new_n281), .B2(new_n274), .ZN(new_n282));
  INV_X1    g0082(.A(G116), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n283), .B1(new_n205), .B2(G33), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n280), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n277), .A2(G20), .A3(new_n283), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n273), .A2(new_n214), .B1(G20), .B2(new_n283), .ZN(new_n287));
  NAND2_X1  g0087(.A1(G33), .A2(G283), .ZN(new_n288));
  INV_X1    g0088(.A(G97), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n288), .B(new_n206), .C1(G33), .C2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(KEYINPUT20), .B1(new_n287), .B2(new_n290), .ZN(new_n291));
  AND3_X1   g0091(.A1(new_n287), .A2(KEYINPUT20), .A3(new_n290), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n285), .B(new_n286), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n272), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT21), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT21), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n272), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n259), .A2(new_n271), .ZN(new_n298));
  INV_X1    g0098(.A(G179), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n295), .A2(new_n297), .B1(new_n293), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT83), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n298), .A2(G200), .ZN(new_n303));
  INV_X1    g0103(.A(new_n293), .ZN(new_n304));
  INV_X1    g0104(.A(G190), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n303), .B(new_n304), .C1(new_n305), .C2(new_n298), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n301), .A2(new_n302), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n300), .A2(new_n293), .ZN(new_n308));
  INV_X1    g0108(.A(new_n297), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n296), .B1(new_n272), .B2(new_n293), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n306), .B(new_n308), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT83), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n254), .A2(G1698), .ZN(new_n314));
  INV_X1    g0114(.A(G223), .ZN(new_n315));
  OAI22_X1  g0115(.A1(new_n314), .A2(new_n315), .B1(new_n217), .B2(new_n254), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n254), .A2(G222), .A3(new_n248), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT69), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n254), .A2(KEYINPUT69), .A3(G222), .A4(new_n248), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n257), .B1(new_n317), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G41), .ZN(new_n324));
  AOI21_X1  g0124(.A(G1), .B1(new_n324), .B2(new_n261), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n325), .A2(new_n257), .A3(G274), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n261), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n205), .A2(new_n327), .B1(new_n263), .B2(new_n256), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G226), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n326), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n247), .B1(new_n323), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n205), .A2(G20), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n275), .A2(new_n333), .ZN(new_n334));
  MUX2_X1   g0134(.A(new_n278), .B(new_n334), .S(G50), .Z(new_n335));
  OAI21_X1  g0135(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n336));
  INV_X1    g0136(.A(G150), .ZN(new_n337));
  NOR2_X1   g0137(.A1(G20), .A2(G33), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n336), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT8), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G58), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n342), .B(KEYINPUT71), .ZN(new_n343));
  INV_X1    g0143(.A(G58), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT8), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT70), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n344), .A2(KEYINPUT70), .A3(KEYINPUT8), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n343), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G33), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n350), .A2(G20), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n340), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n335), .B1(new_n352), .B2(new_n275), .ZN(new_n353));
  INV_X1    g0153(.A(new_n331), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n316), .B1(new_n320), .B2(new_n321), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n299), .B(new_n354), .C1(new_n355), .C2(new_n257), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n332), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT74), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT9), .ZN(new_n359));
  AND3_X1   g0159(.A1(new_n353), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n358), .B1(new_n353), .B2(new_n359), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(G200), .B1(new_n323), .B2(new_n331), .ZN(new_n363));
  OAI211_X1 g0163(.A(G190), .B(new_n354), .C1(new_n355), .C2(new_n257), .ZN(new_n364));
  OAI211_X1 g0164(.A(KEYINPUT9), .B(new_n335), .C1(new_n352), .C2(new_n275), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NOR3_X1   g0166(.A1(new_n362), .A2(KEYINPUT10), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT10), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n353), .A2(new_n359), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT74), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n353), .A2(new_n358), .A3(new_n359), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n366), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n368), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n357), .B1(new_n367), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n315), .A2(new_n248), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n330), .A2(G1698), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n376), .B(new_n377), .C1(new_n249), .C2(new_n250), .ZN(new_n378));
  NAND2_X1  g0178(.A1(G33), .A2(G87), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n258), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n257), .A2(G232), .A3(new_n382), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n326), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n381), .A2(new_n384), .A3(G179), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n257), .B1(new_n378), .B2(new_n379), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n326), .A2(new_n383), .ZN(new_n387));
  OAI21_X1  g0187(.A(G169), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AND3_X1   g0188(.A1(new_n385), .A2(KEYINPUT78), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT78), .B1(new_n385), .B2(new_n388), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT18), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT16), .ZN(new_n393));
  INV_X1    g0193(.A(G159), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n339), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G68), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT64), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT64), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G68), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n201), .B1(new_n401), .B2(G58), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n396), .B1(new_n402), .B2(new_n206), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT3), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n350), .ZN(new_n405));
  NAND2_X1  g0205(.A1(KEYINPUT3), .A2(G33), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n206), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT7), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n405), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n406), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n219), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n393), .B1(new_n403), .B2(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n249), .A2(new_n250), .ZN(new_n413));
  AOI21_X1  g0213(.A(KEYINPUT7), .B1(new_n413), .B2(new_n206), .ZN(new_n414));
  INV_X1    g0214(.A(new_n410), .ZN(new_n415));
  OAI21_X1  g0215(.A(G68), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n202), .B1(new_n219), .B2(new_n344), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n395), .B1(new_n417), .B2(G20), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n416), .A2(new_n418), .A3(KEYINPUT16), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n412), .A2(new_n419), .A3(new_n274), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n349), .A2(new_n334), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n343), .A2(new_n278), .A3(new_n347), .A4(new_n348), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n391), .A2(new_n392), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n392), .B1(new_n391), .B2(new_n424), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(G200), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(new_n381), .B2(new_n384), .ZN(new_n430));
  NOR3_X1   g0230(.A1(new_n386), .A2(new_n387), .A3(new_n305), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n420), .A2(new_n423), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT17), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n420), .A2(KEYINPUT17), .A3(new_n423), .A4(new_n432), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(G20), .A2(G77), .ZN(new_n438));
  XNOR2_X1  g0238(.A(KEYINPUT15), .B(G87), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n206), .A2(G33), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n342), .A2(new_n345), .ZN(new_n441));
  OAI221_X1 g0241(.A(new_n438), .B1(new_n439), .B2(new_n440), .C1(new_n441), .C2(new_n339), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n274), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n280), .A2(new_n282), .A3(G77), .A4(new_n333), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n281), .A2(new_n217), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT73), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n442), .A2(new_n274), .B1(new_n217), .B2(new_n281), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT73), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(new_n449), .A3(new_n444), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(G232), .A2(G1698), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n248), .A2(G238), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n254), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n454), .B(new_n258), .C1(G107), .C2(new_n254), .ZN(new_n455));
  INV_X1    g0255(.A(new_n218), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n328), .A2(new_n456), .B1(new_n270), .B2(new_n325), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(G179), .ZN(new_n459));
  AOI21_X1  g0259(.A(G169), .B1(new_n455), .B2(new_n457), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n451), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n458), .A2(G200), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n455), .A2(G190), .A3(new_n457), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n447), .A2(new_n450), .A3(new_n463), .A4(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n428), .A2(new_n437), .A3(new_n462), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n219), .A2(G20), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n351), .A2(G77), .B1(new_n338), .B2(G50), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n275), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  XOR2_X1   g0269(.A(new_n469), .B(KEYINPUT11), .Z(new_n470));
  NAND4_X1  g0270(.A1(new_n280), .A2(new_n282), .A3(G68), .A4(new_n333), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT12), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n205), .A2(G13), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n467), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT12), .B1(new_n281), .B2(new_n397), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n470), .A2(new_n471), .A3(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n326), .B1(new_n329), .B2(new_n220), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT13), .ZN(new_n480));
  OAI211_X1 g0280(.A(G226), .B(new_n248), .C1(new_n249), .C2(new_n250), .ZN(new_n481));
  NAND2_X1  g0281(.A1(G33), .A2(G97), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g0283(.A(G232), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT75), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n254), .A2(KEYINPUT75), .A3(G232), .A4(G1698), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n483), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n479), .B(new_n480), .C1(new_n257), .C2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT76), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n486), .A2(new_n487), .ZN(new_n491));
  INV_X1    g0291(.A(new_n483), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n257), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT13), .B1(new_n493), .B2(new_n478), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n491), .A2(new_n492), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n258), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT76), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n496), .A2(new_n497), .A3(new_n480), .A4(new_n479), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n490), .A2(new_n494), .A3(G179), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n494), .A2(new_n489), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT77), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT14), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n500), .A2(G169), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n502), .B1(new_n500), .B2(G169), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n477), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n490), .A2(new_n494), .A3(G190), .A4(new_n498), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n500), .A2(G200), .ZN(new_n508));
  INV_X1    g0308(.A(new_n477), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n375), .A2(new_n466), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G294), .ZN(new_n513));
  INV_X1    g0313(.A(G257), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G1698), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(G250), .B2(G1698), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n513), .B1(new_n516), .B2(new_n413), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n258), .A2(new_n517), .B1(new_n264), .B2(G264), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT84), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n268), .A2(new_n270), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n267), .ZN(new_n522));
  NOR2_X1   g0322(.A1(KEYINPUT5), .A2(G41), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n262), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n524), .A2(G264), .A3(new_n257), .ZN(new_n525));
  NOR2_X1   g0325(.A1(G250), .A2(G1698), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n526), .B1(new_n514), .B2(G1698), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n527), .A2(new_n254), .B1(G33), .B2(G294), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n520), .B(new_n525), .C1(new_n528), .C2(new_n257), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(KEYINPUT84), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n521), .A2(new_n530), .A3(G169), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n518), .A2(G179), .A3(new_n520), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n206), .B(G87), .C1(new_n249), .C2(new_n250), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT22), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT22), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n254), .A2(new_n536), .A3(new_n206), .A4(G87), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT24), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT23), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n206), .B2(G107), .ZN(new_n541));
  INV_X1    g0341(.A(G107), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n542), .A2(KEYINPUT23), .A3(G20), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n350), .A2(new_n283), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n541), .A2(new_n543), .B1(new_n544), .B2(new_n206), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n538), .A2(new_n539), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n539), .B1(new_n538), .B2(new_n545), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n274), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n281), .A2(new_n274), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n205), .A2(G33), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT25), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n278), .B2(G107), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n281), .A2(KEYINPUT25), .A3(new_n542), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n552), .A2(G107), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n548), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n533), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n558), .A2(KEYINPUT85), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT85), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n560), .B1(new_n533), .B2(new_n557), .ZN(new_n561));
  AOI21_X1  g0361(.A(G190), .B1(new_n521), .B2(new_n530), .ZN(new_n562));
  AOI21_X1  g0362(.A(G200), .B1(new_n518), .B2(new_n520), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n564), .A2(new_n557), .ZN(new_n565));
  NOR3_X1   g0365(.A1(new_n559), .A2(new_n561), .A3(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT81), .ZN(new_n567));
  OAI21_X1  g0367(.A(G107), .B1(new_n414), .B2(new_n415), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n339), .A2(new_n217), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT6), .ZN(new_n570));
  AND2_X1   g0370(.A1(G97), .A2(G107), .ZN(new_n571));
  NOR2_X1   g0371(.A1(G97), .A2(G107), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n542), .A2(KEYINPUT6), .A3(G97), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n569), .B1(new_n575), .B2(G20), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n275), .B1(new_n568), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n278), .A2(G97), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n551), .B2(new_n289), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(G244), .B(new_n248), .C1(new_n249), .C2(new_n250), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT4), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n288), .ZN(new_n585));
  NAND2_X1  g0385(.A1(G250), .A2(G1698), .ZN(new_n586));
  NAND2_X1  g0386(.A1(KEYINPUT4), .A2(G244), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n586), .B1(new_n587), .B2(G1698), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n585), .B1(new_n254), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n257), .B1(new_n584), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n524), .A2(G257), .A3(new_n257), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n520), .ZN(new_n592));
  OAI21_X1  g0392(.A(G200), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT79), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT79), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n595), .B(G200), .C1(new_n590), .C2(new_n592), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n590), .A2(new_n592), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G190), .ZN(new_n598));
  AND4_X1   g0398(.A1(new_n581), .A2(new_n594), .A3(new_n596), .A4(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(KEYINPUT80), .B1(new_n577), .B2(new_n580), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n542), .A2(KEYINPUT6), .A3(G97), .ZN(new_n601));
  XNOR2_X1  g0401(.A(G97), .B(G107), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n601), .B1(new_n602), .B2(new_n570), .ZN(new_n603));
  OAI22_X1  g0403(.A1(new_n603), .A2(new_n206), .B1(new_n217), .B2(new_n339), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n542), .B1(new_n409), .B2(new_n410), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n274), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n580), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT80), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(G169), .B1(new_n590), .B2(new_n592), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n584), .A2(new_n589), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n258), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n591), .A2(new_n520), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(G179), .A3(new_n613), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n600), .A2(new_n609), .B1(new_n610), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n567), .B1(new_n599), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n600), .A2(new_n609), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n614), .A2(new_n610), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n581), .A2(new_n594), .A3(new_n596), .A4(new_n598), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(KEYINPUT81), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n220), .A2(new_n248), .ZN(new_n622));
  INV_X1    g0422(.A(G244), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(G1698), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n622), .B(new_n624), .C1(new_n249), .C2(new_n250), .ZN(new_n625));
  INV_X1    g0425(.A(new_n544), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n257), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n257), .A2(G274), .A3(new_n262), .ZN(new_n628));
  INV_X1    g0428(.A(G250), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(new_n205), .B2(G45), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n257), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n247), .B1(new_n627), .B2(new_n632), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n270), .A2(new_n262), .B1(new_n257), .B2(new_n630), .ZN(new_n634));
  NOR2_X1   g0434(.A1(G238), .A2(G1698), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n635), .B1(new_n623), .B2(G1698), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n544), .B1(new_n636), .B2(new_n254), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n634), .B(new_n299), .C1(new_n637), .C2(new_n257), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n206), .ZN(new_n641));
  INV_X1    g0441(.A(G87), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n572), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n206), .B(G68), .C1(new_n249), .C2(new_n250), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT19), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n440), .B2(new_n289), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n644), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n648), .A2(new_n274), .B1(new_n281), .B2(new_n439), .ZN(new_n649));
  INV_X1    g0449(.A(new_n439), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n549), .A2(new_n550), .A3(new_n650), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n649), .A2(KEYINPUT82), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(KEYINPUT82), .B1(new_n649), .B2(new_n651), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n639), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n627), .A2(new_n632), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(G190), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n634), .B1(new_n637), .B2(new_n257), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G200), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n552), .A2(G87), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n656), .A2(new_n658), .A3(new_n649), .A4(new_n659), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n654), .A2(new_n660), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n616), .A2(new_n621), .A3(new_n661), .ZN(new_n662));
  AND4_X1   g0462(.A1(new_n313), .A2(new_n512), .A3(new_n566), .A4(new_n662), .ZN(G372));
  INV_X1    g0463(.A(new_n357), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n385), .A2(new_n388), .ZN(new_n665));
  AOI211_X1 g0465(.A(KEYINPUT18), .B(new_n665), .C1(new_n420), .C2(new_n423), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n385), .A2(new_n388), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n392), .B1(new_n424), .B2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n450), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n449), .B1(new_n448), .B2(new_n444), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n461), .B(KEYINPUT86), .C1(new_n670), .C2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(KEYINPUT86), .B1(new_n451), .B2(new_n461), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n505), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n676), .A2(new_n499), .A3(new_n503), .ZN(new_n677));
  AOI22_X1  g0477(.A1(new_n510), .A2(new_n675), .B1(new_n677), .B2(new_n477), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n435), .A2(new_n436), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n669), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT10), .B1(new_n362), .B2(new_n366), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n372), .A2(new_n368), .A3(new_n373), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n664), .B1(new_n680), .B2(new_n683), .ZN(new_n684));
  AOI22_X1  g0484(.A1(new_n614), .A2(new_n610), .B1(new_n606), .B2(new_n607), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT26), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n654), .A2(new_n660), .A3(new_n685), .A4(new_n686), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n687), .A2(new_n654), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n654), .A2(new_n660), .ZN(new_n689));
  OAI21_X1  g0489(.A(KEYINPUT26), .B1(new_n619), .B2(new_n689), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n548), .B(new_n556), .C1(new_n562), .C2(new_n563), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n661), .A2(new_n691), .A3(new_n619), .A4(new_n620), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n532), .A2(new_n531), .B1(new_n548), .B2(new_n556), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n688), .B(new_n690), .C1(new_n692), .C2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n512), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n684), .A2(new_n697), .ZN(G369));
  INV_X1    g0498(.A(new_n561), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n694), .A2(new_n560), .ZN(new_n700));
  OR3_X1    g0500(.A1(new_n473), .A2(KEYINPUT27), .A3(G20), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT27), .B1(new_n473), .B2(G20), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n701), .A2(G213), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g0503(.A(KEYINPUT87), .B(G343), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT88), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n557), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n699), .A2(new_n700), .A3(new_n691), .A4(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n694), .A2(new_n707), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT89), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n307), .A2(new_n312), .B1(new_n293), .B2(new_n707), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n707), .A2(new_n293), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n301), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(G330), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n713), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI211_X1 g0519(.A(KEYINPUT89), .B(G330), .C1(new_n714), .C2(new_n716), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n712), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n559), .A2(new_n561), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n301), .A2(new_n707), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n722), .A2(new_n691), .A3(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n707), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n694), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n721), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT90), .ZN(G399));
  INV_X1    g0529(.A(new_n209), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(G41), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n643), .A2(G116), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n732), .A2(G1), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(new_n212), .B2(new_n732), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT28), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n692), .B1(new_n722), .B2(new_n301), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n661), .A2(new_n685), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(KEYINPUT26), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n661), .A2(new_n686), .A3(new_n615), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n739), .A2(new_n740), .A3(new_n654), .ZN(new_n741));
  OAI211_X1 g0541(.A(KEYINPUT29), .B(new_n725), .C1(new_n737), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n696), .A2(new_n725), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT29), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n662), .A2(new_n566), .A3(new_n313), .A4(new_n725), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n518), .A2(new_n655), .A3(new_n259), .A4(new_n271), .ZN(new_n748));
  OAI21_X1  g0548(.A(KEYINPUT91), .B1(new_n748), .B2(new_n614), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n590), .A2(new_n592), .A3(new_n299), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n525), .B1(new_n528), .B2(new_n257), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n657), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT91), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n524), .A2(G270), .A3(new_n257), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n520), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n755), .B1(new_n258), .B2(new_n255), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n750), .A2(new_n752), .A3(new_n753), .A4(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT30), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n749), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n750), .A2(new_n752), .A3(KEYINPUT30), .A4(new_n756), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n657), .B(KEYINPUT92), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n756), .A2(new_n597), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n761), .A2(new_n762), .A3(new_n299), .A4(new_n529), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n759), .A2(new_n760), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(KEYINPUT31), .B1(new_n764), .B2(new_n707), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n759), .A2(new_n763), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(KEYINPUT93), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT93), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n759), .A2(new_n768), .A3(new_n763), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n767), .A2(new_n760), .A3(new_n769), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n707), .A2(KEYINPUT31), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n765), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n718), .B1(new_n747), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n746), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n736), .B1(new_n774), .B2(G1), .ZN(G364));
  NOR2_X1   g0575(.A1(new_n276), .A2(G20), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n205), .B1(new_n776), .B2(G45), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n731), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(new_n717), .B2(new_n718), .ZN(new_n780));
  AND3_X1   g0580(.A1(new_n719), .A2(new_n780), .A3(new_n720), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n214), .B1(G20), .B2(new_n247), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n206), .A2(new_n299), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n784), .A2(new_n305), .A3(G200), .ZN(new_n785));
  INV_X1    g0585(.A(new_n784), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n786), .A2(new_n305), .A3(new_n429), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G50), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n254), .B1(new_n397), .B2(new_n785), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT32), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n206), .A2(G179), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G190), .A2(G200), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n791), .B1(new_n794), .B2(new_n394), .ZN(new_n795));
  INV_X1    g0595(.A(new_n794), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n796), .A2(KEYINPUT32), .A3(G159), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n790), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n792), .A2(new_n305), .A3(G200), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n542), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n784), .A2(G190), .A3(new_n429), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n792), .A2(G190), .A3(G200), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n801), .A2(new_n344), .B1(new_n802), .B2(new_n642), .ZN(new_n803));
  NOR3_X1   g0603(.A1(new_n305), .A2(G179), .A3(G200), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n206), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n800), .B(new_n803), .C1(G97), .C2(new_n806), .ZN(new_n807));
  AND3_X1   g0607(.A1(new_n784), .A2(KEYINPUT95), .A3(new_n793), .ZN(new_n808));
  AOI21_X1  g0608(.A(KEYINPUT95), .B1(new_n784), .B2(new_n793), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n810), .A2(KEYINPUT96), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n810), .A2(KEYINPUT96), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n798), .B(new_n807), .C1(new_n217), .C2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n254), .B1(new_n796), .B2(G329), .ZN(new_n815));
  XOR2_X1   g0615(.A(KEYINPUT33), .B(G317), .Z(new_n816));
  OAI21_X1  g0616(.A(new_n815), .B1(new_n785), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n810), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n817), .B1(new_n818), .B2(G311), .ZN(new_n819));
  INV_X1    g0619(.A(G294), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n805), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G322), .ZN(new_n822));
  INV_X1    g0622(.A(G283), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n801), .A2(new_n822), .B1(new_n799), .B2(new_n823), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n821), .B(new_n824), .C1(G326), .C2(new_n787), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n802), .B(KEYINPUT97), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n819), .B(new_n825), .C1(new_n253), .C2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n783), .B1(new_n814), .B2(new_n828), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n779), .B(KEYINPUT94), .Z(new_n830));
  NOR2_X1   g0630(.A1(new_n730), .A2(new_n413), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(G355), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(G116), .B2(new_n209), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n245), .A2(new_n261), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n730), .A2(new_n254), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(new_n261), .B2(new_n213), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n833), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(G13), .A2(G33), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(G20), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n841), .A2(new_n782), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n830), .B1(new_n838), .B2(new_n843), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n829), .B(new_n844), .C1(new_n717), .C2(new_n841), .ZN(new_n845));
  OR2_X1    g0645(.A1(new_n781), .A2(new_n845), .ZN(G396));
  INV_X1    g0646(.A(KEYINPUT86), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n462), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n707), .B1(new_n670), .B2(new_n671), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n848), .A2(new_n850), .A3(new_n672), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n462), .A2(new_n849), .A3(new_n465), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n696), .A2(new_n725), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(KEYINPUT100), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT100), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n696), .A2(new_n856), .A3(new_n853), .A4(new_n725), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n687), .A2(new_n654), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n661), .A2(new_n615), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n859), .B1(KEYINPUT26), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n301), .A2(new_n558), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n599), .A2(new_n615), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n862), .A2(new_n863), .A3(new_n691), .A4(new_n661), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n707), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n858), .B1(new_n865), .B2(new_n853), .ZN(new_n866));
  INV_X1    g0666(.A(new_n773), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n779), .B1(new_n866), .B2(new_n867), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n462), .A2(new_n849), .A3(new_n465), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n675), .B2(new_n850), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n839), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n783), .A2(new_n840), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n830), .B1(G77), .B2(new_n874), .ZN(new_n875));
  XOR2_X1   g0675(.A(new_n875), .B(KEYINPUT98), .Z(new_n876));
  INV_X1    g0676(.A(G311), .ZN(new_n877));
  OAI22_X1  g0677(.A1(new_n785), .A2(new_n823), .B1(new_n794), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n801), .ZN(new_n879));
  INV_X1    g0679(.A(new_n799), .ZN(new_n880));
  AOI22_X1  g0680(.A1(G294), .A2(new_n879), .B1(new_n880), .B2(G87), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n253), .B2(new_n788), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n878), .B(new_n882), .C1(G97), .C2(new_n806), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n254), .B1(new_n826), .B2(G107), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n884), .B(KEYINPUT99), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n883), .B(new_n885), .C1(new_n283), .C2(new_n813), .ZN(new_n886));
  INV_X1    g0686(.A(new_n785), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n787), .A2(G137), .B1(new_n887), .B2(G150), .ZN(new_n888));
  INV_X1    g0688(.A(G143), .ZN(new_n889));
  OAI221_X1 g0689(.A(new_n888), .B1(new_n889), .B2(new_n801), .C1(new_n813), .C2(new_n394), .ZN(new_n890));
  XOR2_X1   g0690(.A(new_n890), .B(KEYINPUT34), .Z(new_n891));
  NOR2_X1   g0691(.A1(new_n799), .A2(new_n397), .ZN(new_n892));
  INV_X1    g0692(.A(G132), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n254), .B1(new_n794), .B2(new_n893), .ZN(new_n894));
  AOI211_X1 g0694(.A(new_n892), .B(new_n894), .C1(G58), .C2(new_n806), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(new_n789), .B2(new_n827), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n886), .B1(new_n891), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n876), .B1(new_n897), .B2(new_n782), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n869), .A2(new_n870), .B1(new_n873), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(G384));
  NOR2_X1   g0700(.A1(new_n776), .A2(new_n205), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n397), .B1(new_n409), .B2(new_n410), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n393), .B1(new_n403), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(new_n419), .A3(new_n274), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n423), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n703), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT101), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT101), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n905), .A2(new_n908), .A3(new_n703), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n421), .A2(new_n422), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n403), .A2(new_n902), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n275), .B1(new_n912), .B2(KEYINPUT16), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n911), .B1(new_n913), .B2(new_n412), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT78), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n667), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n385), .A2(KEYINPUT78), .A3(new_n388), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(KEYINPUT18), .B1(new_n914), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n425), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n910), .B1(new_n920), .B2(new_n679), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT37), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n908), .B1(new_n905), .B2(new_n703), .ZN(new_n923));
  INV_X1    g0723(.A(new_n703), .ZN(new_n924));
  AOI211_X1 g0724(.A(KEYINPUT101), .B(new_n924), .C1(new_n904), .C2(new_n423), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n905), .A2(new_n667), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n927), .A2(new_n433), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n922), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT37), .B1(new_n391), .B2(new_n424), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n424), .A2(new_n703), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n930), .A2(new_n433), .A3(new_n931), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n921), .B(KEYINPUT38), .C1(new_n929), .C2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT38), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n931), .B1(new_n669), .B2(new_n437), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n424), .A2(new_n667), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n936), .A2(new_n931), .A3(new_n433), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n420), .A2(new_n423), .A3(new_n432), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n924), .B1(new_n420), .B2(new_n423), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n937), .A2(KEYINPUT37), .B1(new_n940), .B2(new_n930), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n934), .B1(new_n935), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n933), .A2(new_n942), .ZN(new_n943));
  OR2_X1    g0743(.A1(KEYINPUT103), .A2(KEYINPUT31), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n764), .A2(new_n707), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n944), .B1(new_n764), .B2(new_n707), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n747), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n510), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n477), .B(new_n707), .C1(new_n677), .C2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n477), .A2(new_n707), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n506), .A2(new_n510), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n872), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n943), .A2(new_n948), .A3(KEYINPUT40), .A4(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT104), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT40), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n933), .B2(new_n942), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n958), .A2(KEYINPUT104), .A3(new_n953), .A4(new_n948), .ZN(new_n959));
  INV_X1    g0759(.A(new_n933), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n940), .A2(new_n930), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n927), .A2(new_n433), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n962), .A2(new_n925), .A3(new_n923), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n961), .B1(new_n963), .B2(new_n922), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT38), .B1(new_n964), .B2(new_n921), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n953), .B(new_n948), .C1(new_n960), .C2(new_n965), .ZN(new_n966));
  XOR2_X1   g0766(.A(KEYINPUT102), .B(KEYINPUT40), .Z(new_n967));
  AOI22_X1  g0767(.A1(new_n956), .A2(new_n959), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n512), .A2(new_n948), .ZN(new_n969));
  OAI21_X1  g0769(.A(G330), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT105), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n968), .A2(new_n969), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(new_n971), .B2(new_n970), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n950), .A2(new_n952), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n462), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n725), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n978), .B1(new_n858), .B2(new_n980), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n907), .A2(new_n433), .A3(new_n909), .A4(new_n927), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n932), .B1(KEYINPUT37), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n926), .B1(new_n428), .B2(new_n437), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n934), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n933), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n981), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n924), .B1(new_n666), .B2(new_n668), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n677), .A2(new_n477), .A3(new_n725), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT39), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n943), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n985), .A2(KEYINPUT39), .A3(new_n933), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n987), .B(new_n988), .C1(new_n989), .C2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n746), .A2(new_n512), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n684), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n994), .B(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n901), .B1(new_n976), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n997), .B2(new_n976), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n575), .A2(KEYINPUT35), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n575), .A2(KEYINPUT35), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n1000), .A2(new_n1001), .A3(G116), .A4(new_n215), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT36), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n213), .B(G77), .C1(new_n344), .C2(new_n219), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(G50), .B2(new_n397), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1005), .A2(G1), .A3(new_n276), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n999), .A2(new_n1003), .A3(new_n1006), .ZN(G367));
  NAND2_X1  g0807(.A1(new_n659), .A2(new_n649), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n707), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n661), .A2(new_n1009), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1010), .A2(KEYINPUT106), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(KEYINPUT106), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1011), .B(new_n1012), .C1(new_n654), .C2(new_n1009), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1013), .A2(KEYINPUT107), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(KEYINPUT107), .ZN(new_n1015));
  XOR2_X1   g0815(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n1016));
  NAND3_X1  g0816(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n619), .B(new_n620), .C1(new_n581), .C2(new_n725), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n685), .A2(new_n707), .ZN(new_n1019));
  AND3_X1   g0819(.A1(new_n1018), .A2(KEYINPUT109), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(KEYINPUT109), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n721), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1024));
  OAI21_X1  g0824(.A(KEYINPUT42), .B1(new_n1024), .B2(new_n724), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT42), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1022), .A2(new_n1026), .A3(new_n566), .A4(new_n723), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n699), .A2(new_n700), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n615), .B1(new_n1022), .B2(new_n1028), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1025), .B(new_n1027), .C1(new_n1029), .C2(new_n707), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1013), .A2(KEYINPUT43), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1023), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1023), .B1(new_n1031), .B2(new_n1030), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1017), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1036), .A2(new_n721), .A3(new_n1022), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1017), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1037), .A2(new_n1038), .A3(new_n1032), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1035), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n731), .B(KEYINPUT41), .Z(new_n1042));
  OR2_X1    g0842(.A1(new_n711), .A2(new_n723), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n724), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n719), .A2(new_n720), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT110), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1044), .A2(KEYINPUT110), .A3(new_n719), .A4(new_n720), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1048), .A2(new_n774), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n721), .A2(KEYINPUT111), .ZN(new_n1052));
  AND2_X1   g0852(.A1(new_n724), .A2(new_n726), .ZN(new_n1053));
  AOI21_X1  g0853(.A(KEYINPUT45), .B1(new_n1053), .B2(new_n1022), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT45), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n727), .A2(new_n1024), .A3(new_n1055), .ZN(new_n1056));
  AND3_X1   g0856(.A1(new_n727), .A2(new_n1024), .A3(KEYINPUT44), .ZN(new_n1057));
  AOI21_X1  g0857(.A(KEYINPUT44), .B1(new_n727), .B2(new_n1024), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n1054), .A2(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT111), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n1060), .B(new_n712), .C1(new_n719), .C2(new_n720), .ZN(new_n1061));
  NOR3_X1   g0861(.A1(new_n1052), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1058), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n727), .A2(new_n1024), .A3(KEYINPUT44), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1053), .A2(new_n1022), .A3(KEYINPUT45), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1055), .B1(new_n727), .B2(new_n1024), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1063), .A2(new_n1064), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NOR3_X1   g0867(.A1(new_n1067), .A2(KEYINPUT111), .A3(new_n721), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1051), .B1(new_n1062), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1042), .B1(new_n1069), .B2(new_n774), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1041), .B1(new_n1070), .B2(new_n778), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n842), .B1(new_n209), .B2(new_n439), .C1(new_n836), .C2(new_n236), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n830), .A2(new_n1072), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n802), .A2(KEYINPUT46), .A3(new_n283), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n826), .A2(G116), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1074), .B1(new_n1075), .B2(KEYINPUT46), .ZN(new_n1076));
  INV_X1    g0876(.A(G317), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n413), .B1(new_n794), .B2(new_n1077), .C1(new_n785), .C2(new_n820), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n788), .A2(new_n877), .B1(new_n542), .B2(new_n805), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n801), .A2(new_n253), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n799), .A2(new_n289), .ZN(new_n1081));
  OR4_X1    g0881(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .A4(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n813), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1076), .B(new_n1082), .C1(G283), .C2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(G137), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n254), .B1(new_n794), .B2(new_n1085), .C1(new_n785), .C2(new_n394), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n344), .A2(new_n802), .B1(new_n799), .B2(new_n217), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n1086), .B(new_n1087), .C1(new_n1083), .C2(G50), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n801), .A2(new_n337), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n805), .A2(new_n397), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n1089), .B(new_n1090), .C1(G143), .C2(new_n787), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT112), .Z(new_n1092));
  AOI21_X1  g0892(.A(new_n1084), .B1(new_n1088), .B2(new_n1092), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT47), .Z(new_n1094));
  AOI21_X1  g0894(.A(new_n1073), .B1(new_n1094), .B2(new_n782), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n841), .ZN(new_n1096));
  OR2_X1    g0896(.A1(new_n1013), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1071), .A2(new_n1098), .ZN(G387));
  NAND2_X1  g0899(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n774), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1102), .A2(new_n731), .A3(new_n1050), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n805), .A2(new_n439), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n788), .A2(new_n394), .B1(new_n802), .B2(new_n217), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1104), .B(new_n1105), .C1(G50), .C2(new_n879), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n818), .A2(G68), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n349), .A2(new_n887), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n413), .B(new_n1081), .C1(G150), .C2(new_n796), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n254), .B1(new_n796), .B2(G326), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n805), .A2(new_n823), .B1(new_n802), .B2(new_n820), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(G311), .A2(new_n887), .B1(new_n879), .B2(G317), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1113), .B1(new_n822), .B2(new_n788), .C1(new_n813), .C2(new_n253), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT48), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1112), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n1115), .B2(new_n1114), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT49), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1111), .B1(new_n283), .B2(new_n799), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1110), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n783), .B1(new_n1121), .B2(KEYINPUT113), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(KEYINPUT113), .B2(new_n1121), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n830), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n733), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n831), .A2(new_n1125), .B1(new_n542), .B2(new_n730), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n233), .A2(new_n261), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n441), .A2(G50), .ZN(new_n1128));
  XOR2_X1   g0928(.A(new_n1128), .B(KEYINPUT50), .Z(new_n1129));
  OAI211_X1 g0929(.A(new_n733), .B(new_n261), .C1(new_n397), .C2(new_n217), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n835), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1126), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1124), .B1(new_n1132), .B2(new_n842), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1123), .B(new_n1133), .C1(new_n711), .C2(new_n1096), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1103), .B(new_n1134), .C1(new_n777), .C2(new_n1100), .ZN(G393));
  OAI21_X1  g0935(.A(new_n778), .B1(new_n1062), .B2(new_n1068), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n835), .A2(new_n240), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n843), .B1(G97), .B2(new_n730), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1124), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n787), .A2(G150), .B1(new_n879), .B2(G159), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT51), .Z(new_n1141));
  OAI22_X1  g0941(.A1(new_n642), .A2(new_n799), .B1(new_n802), .B2(new_n219), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n254), .B1(new_n794), .B2(new_n889), .C1(new_n785), .C2(new_n789), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n1142), .B(new_n1143), .C1(G77), .C2(new_n806), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1141), .B(new_n1144), .C1(new_n441), .C2(new_n813), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT114), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n787), .A2(G317), .B1(new_n879), .B2(G311), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n1147), .B(KEYINPUT52), .Z(new_n1148));
  NOR2_X1   g0948(.A1(new_n802), .A2(new_n823), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n800), .B(new_n1149), .C1(G116), .C2(new_n806), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n413), .B1(new_n794), .B2(new_n822), .C1(new_n785), .C2(new_n253), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n818), .B2(G294), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1148), .A2(new_n1150), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1146), .A2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT115), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n1139), .B1(new_n1096), .B2(new_n1022), .C1(new_n1155), .C2(new_n783), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1136), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1046), .A2(new_n711), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n1060), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n721), .A2(KEYINPUT111), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1159), .A2(new_n1160), .A3(new_n1067), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1059), .A2(new_n1060), .A3(new_n1158), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1161), .A2(new_n1050), .A3(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1069), .A2(new_n731), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1157), .A2(new_n1164), .ZN(G390));
  NAND2_X1  g0965(.A1(new_n943), .A2(new_n989), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n725), .B1(new_n737), .B2(new_n741), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n980), .B1(new_n1167), .B2(new_n872), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1166), .B1(new_n1168), .B2(new_n977), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n718), .B(new_n872), .C1(new_n747), .C2(new_n772), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n977), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n989), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n856), .B1(new_n865), .B2(new_n853), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n857), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n980), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1173), .B1(new_n1176), .B2(new_n977), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n993), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1170), .B(new_n1172), .C1(new_n1177), .C2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n980), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n855), .B2(new_n857), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n989), .B1(new_n1181), .B2(new_n978), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1169), .B1(new_n1182), .B2(new_n993), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n718), .B1(new_n747), .B2(new_n947), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(new_n953), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1179), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1184), .A2(new_n853), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n978), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n741), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n692), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n1028), .B2(new_n693), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n707), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1180), .B1(new_n1192), .B2(new_n853), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1188), .A2(new_n1172), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n977), .B1(new_n773), .B2(new_n853), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n948), .A2(G330), .A3(new_n953), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(KEYINPUT116), .B1(new_n1197), .B2(new_n1181), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT116), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1199), .B(new_n1176), .C1(new_n1195), .C2(new_n1196), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1194), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1184), .A2(new_n512), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n995), .A2(new_n684), .A3(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1186), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1182), .A2(new_n993), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n1170), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(new_n1196), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1188), .A2(new_n1172), .A3(new_n1193), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1200), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1185), .B1(new_n1171), .B2(new_n977), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1199), .B1(new_n1210), .B2(new_n1176), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1208), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1203), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1207), .A2(new_n1212), .A3(new_n1179), .A4(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1204), .A2(new_n1214), .A3(new_n731), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1207), .A2(new_n778), .A3(new_n1179), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n788), .A2(new_n823), .B1(new_n542), .B2(new_n785), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n1083), .B2(G97), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT117), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n254), .B1(new_n826), .B2(G87), .ZN(new_n1220));
  XOR2_X1   g1020(.A(new_n1220), .B(KEYINPUT118), .Z(new_n1221));
  NOR2_X1   g1021(.A1(new_n794), .A2(new_n820), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n805), .A2(new_n217), .B1(new_n801), .B2(new_n283), .ZN(new_n1223));
  NOR4_X1   g1023(.A1(new_n1221), .A2(new_n892), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(KEYINPUT54), .B(G143), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1083), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n802), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(G150), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1229), .B(KEYINPUT53), .ZN(new_n1230));
  INV_X1    g1030(.A(G128), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n788), .A2(new_n1231), .B1(new_n799), .B2(new_n789), .ZN(new_n1232));
  INV_X1    g1032(.A(G125), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n254), .B1(new_n794), .B2(new_n1233), .C1(new_n785), .C2(new_n1085), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n805), .A2(new_n394), .B1(new_n801), .B2(new_n893), .ZN(new_n1235));
  NOR4_X1   g1035(.A1(new_n1230), .A2(new_n1232), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n1219), .A2(new_n1224), .B1(new_n1227), .B2(new_n1236), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n830), .B1(new_n349), .B2(new_n874), .C1(new_n1237), .C2(new_n783), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n993), .B2(new_n839), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1239), .B(KEYINPUT119), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1216), .A2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1215), .A2(new_n1241), .ZN(G378));
  OAI21_X1  g1042(.A(new_n988), .B1(new_n993), .B2(new_n989), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n986), .B2(new_n981), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n956), .A2(new_n959), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n718), .B1(new_n966), .B2(new_n967), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT122), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n353), .A2(new_n703), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT55), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1248), .B(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n683), .B2(new_n357), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n664), .B(new_n1250), .C1(new_n681), .C2(new_n682), .ZN(new_n1253));
  XOR2_X1   g1053(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1252), .A2(new_n1253), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n375), .A2(new_n1250), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n683), .A2(new_n357), .A3(new_n1251), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1254), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1247), .B1(new_n1256), .B2(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1255), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1257), .A2(new_n1254), .A3(new_n1258), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1261), .A2(new_n1262), .A3(KEYINPUT122), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1260), .A2(new_n1263), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1245), .A2(new_n1246), .A3(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1256), .A2(new_n1259), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1244), .B1(new_n1265), .B2(new_n1268), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n948), .A2(new_n953), .ZN(new_n1270));
  AOI21_X1  g1070(.A(KEYINPUT104), .B1(new_n1270), .B2(new_n958), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n954), .A2(new_n955), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1246), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1266), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1245), .A2(new_n1264), .A3(new_n1246), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1274), .A2(new_n994), .A3(new_n1275), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1269), .A2(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1213), .B1(new_n1186), .B2(new_n1201), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1277), .A2(KEYINPUT57), .A3(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n773), .A2(new_n853), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1280), .A2(new_n978), .ZN(new_n1281));
  AOI211_X1 g1081(.A(new_n1281), .B(new_n1169), .C1(new_n993), .C2(new_n1182), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1185), .B1(new_n1205), .B2(new_n1170), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1203), .B1(new_n1284), .B2(new_n1212), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1269), .A2(new_n1276), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n731), .B(new_n1279), .C1(new_n1287), .C2(KEYINPUT57), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1260), .A2(new_n839), .A3(new_n1263), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n779), .B1(G50), .B2(new_n874), .ZN(new_n1290));
  OAI22_X1  g1090(.A1(new_n788), .A2(new_n1233), .B1(new_n337), .B2(new_n805), .ZN(new_n1291));
  AOI22_X1  g1091(.A1(G132), .A2(new_n887), .B1(new_n1228), .B2(new_n1226), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1292), .B1(new_n810), .B2(new_n1085), .ZN(new_n1293));
  AOI211_X1 g1093(.A(new_n1291), .B(new_n1293), .C1(G128), .C2(new_n879), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  OR2_X1    g1095(.A1(new_n1295), .A2(KEYINPUT59), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(KEYINPUT59), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n880), .A2(G159), .ZN(new_n1298));
  AOI211_X1 g1098(.A(G33), .B(G41), .C1(new_n796), .C2(G124), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1296), .A2(new_n1297), .A3(new_n1298), .A4(new_n1299), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n254), .A2(G41), .ZN(new_n1301));
  OAI221_X1 g1101(.A(new_n1301), .B1(new_n823), .B2(new_n794), .C1(new_n289), .C2(new_n785), .ZN(new_n1302));
  AOI211_X1 g1102(.A(new_n1090), .B(new_n1302), .C1(G77), .C2(new_n1228), .ZN(new_n1303));
  OAI22_X1  g1103(.A1(new_n788), .A2(new_n283), .B1(new_n542), .B2(new_n801), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1304), .B1(G58), .B2(new_n880), .ZN(new_n1305));
  OAI211_X1 g1105(.A(new_n1303), .B(new_n1305), .C1(new_n439), .C2(new_n810), .ZN(new_n1306));
  XOR2_X1   g1106(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1301), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1309), .B(new_n789), .C1(G33), .C2(G41), .ZN(new_n1310));
  OR2_X1    g1110(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1300), .A2(new_n1308), .A3(new_n1310), .A4(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1290), .B1(new_n1312), .B2(new_n782), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1289), .A2(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1314), .B1(new_n1286), .B2(new_n777), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1288), .A2(new_n1316), .ZN(G375));
  NAND2_X1  g1117(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1042), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1203), .B(new_n1208), .C1(new_n1209), .C2(new_n1211), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1318), .A2(new_n1319), .A3(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n978), .A2(new_n839), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n830), .B1(G68), .B2(new_n874), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n805), .A2(new_n789), .ZN(new_n1324));
  OAI22_X1  g1124(.A1(new_n801), .A2(new_n1085), .B1(new_n799), .B2(new_n344), .ZN(new_n1325));
  AOI211_X1 g1125(.A(new_n1324), .B(new_n1325), .C1(G132), .C2(new_n787), .ZN(new_n1326));
  OAI221_X1 g1126(.A(new_n254), .B1(new_n794), .B2(new_n1231), .C1(new_n785), .C2(new_n1225), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1327), .B1(new_n818), .B2(G150), .ZN(new_n1328));
  OAI211_X1 g1128(.A(new_n1326), .B(new_n1328), .C1(new_n394), .C2(new_n827), .ZN(new_n1329));
  OAI22_X1  g1129(.A1(new_n788), .A2(new_n820), .B1(new_n823), .B2(new_n801), .ZN(new_n1330));
  OAI22_X1  g1130(.A1(new_n785), .A2(new_n283), .B1(new_n794), .B2(new_n253), .ZN(new_n1331));
  NOR3_X1   g1131(.A1(new_n1330), .A2(new_n1331), .A3(new_n1104), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n413), .B1(new_n799), .B2(new_n217), .ZN(new_n1333));
  XOR2_X1   g1133(.A(new_n1333), .B(KEYINPUT123), .Z(new_n1334));
  OAI211_X1 g1134(.A(new_n1332), .B(new_n1334), .C1(new_n289), .C2(new_n827), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n813), .A2(new_n542), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1329), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1323), .B1(new_n1337), .B2(new_n782), .ZN(new_n1338));
  AOI22_X1  g1138(.A1(new_n1212), .A2(new_n778), .B1(new_n1322), .B2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1321), .A2(new_n1339), .ZN(G381));
  INV_X1    g1140(.A(KEYINPUT124), .ZN(new_n1341));
  XNOR2_X1  g1141(.A(G375), .B(new_n1341), .ZN(new_n1342));
  OR3_X1    g1142(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1343));
  OR4_X1    g1143(.A1(G387), .A2(new_n1343), .A3(G381), .A4(G390), .ZN(new_n1344));
  OR3_X1    g1144(.A1(new_n1342), .A2(G378), .A3(new_n1344), .ZN(G407));
  NAND2_X1  g1145(.A1(new_n1216), .A2(new_n1240), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n732), .B1(new_n1318), .B2(new_n1186), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1346), .B1(new_n1347), .B2(new_n1214), .ZN(new_n1348));
  INV_X1    g1148(.A(G213), .ZN(new_n1349));
  NOR2_X1   g1149(.A1(new_n704), .A2(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1348), .A2(new_n1350), .ZN(new_n1351));
  OAI211_X1 g1151(.A(G407), .B(G213), .C1(new_n1342), .C2(new_n1351), .ZN(G409));
  NAND3_X1  g1152(.A1(new_n1269), .A2(new_n1276), .A3(KEYINPUT57), .ZN(new_n1353));
  OAI21_X1  g1153(.A(new_n731), .B1(new_n1285), .B2(new_n1353), .ZN(new_n1354));
  AOI21_X1  g1154(.A(KEYINPUT57), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1355));
  OAI211_X1 g1155(.A(G378), .B(new_n1316), .C1(new_n1354), .C2(new_n1355), .ZN(new_n1356));
  NOR3_X1   g1156(.A1(new_n1285), .A2(new_n1042), .A3(new_n1286), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1348), .B1(new_n1357), .B2(new_n1315), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1356), .A2(new_n1358), .ZN(new_n1359));
  INV_X1    g1159(.A(new_n1350), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1359), .A2(new_n1360), .ZN(new_n1361));
  AOI21_X1  g1161(.A(new_n732), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1201), .A2(KEYINPUT60), .A3(new_n1203), .ZN(new_n1363));
  INV_X1    g1163(.A(KEYINPUT60), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1320), .A2(new_n1364), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1362), .A2(new_n1363), .A3(new_n1365), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1366), .A2(new_n1339), .ZN(new_n1367));
  INV_X1    g1167(.A(KEYINPUT125), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1367), .A2(new_n1368), .ZN(new_n1369));
  NAND3_X1  g1169(.A1(new_n1366), .A2(KEYINPUT125), .A3(new_n1339), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1369), .A2(new_n899), .A3(new_n1370), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1350), .A2(G2897), .ZN(new_n1372));
  NAND3_X1  g1172(.A1(new_n1367), .A2(new_n1368), .A3(G384), .ZN(new_n1373));
  AND3_X1   g1173(.A1(new_n1371), .A2(new_n1372), .A3(new_n1373), .ZN(new_n1374));
  AOI21_X1  g1174(.A(new_n1372), .B1(new_n1371), .B2(new_n1373), .ZN(new_n1375));
  OAI21_X1  g1175(.A(new_n1361), .B1(new_n1374), .B2(new_n1375), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1371), .A2(new_n1373), .ZN(new_n1377));
  NAND3_X1  g1177(.A1(new_n1377), .A2(new_n1359), .A3(new_n1360), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1378), .A2(KEYINPUT62), .ZN(new_n1379));
  INV_X1    g1179(.A(KEYINPUT61), .ZN(new_n1380));
  INV_X1    g1180(.A(KEYINPUT62), .ZN(new_n1381));
  NAND4_X1  g1181(.A1(new_n1377), .A2(new_n1359), .A3(new_n1381), .A4(new_n1360), .ZN(new_n1382));
  NAND4_X1  g1182(.A1(new_n1376), .A2(new_n1379), .A3(new_n1380), .A4(new_n1382), .ZN(new_n1383));
  XNOR2_X1  g1183(.A(G393), .B(G396), .ZN(new_n1384));
  AND2_X1   g1184(.A1(new_n1157), .A2(new_n1164), .ZN(new_n1385));
  AOI21_X1  g1185(.A(new_n1050), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1386));
  OAI21_X1  g1186(.A(new_n1319), .B1(new_n1386), .B2(new_n1101), .ZN(new_n1387));
  AOI21_X1  g1187(.A(new_n1040), .B1(new_n1387), .B2(new_n777), .ZN(new_n1388));
  INV_X1    g1188(.A(new_n1098), .ZN(new_n1389));
  NOR3_X1   g1189(.A1(new_n1385), .A2(new_n1388), .A3(new_n1389), .ZN(new_n1390));
  AOI21_X1  g1190(.A(G390), .B1(new_n1071), .B2(new_n1098), .ZN(new_n1391));
  OAI21_X1  g1191(.A(new_n1384), .B1(new_n1390), .B2(new_n1391), .ZN(new_n1392));
  INV_X1    g1192(.A(new_n1384), .ZN(new_n1393));
  OAI21_X1  g1193(.A(new_n1385), .B1(new_n1388), .B2(new_n1389), .ZN(new_n1394));
  NAND3_X1  g1194(.A1(new_n1071), .A2(new_n1098), .A3(G390), .ZN(new_n1395));
  NAND3_X1  g1195(.A1(new_n1393), .A2(new_n1394), .A3(new_n1395), .ZN(new_n1396));
  NAND2_X1  g1196(.A1(new_n1392), .A2(new_n1396), .ZN(new_n1397));
  NAND2_X1  g1197(.A1(new_n1383), .A2(new_n1397), .ZN(new_n1398));
  INV_X1    g1198(.A(KEYINPUT126), .ZN(new_n1399));
  NAND2_X1  g1199(.A1(new_n1378), .A2(new_n1399), .ZN(new_n1400));
  NAND2_X1  g1200(.A1(new_n1400), .A2(KEYINPUT63), .ZN(new_n1401));
  INV_X1    g1201(.A(KEYINPUT63), .ZN(new_n1402));
  NAND3_X1  g1202(.A1(new_n1378), .A2(new_n1399), .A3(new_n1402), .ZN(new_n1403));
  NAND3_X1  g1203(.A1(new_n1392), .A2(new_n1380), .A3(new_n1396), .ZN(new_n1404));
  NAND2_X1  g1204(.A1(new_n1404), .A2(KEYINPUT127), .ZN(new_n1405));
  INV_X1    g1205(.A(KEYINPUT127), .ZN(new_n1406));
  NAND4_X1  g1206(.A1(new_n1392), .A2(new_n1406), .A3(new_n1396), .A4(new_n1380), .ZN(new_n1407));
  NAND2_X1  g1207(.A1(new_n1405), .A2(new_n1407), .ZN(new_n1408));
  NAND4_X1  g1208(.A1(new_n1401), .A2(new_n1376), .A3(new_n1403), .A4(new_n1408), .ZN(new_n1409));
  NAND2_X1  g1209(.A1(new_n1398), .A2(new_n1409), .ZN(G405));
  NAND2_X1  g1210(.A1(new_n1370), .A2(new_n899), .ZN(new_n1411));
  AOI21_X1  g1211(.A(KEYINPUT125), .B1(new_n1366), .B2(new_n1339), .ZN(new_n1412));
  NOR2_X1   g1212(.A1(new_n1411), .A2(new_n1412), .ZN(new_n1413));
  INV_X1    g1213(.A(new_n1373), .ZN(new_n1414));
  NOR2_X1   g1214(.A1(new_n1413), .A2(new_n1414), .ZN(new_n1415));
  INV_X1    g1215(.A(new_n1356), .ZN(new_n1416));
  AOI21_X1  g1216(.A(G378), .B1(new_n1288), .B2(new_n1316), .ZN(new_n1417));
  OR3_X1    g1217(.A1(new_n1415), .A2(new_n1416), .A3(new_n1417), .ZN(new_n1418));
  INV_X1    g1218(.A(new_n1397), .ZN(new_n1419));
  OAI21_X1  g1219(.A(new_n1415), .B1(new_n1416), .B2(new_n1417), .ZN(new_n1420));
  AND3_X1   g1220(.A1(new_n1418), .A2(new_n1419), .A3(new_n1420), .ZN(new_n1421));
  AOI21_X1  g1221(.A(new_n1419), .B1(new_n1418), .B2(new_n1420), .ZN(new_n1422));
  NOR2_X1   g1222(.A1(new_n1421), .A2(new_n1422), .ZN(G402));
endmodule


