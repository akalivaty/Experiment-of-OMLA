//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 1 0 0 0 1 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 0 0 0 0 0 0 0 1 1 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n564,
    new_n566, new_n567, new_n568, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n629, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1215, new_n1216, new_n1217;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT64), .Z(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  OR2_X1    g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  OAI21_X1  g042(.A(G2105), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  OAI211_X1 g047(.A(G137), .B(new_n470), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G101), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n476));
  INV_X1    g051(.A(G2104), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(G2105), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n470), .A2(KEYINPUT65), .A3(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n475), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR3_X1   g055(.A1(new_n469), .A2(new_n474), .A3(new_n480), .ZN(G160));
  XNOR2_X1  g056(.A(KEYINPUT3), .B(G2104), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(new_n470), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT66), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n485), .B(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G112), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n477), .B1(new_n490), .B2(G2105), .ZN(new_n491));
  AOI22_X1  g066(.A1(new_n488), .A2(G136), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n487), .A2(new_n492), .ZN(G162));
  OAI211_X1 g068(.A(G138), .B(new_n470), .C1(new_n471), .C2(new_n472), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n482), .A2(KEYINPUT4), .A3(G138), .A4(new_n470), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  XNOR2_X1  g075(.A(KEYINPUT67), .B(G114), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(new_n470), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n482), .A2(G126), .A3(G2105), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n498), .A2(new_n504), .ZN(G164));
  NAND2_X1  g080(.A1(KEYINPUT68), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT68), .A3(G543), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n507), .A2(new_n509), .A3(G62), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT69), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT69), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n507), .A2(new_n509), .A3(new_n512), .A4(G62), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n511), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G651), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT6), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G651), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n507), .A2(new_n509), .A3(new_n518), .A4(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n518), .A2(new_n520), .A3(G543), .ZN(new_n523));
  INV_X1    g098(.A(G50), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n521), .A2(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n516), .A2(new_n526), .A3(KEYINPUT70), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n528));
  INV_X1    g103(.A(new_n514), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n529), .B1(new_n510), .B2(KEYINPUT69), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n517), .B1(new_n530), .B2(new_n513), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n528), .B1(new_n531), .B2(new_n525), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n527), .A2(new_n532), .ZN(G166));
  INV_X1    g108(.A(new_n521), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G89), .ZN(new_n535));
  INV_X1    g110(.A(new_n523), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G51), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n507), .A2(new_n509), .A3(G63), .A4(G651), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  NAND4_X1  g115(.A1(new_n535), .A2(new_n537), .A3(new_n538), .A4(new_n540), .ZN(G286));
  INV_X1    g116(.A(G286), .ZN(G168));
  NAND3_X1  g117(.A1(new_n507), .A2(new_n509), .A3(G64), .ZN(new_n543));
  NAND2_X1  g118(.A1(G77), .A2(G543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n517), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n534), .A2(G90), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT71), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n536), .A2(G52), .ZN(new_n549));
  NAND4_X1  g124(.A1(new_n546), .A2(new_n547), .A3(new_n548), .A4(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(G90), .ZN(new_n551));
  INV_X1    g126(.A(G52), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n521), .A2(new_n551), .B1(new_n523), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g128(.A(KEYINPUT71), .B1(new_n553), .B2(new_n545), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n550), .A2(new_n554), .ZN(G171));
  INV_X1    g130(.A(G81), .ZN(new_n556));
  INV_X1    g131(.A(G43), .ZN(new_n557));
  OAI22_X1  g132(.A1(new_n521), .A2(new_n556), .B1(new_n523), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n507), .A2(new_n509), .A3(G56), .ZN(new_n559));
  NAND2_X1  g134(.A1(G68), .A2(G543), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n517), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n564));
  XOR2_X1   g139(.A(new_n564), .B(KEYINPUT72), .Z(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT73), .ZN(G188));
  NAND4_X1  g144(.A1(new_n518), .A2(new_n520), .A3(G53), .A4(G543), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT9), .ZN(new_n571));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n507), .A2(new_n509), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G651), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n534), .A2(G91), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n571), .A2(new_n576), .A3(new_n577), .ZN(G299));
  INV_X1    g153(.A(G171), .ZN(G301));
  INV_X1    g154(.A(KEYINPUT74), .ZN(new_n580));
  AOI21_X1  g155(.A(KEYINPUT70), .B1(new_n516), .B2(new_n526), .ZN(new_n581));
  NOR3_X1   g156(.A1(new_n531), .A2(new_n528), .A3(new_n525), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n527), .A2(new_n532), .A3(KEYINPUT74), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n583), .A2(new_n584), .ZN(G303));
  INV_X1    g160(.A(G87), .ZN(new_n586));
  INV_X1    g161(.A(G49), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n521), .A2(new_n586), .B1(new_n523), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(G74), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n517), .B1(new_n573), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G288));
  NAND3_X1  g167(.A1(new_n507), .A2(new_n509), .A3(G61), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n593), .A2(KEYINPUT75), .B1(G73), .B2(G543), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT75), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n507), .A2(new_n509), .A3(new_n595), .A4(G61), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n517), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(G86), .ZN(new_n598));
  INV_X1    g173(.A(G48), .ZN(new_n599));
  OAI22_X1  g174(.A1(new_n521), .A2(new_n598), .B1(new_n523), .B2(new_n599), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n597), .A2(new_n600), .ZN(G305));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  XOR2_X1   g177(.A(KEYINPUT76), .B(G47), .Z(new_n603));
  OAI22_X1  g178(.A1(new_n521), .A2(new_n602), .B1(new_n603), .B2(new_n523), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n507), .A2(new_n509), .A3(G60), .ZN(new_n605));
  NAND2_X1  g180(.A1(G72), .A2(G543), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n517), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(G290));
  NAND3_X1  g184(.A1(new_n507), .A2(new_n509), .A3(G66), .ZN(new_n610));
  NAND2_X1  g185(.A1(G79), .A2(G543), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G651), .ZN(new_n613));
  INV_X1    g188(.A(G54), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n523), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n613), .A2(KEYINPUT77), .A3(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT77), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n517), .B1(new_n610), .B2(new_n611), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n615), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(G92), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n521), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT10), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  MUX2_X1   g200(.A(new_n625), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g201(.A(new_n625), .B(G301), .S(G868), .Z(G321));
  NAND2_X1  g202(.A1(G286), .A2(G868), .ZN(new_n628));
  INV_X1    g203(.A(G299), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(G868), .ZN(G297));
  OAI21_X1  g205(.A(new_n628), .B1(new_n629), .B2(G868), .ZN(G280));
  AND2_X1   g206(.A1(new_n621), .A2(new_n624), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT78), .B(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(G860), .B2(new_n633), .ZN(G148));
  INV_X1    g209(.A(KEYINPUT80), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n632), .A2(new_n633), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT79), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(G868), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n635), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n637), .A2(KEYINPUT80), .A3(G868), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n640), .B(new_n641), .C1(G868), .C2(new_n562), .ZN(G323));
  XNOR2_X1  g217(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g218(.A1(new_n478), .A2(new_n479), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(new_n482), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT13), .Z(new_n648));
  INV_X1    g223(.A(G2100), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n484), .A2(G123), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n488), .A2(G135), .ZN(new_n653));
  NOR2_X1   g228(.A1(G99), .A2(G2105), .ZN(new_n654));
  OAI21_X1  g229(.A(G2104), .B1(new_n470), .B2(G111), .ZN(new_n655));
  OAI211_X1 g230(.A(new_n652), .B(new_n653), .C1(new_n654), .C2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(G2096), .Z(new_n657));
  NAND3_X1  g232(.A1(new_n650), .A2(new_n651), .A3(new_n657), .ZN(G156));
  XNOR2_X1  g233(.A(KEYINPUT15), .B(G2435), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2438), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2427), .B(G2430), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT82), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(KEYINPUT14), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT83), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n665), .B1(new_n660), .B2(new_n662), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2443), .B(G2446), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n666), .B(new_n667), .Z(new_n668));
  XNOR2_X1  g243(.A(G2451), .B(G2454), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT16), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n666), .B(new_n667), .ZN(new_n672));
  INV_X1    g247(.A(new_n670), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1341), .B(G1348), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n671), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT84), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n675), .B1(new_n671), .B2(new_n674), .ZN(new_n679));
  INV_X1    g254(.A(G14), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n678), .A2(new_n681), .ZN(G401));
  XOR2_X1   g257(.A(G2072), .B(G2078), .Z(new_n683));
  XOR2_X1   g258(.A(G2084), .B(G2090), .Z(new_n684));
  XNOR2_X1  g259(.A(G2067), .B(G2678), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT85), .B(KEYINPUT18), .Z(new_n687));
  AOI21_X1  g262(.A(new_n683), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n686), .A2(KEYINPUT17), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n684), .A2(new_n685), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n687), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  MUX2_X1   g266(.A(new_n688), .B(new_n683), .S(new_n691), .Z(new_n692));
  XNOR2_X1  g267(.A(G2096), .B(G2100), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(G227));
  XOR2_X1   g269(.A(G1971), .B(G1976), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT86), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT19), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1956), .B(G2474), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1961), .B(G1966), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT20), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n698), .A2(new_n699), .ZN(new_n703));
  NOR3_X1   g278(.A1(new_n697), .A2(new_n700), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(new_n697), .B2(new_n703), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1991), .B(G1996), .ZN(new_n706));
  INV_X1    g281(.A(G1986), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n702), .A2(new_n705), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n708), .B1(new_n702), .B2(new_n705), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT87), .B(G1981), .ZN(new_n712));
  NOR3_X1   g287(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT88), .Z(new_n716));
  OAI21_X1  g291(.A(new_n712), .B1(new_n710), .B2(new_n711), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n714), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n716), .ZN(new_n719));
  INV_X1    g294(.A(new_n712), .ZN(new_n720));
  INV_X1    g295(.A(new_n711), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(new_n709), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n719), .B1(new_n722), .B2(new_n713), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n718), .A2(new_n723), .ZN(G229));
  INV_X1    g299(.A(KEYINPUT90), .ZN(new_n725));
  OR3_X1    g300(.A1(new_n725), .A2(G16), .A3(G23), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(G16), .B2(G23), .ZN(new_n727));
  INV_X1    g302(.A(G16), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n726), .B(new_n727), .C1(G288), .C2(new_n728), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT33), .B(G1976), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n728), .A2(G6), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G305), .B2(G16), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT32), .B(G1981), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT89), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n731), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n728), .A2(G22), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G166), .B2(new_n728), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G1971), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(G1971), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n734), .A2(new_n736), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n738), .A2(new_n741), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n744), .A2(KEYINPUT34), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(KEYINPUT34), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n484), .A2(G119), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n488), .A2(G131), .ZN(new_n748));
  NOR2_X1   g323(.A1(G95), .A2(G2105), .ZN(new_n749));
  OAI21_X1  g324(.A(G2104), .B1(new_n470), .B2(G107), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n747), .B(new_n748), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  MUX2_X1   g326(.A(G25), .B(new_n751), .S(G29), .Z(new_n752));
  XOR2_X1   g327(.A(KEYINPUT35), .B(G1991), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G16), .A2(G24), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n608), .B2(G16), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n754), .B1(G1986), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G1986), .B2(new_n756), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n745), .A2(new_n746), .A3(new_n758), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT36), .Z(new_n760));
  INV_X1    g335(.A(G28), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n761), .A2(KEYINPUT30), .ZN(new_n762));
  AOI21_X1  g337(.A(G29), .B1(new_n761), .B2(KEYINPUT30), .ZN(new_n763));
  OR2_X1    g338(.A1(KEYINPUT31), .A2(G11), .ZN(new_n764));
  NAND2_X1  g339(.A1(KEYINPUT31), .A2(G11), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n762), .A2(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(G29), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n766), .B1(new_n656), .B2(new_n767), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT95), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n728), .A2(G19), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n562), .B2(new_n728), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(G1341), .Z(new_n772));
  NOR2_X1   g347(.A1(G168), .A2(new_n728), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n728), .B2(G21), .ZN(new_n774));
  INV_X1    g349(.A(G1966), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n769), .A2(new_n772), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n767), .A2(G26), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT28), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n484), .A2(G128), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n488), .A2(G140), .ZN(new_n781));
  OR2_X1    g356(.A1(G104), .A2(G2105), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n782), .B(G2104), .C1(G116), .C2(new_n470), .ZN(new_n783));
  AND3_X1   g358(.A1(new_n780), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n779), .B1(new_n784), .B2(new_n767), .ZN(new_n785));
  INV_X1    g360(.A(G2067), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n767), .A2(G27), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G164), .B2(new_n767), .ZN(new_n789));
  INV_X1    g364(.A(G2078), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n787), .B(new_n791), .C1(new_n775), .C2(new_n774), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n728), .A2(G20), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT23), .Z(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G299), .B2(G16), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(G1956), .Z(new_n796));
  NOR3_X1   g371(.A1(new_n777), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n767), .A2(G32), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT94), .B(KEYINPUT26), .ZN(new_n799));
  NAND3_X1  g374(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G105), .B2(new_n644), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n484), .A2(G129), .B1(G141), .B2(new_n488), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n798), .B1(new_n805), .B2(new_n767), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT27), .B(G1996), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n767), .A2(G33), .ZN(new_n809));
  NAND2_X1  g384(.A1(G115), .A2(G2104), .ZN(new_n810));
  INV_X1    g385(.A(G127), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n483), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n470), .B1(new_n812), .B2(KEYINPUT93), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(KEYINPUT93), .B2(new_n812), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT91), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT25), .ZN(new_n817));
  AOI21_X1  g392(.A(KEYINPUT92), .B1(new_n488), .B2(G139), .ZN(new_n818));
  AND3_X1   g393(.A1(new_n488), .A2(KEYINPUT92), .A3(G139), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n814), .B(new_n817), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n809), .B1(new_n820), .B2(G29), .ZN(new_n821));
  INV_X1    g396(.A(G2072), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n821), .A2(new_n822), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT24), .ZN(new_n825));
  INV_X1    g400(.A(G34), .ZN(new_n826));
  AOI21_X1  g401(.A(G29), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n825), .B2(new_n826), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G160), .B2(new_n767), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(G2084), .ZN(new_n830));
  NOR4_X1   g405(.A1(new_n808), .A2(new_n823), .A3(new_n824), .A4(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(G5), .A2(G16), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT96), .Z(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(G301), .B2(new_n728), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(G1961), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n797), .A2(new_n831), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n767), .A2(G35), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(G162), .B2(new_n767), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT97), .Z(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT29), .ZN(new_n840));
  INV_X1    g415(.A(G2090), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n728), .A2(G4), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n632), .B2(new_n728), .ZN(new_n844));
  INV_X1    g419(.A(G1348), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n840), .A2(new_n841), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n842), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NOR3_X1   g423(.A1(new_n760), .A2(new_n836), .A3(new_n848), .ZN(G311));
  INV_X1    g424(.A(G311), .ZN(G150));
  NAND2_X1  g425(.A1(G80), .A2(G543), .ZN(new_n851));
  INV_X1    g426(.A(G67), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n851), .B1(new_n573), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(KEYINPUT98), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT98), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n855), .B(new_n851), .C1(new_n573), .C2(new_n852), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n854), .A2(G651), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(KEYINPUT99), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n854), .A2(new_n859), .A3(G651), .A4(new_n856), .ZN(new_n860));
  INV_X1    g435(.A(G93), .ZN(new_n861));
  INV_X1    g436(.A(G55), .ZN(new_n862));
  OAI22_X1  g437(.A1(new_n521), .A2(new_n861), .B1(new_n523), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(KEYINPUT100), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT100), .ZN(new_n865));
  OAI221_X1 g440(.A(new_n865), .B1(new_n523), .B2(new_n862), .C1(new_n521), .C2(new_n861), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n858), .A2(new_n860), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n562), .A2(KEYINPUT101), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n871));
  NOR3_X1   g446(.A1(new_n558), .A2(new_n561), .A3(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n868), .A2(new_n870), .A3(new_n873), .ZN(new_n874));
  AOI22_X1  g449(.A1(new_n857), .A2(KEYINPUT99), .B1(new_n866), .B2(new_n864), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n875), .A2(KEYINPUT101), .A3(new_n562), .A4(new_n860), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT38), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n632), .A2(G559), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n878), .B(new_n879), .Z(new_n880));
  AND2_X1   g455(.A1(new_n880), .A2(KEYINPUT39), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(KEYINPUT39), .ZN(new_n882));
  NOR3_X1   g457(.A1(new_n881), .A2(new_n882), .A3(G860), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n868), .A2(G860), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT37), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n883), .A2(new_n885), .ZN(G145));
  INV_X1    g461(.A(KEYINPUT103), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n820), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n889));
  AOI21_X1  g464(.A(KEYINPUT4), .B1(new_n488), .B2(G138), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n494), .A2(new_n495), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n504), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT102), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n780), .A2(new_n781), .A3(new_n783), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n888), .B(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n647), .ZN(new_n899));
  OR2_X1    g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n484), .A2(G130), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n488), .A2(G142), .ZN(new_n902));
  NOR2_X1   g477(.A1(G106), .A2(G2105), .ZN(new_n903));
  OAI21_X1  g478(.A(G2104), .B1(new_n470), .B2(G118), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n901), .B(new_n902), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  XOR2_X1   g480(.A(new_n751), .B(new_n905), .Z(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(new_n805), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n898), .A2(new_n899), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n900), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n907), .B1(new_n900), .B2(new_n908), .ZN(new_n910));
  XNOR2_X1  g485(.A(G162), .B(G160), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(new_n656), .ZN(new_n912));
  OR3_X1    g487(.A1(new_n909), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(G37), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n912), .B1(new_n909), .B2(new_n910), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g492(.A1(new_n868), .A2(new_n639), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n625), .A2(new_n629), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n621), .A2(new_n624), .A3(G299), .ZN(new_n920));
  XOR2_X1   g495(.A(KEYINPUT104), .B(KEYINPUT41), .Z(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n920), .ZN(new_n924));
  AOI21_X1  g499(.A(G299), .B1(new_n621), .B2(new_n624), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n923), .B1(new_n926), .B2(KEYINPUT41), .ZN(new_n927));
  INV_X1    g502(.A(new_n926), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n637), .B(new_n877), .ZN(new_n929));
  MUX2_X1   g504(.A(new_n927), .B(new_n928), .S(new_n929), .Z(new_n930));
  NOR2_X1   g505(.A1(new_n597), .A2(new_n600), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(G290), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n608), .B1(new_n597), .B2(new_n600), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n527), .A2(new_n532), .A3(G288), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(G288), .B1(new_n527), .B2(new_n532), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(G166), .A2(new_n591), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n939), .A2(new_n935), .A3(new_n932), .A4(new_n933), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT42), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n938), .A2(new_n940), .A3(KEYINPUT105), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT105), .B1(new_n938), .B2(new_n940), .ZN(new_n943));
  OR2_X1    g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n941), .B1(new_n944), .B2(KEYINPUT42), .ZN(new_n945));
  XOR2_X1   g520(.A(new_n930), .B(new_n945), .Z(new_n946));
  OAI21_X1  g521(.A(new_n918), .B1(new_n946), .B2(new_n639), .ZN(G295));
  OAI21_X1  g522(.A(new_n918), .B1(new_n946), .B2(new_n639), .ZN(G331));
  NOR2_X1   g523(.A1(new_n942), .A2(new_n943), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n550), .A2(new_n554), .A3(G286), .ZN(new_n950));
  AOI21_X1  g525(.A(G286), .B1(new_n550), .B2(new_n554), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n874), .A2(new_n952), .A3(new_n876), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n952), .B1(new_n874), .B2(new_n876), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n927), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n952), .ZN(new_n956));
  AOI211_X1 g531(.A(new_n872), .B(new_n869), .C1(new_n875), .C2(new_n860), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n873), .B1(new_n868), .B2(new_n870), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n874), .A2(new_n952), .A3(new_n876), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(new_n928), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n955), .A2(new_n961), .A3(KEYINPUT106), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT106), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n959), .A2(new_n963), .A3(new_n928), .A4(new_n960), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n949), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n914), .B1(new_n965), .B2(KEYINPUT107), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT107), .ZN(new_n967));
  AOI211_X1 g542(.A(new_n967), .B(new_n949), .C1(new_n962), .C2(new_n964), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n962), .A2(new_n949), .A3(new_n964), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT43), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(KEYINPUT108), .B1(new_n926), .B2(new_n922), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT41), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n972), .B1(new_n973), .B2(new_n928), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n926), .A2(KEYINPUT108), .A3(new_n922), .ZN(new_n975));
  OAI22_X1  g550(.A1(new_n974), .A2(new_n975), .B1(new_n953), .B2(new_n954), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n944), .B1(new_n976), .B2(new_n961), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT43), .ZN(new_n978));
  NOR4_X1   g553(.A1(new_n966), .A2(new_n968), .A3(new_n977), .A4(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT44), .B1(new_n971), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n978), .B1(new_n969), .B2(new_n970), .ZN(new_n982));
  NOR4_X1   g557(.A1(new_n966), .A2(new_n968), .A3(new_n977), .A4(KEYINPUT43), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n980), .A2(new_n984), .ZN(G397));
  INV_X1    g560(.A(G1384), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT45), .B1(new_n895), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n480), .ZN(new_n988));
  XOR2_X1   g563(.A(KEYINPUT109), .B(G40), .Z(new_n989));
  NAND4_X1  g564(.A1(new_n468), .A2(new_n988), .A3(new_n473), .A4(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  OR3_X1    g567(.A1(new_n992), .A2(KEYINPUT112), .A3(G1996), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT112), .B1(new_n992), .B2(G1996), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n804), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n784), .A2(new_n786), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n896), .A2(G2067), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n998), .B(KEYINPUT113), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n804), .A2(G1996), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n992), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n995), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n992), .ZN(new_n1003));
  INV_X1    g578(.A(new_n753), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n751), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n751), .A2(new_n1004), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1003), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  AND2_X1   g582(.A1(new_n1002), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(G290), .A2(G1986), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1009), .A2(KEYINPUT110), .ZN(new_n1010));
  NAND2_X1  g585(.A1(G290), .A2(G1986), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1012), .A2(new_n992), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n1013), .B(KEYINPUT111), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1008), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n1016));
  INV_X1    g591(.A(G8), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g593(.A(KEYINPUT45), .B(new_n986), .C1(new_n498), .C2(new_n504), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(new_n991), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n775), .B1(new_n987), .B2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g596(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n895), .A2(new_n986), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G2084), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n986), .B1(new_n498), .B2(new_n504), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n990), .B1(new_n1025), .B2(KEYINPUT50), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1023), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n1021), .A2(G286), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(G286), .B1(new_n1021), .B2(new_n1027), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1018), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1021), .A2(G168), .A3(new_n1027), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n1031), .A2(G8), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1030), .B(KEYINPUT62), .C1(KEYINPUT51), .C2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT62), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1018), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT102), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT102), .B1(new_n496), .B2(new_n497), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n1037), .A2(new_n1038), .A3(new_n504), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1036), .B1(new_n1039), .B2(G1384), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1019), .A2(new_n991), .ZN(new_n1041));
  AOI21_X1  g616(.A(G1966), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n1023), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1043));
  OAI21_X1  g618(.A(G168), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1021), .A2(G286), .A3(new_n1027), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1035), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT51), .B1(new_n1031), .B2(G8), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1034), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1038), .A2(new_n504), .ZN(new_n1049));
  AOI21_X1  g624(.A(G1384), .B1(new_n1049), .B2(new_n894), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1041), .B(new_n790), .C1(new_n1050), .C2(KEYINPUT45), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT120), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT120), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1040), .A2(new_n1053), .A3(new_n790), .A4(new_n1041), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1052), .A2(KEYINPUT53), .A3(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n895), .A2(KEYINPUT45), .A3(new_n986), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n990), .B1(new_n1025), .B2(new_n1036), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1056), .A2(new_n790), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT53), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1060));
  INV_X1    g635(.A(G1961), .ZN(new_n1061));
  AOI22_X1  g636(.A1(new_n1058), .A2(new_n1059), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(G301), .B1(new_n1055), .B2(new_n1062), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1033), .A2(new_n1048), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT121), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(new_n465), .B2(new_n467), .ZN(new_n1068));
  OAI21_X1  g643(.A(G125), .B1(new_n471), .B2(new_n472), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1069), .A2(KEYINPUT121), .A3(new_n466), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1068), .A2(G2105), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G40), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n474), .A2(new_n480), .A3(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1071), .A2(KEYINPUT122), .A3(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT53), .B1(new_n790), .B2(KEYINPUT123), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1075), .B1(KEYINPUT123), .B2(new_n790), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT122), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1079), .A2(new_n1040), .A3(new_n1056), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1065), .A2(new_n1066), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(G171), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT125), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1055), .A2(G301), .A3(new_n1062), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT125), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1081), .A2(new_n1085), .A3(G171), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1083), .A2(KEYINPUT54), .A3(new_n1084), .A4(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1081), .A2(G171), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1088), .B1(new_n1063), .B2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1087), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT56), .B(G2072), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1056), .A2(new_n1057), .A3(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n991), .B1(new_n1025), .B2(KEYINPUT50), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n895), .A2(new_n986), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1022), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1095), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1094), .B1(new_n1098), .B2(G1956), .ZN(new_n1099));
  XOR2_X1   g674(.A(G299), .B(KEYINPUT57), .Z(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(G1348), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1103));
  AND4_X1   g678(.A1(new_n986), .A2(new_n895), .A3(new_n786), .A4(new_n991), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1102), .B1(new_n625), .B2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1100), .B(new_n1094), .C1(new_n1098), .C2(G1956), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1105), .A2(KEYINPUT60), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT60), .ZN(new_n1110));
  NOR3_X1   g685(.A1(new_n1103), .A2(new_n1110), .A3(new_n1104), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n632), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1060), .A2(new_n845), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1104), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1114), .A2(KEYINPUT60), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1116), .A2(KEYINPUT119), .A3(new_n625), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1109), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(KEYINPUT118), .A2(KEYINPUT61), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1102), .A2(new_n1107), .A3(new_n1122), .ZN(new_n1123));
  OR2_X1    g698(.A1(new_n1107), .A2(new_n1122), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1096), .A2(new_n990), .ZN(new_n1127));
  XNOR2_X1  g702(.A(KEYINPUT58), .B(G1341), .ZN(new_n1128));
  OAI22_X1  g703(.A1(G1996), .A2(new_n1126), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1125), .B1(new_n1129), .B2(new_n562), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1129), .A2(new_n1125), .A3(new_n562), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1123), .B(new_n1124), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1108), .B1(new_n1120), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1064), .B1(new_n1092), .B2(new_n1133), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n583), .A2(KEYINPUT55), .A3(G8), .A4(new_n584), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT115), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT116), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(G303), .A2(KEYINPUT115), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT116), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(G303), .A2(G8), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT55), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1139), .A2(new_n1143), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1126), .ZN(new_n1148));
  OAI22_X1  g723(.A1(new_n1148), .A2(G1971), .B1(G2090), .B2(new_n1060), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1149), .A2(G8), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n1098), .A2(new_n841), .ZN(new_n1152));
  AOI21_X1  g727(.A(G1971), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1153));
  OAI21_X1  g728(.A(G8), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1139), .A2(new_n1143), .A3(new_n1154), .A4(new_n1146), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1127), .A2(new_n1017), .ZN(new_n1156));
  INV_X1    g731(.A(G1976), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1156), .B1(new_n1157), .B2(G288), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(KEYINPUT52), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT52), .B1(G288), .B2(new_n1157), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1156), .B(new_n1160), .C1(new_n1157), .C2(G288), .ZN(new_n1161));
  NAND2_X1  g736(.A1(G305), .A2(G1981), .ZN(new_n1162));
  INV_X1    g737(.A(G1981), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n931), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT49), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1162), .A2(KEYINPUT49), .A3(new_n1164), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1167), .A2(new_n1156), .A3(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1159), .A2(new_n1161), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1170), .ZN(new_n1171));
  AND4_X1   g746(.A1(KEYINPUT124), .A2(new_n1151), .A3(new_n1155), .A4(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1170), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1173));
  AOI21_X1  g748(.A(KEYINPUT124), .B1(new_n1173), .B2(new_n1155), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1134), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1173), .ZN(new_n1176));
  OAI211_X1 g751(.A(G8), .B(new_n1029), .C1(new_n1147), .C2(new_n1149), .ZN(new_n1177));
  OAI21_X1  g752(.A(KEYINPUT63), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g753(.A1(G288), .A2(G1976), .ZN(new_n1179));
  AOI22_X1  g754(.A1(new_n1169), .A2(new_n1179), .B1(new_n1163), .B2(new_n931), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT117), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1156), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1182), .B1(new_n1181), .B2(new_n1180), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1151), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1183), .B1(new_n1184), .B2(new_n1171), .ZN(new_n1185));
  NOR3_X1   g760(.A1(new_n1044), .A2(KEYINPUT63), .A3(new_n1017), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1173), .A2(new_n1155), .A3(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1178), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1015), .B1(new_n1175), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT46), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n993), .A2(new_n1190), .A3(new_n994), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n1191), .B(new_n1192), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1190), .B1(new_n993), .B2(new_n994), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n992), .B1(new_n999), .B2(new_n805), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1193), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT47), .ZN(new_n1198));
  XNOR2_X1  g773(.A(new_n1197), .B(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(new_n996), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n1003), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1003), .A2(new_n1009), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1203), .B(KEYINPUT48), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1008), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1202), .A2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(KEYINPUT127), .B1(new_n1199), .B2(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n1197), .B(KEYINPUT47), .ZN(new_n1208));
  AND2_X1   g783(.A1(new_n1202), .A2(new_n1205), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT127), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1207), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1189), .A2(new_n1212), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g788(.A1(G227), .A2(new_n460), .ZN(new_n1215));
  NAND3_X1  g789(.A1(new_n718), .A2(new_n723), .A3(new_n1215), .ZN(new_n1216));
  AOI21_X1  g790(.A(new_n1216), .B1(new_n678), .B2(new_n681), .ZN(new_n1217));
  OAI211_X1 g791(.A(new_n1217), .B(new_n916), .C1(new_n982), .C2(new_n983), .ZN(G225));
  INV_X1    g792(.A(G225), .ZN(G308));
endmodule


