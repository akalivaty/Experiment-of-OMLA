//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 1 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007;
  INV_X1    g000(.A(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G217), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT69), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(G128), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT23), .A3(G119), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n194), .B(new_n196), .C1(G119), .C2(new_n195), .ZN(new_n197));
  XNOR2_X1  g011(.A(G119), .B(G128), .ZN(new_n198));
  XOR2_X1   g012(.A(KEYINPUT24), .B(G110), .Z(new_n199));
  AOI22_X1  g013(.A1(new_n197), .A2(G110), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G140), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G125), .ZN(new_n202));
  INV_X1    g016(.A(G125), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G140), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT16), .ZN(new_n205));
  OR3_X1    g019(.A1(new_n203), .A2(KEYINPUT16), .A3(G140), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G146), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(G146), .B1(new_n205), .B2(new_n206), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n200), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  OAI22_X1  g024(.A1(new_n197), .A2(G110), .B1(new_n198), .B2(new_n199), .ZN(new_n211));
  AND2_X1   g025(.A1(new_n202), .A2(new_n204), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT64), .B(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n211), .A2(new_n207), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n210), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(G221), .A2(G234), .ZN(new_n217));
  OR3_X1    g031(.A1(new_n217), .A2(KEYINPUT70), .A3(G953), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT22), .B(G137), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT70), .B1(new_n217), .B2(G953), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n219), .B1(new_n218), .B2(new_n220), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n216), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n223), .B1(new_n210), .B2(new_n215), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n191), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT25), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI211_X1 g043(.A(KEYINPUT25), .B(new_n191), .C1(new_n225), .C2(new_n226), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n190), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n216), .B(new_n224), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n189), .A2(G902), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  XOR2_X1   g049(.A(KEYINPUT26), .B(G101), .Z(new_n236));
  NOR2_X1   g050(.A1(G237), .A2(G953), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G210), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n236), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(G134), .B(G137), .ZN(new_n242));
  INV_X1    g056(.A(G131), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT65), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT11), .ZN(new_n245));
  INV_X1    g059(.A(G134), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n245), .B1(new_n246), .B2(G137), .ZN(new_n247));
  INV_X1    g061(.A(G137), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(KEYINPUT11), .A3(G134), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n246), .A2(G137), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n247), .A2(new_n249), .A3(new_n243), .A4(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT65), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n246), .A2(G137), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n248), .A2(G134), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n252), .B(G131), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n244), .A2(new_n251), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G146), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G143), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n258), .B1(new_n213), .B2(G143), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT1), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n260), .B1(new_n213), .B2(G143), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n259), .B1(new_n261), .B2(new_n195), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n257), .A2(KEYINPUT64), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT64), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G146), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n263), .A2(new_n265), .A3(G143), .ZN(new_n266));
  INV_X1    g080(.A(G143), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G146), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n195), .A2(KEYINPUT1), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n266), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n256), .B1(new_n262), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n247), .A2(new_n249), .A3(new_n250), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G131), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n273), .A2(new_n251), .ZN(new_n274));
  AND2_X1   g088(.A1(KEYINPUT0), .A2(G128), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n266), .A2(new_n275), .A3(new_n268), .ZN(new_n276));
  INV_X1    g090(.A(new_n258), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n263), .A2(new_n265), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n277), .B1(new_n278), .B2(new_n267), .ZN(new_n279));
  NOR2_X1   g093(.A1(KEYINPUT0), .A2(G128), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n275), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n276), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n274), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n271), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT28), .ZN(new_n286));
  XOR2_X1   g100(.A(KEYINPUT2), .B(G113), .Z(new_n287));
  INV_X1    g101(.A(KEYINPUT66), .ZN(new_n288));
  XNOR2_X1  g102(.A(G116), .B(G119), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n193), .A2(G116), .ZN(new_n291));
  INV_X1    g105(.A(G116), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G119), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT2), .B(G113), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n294), .A2(new_n295), .A3(KEYINPUT66), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n290), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT67), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n290), .A2(new_n296), .A3(KEYINPUT67), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n285), .A2(new_n286), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n273), .A2(new_n251), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n303), .B(new_n276), .C1(new_n279), .C2(new_n282), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n195), .B1(new_n266), .B2(KEYINPUT1), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n270), .B1(new_n305), .B2(new_n279), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n244), .A2(new_n251), .A3(new_n255), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n301), .A2(new_n304), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT28), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n302), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n308), .A2(new_n304), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n297), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n241), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT30), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n308), .A2(new_n304), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n315), .B1(new_n308), .B2(new_n304), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n297), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(new_n309), .A3(new_n241), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT31), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n309), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT30), .B1(new_n271), .B2(new_n284), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n308), .A2(new_n304), .A3(new_n315), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n322), .B1(new_n325), .B2(new_n297), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n326), .A2(KEYINPUT31), .A3(new_n241), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n314), .B1(new_n321), .B2(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(G472), .A2(G902), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT32), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n311), .A2(new_n313), .ZN(new_n332));
  INV_X1    g146(.A(new_n241), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(KEYINPUT31), .B1(new_n326), .B2(new_n241), .ZN(new_n335));
  AND4_X1   g149(.A1(KEYINPUT31), .A2(new_n318), .A3(new_n309), .A4(new_n241), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT32), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(new_n338), .A3(new_n329), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n331), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n318), .A2(new_n309), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n333), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT29), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n342), .B(new_n343), .C1(new_n332), .C2(new_n333), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n285), .A2(new_n301), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n345), .B1(new_n310), .B2(new_n302), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n333), .A2(new_n343), .ZN(new_n347));
  AOI21_X1  g161(.A(G902), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G472), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n235), .B1(new_n340), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(G214), .B1(G237), .B2(G902), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G101), .ZN(new_n354));
  INV_X1    g168(.A(G107), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n355), .A2(G104), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT71), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n357), .A2(KEYINPUT3), .ZN(new_n358));
  INV_X1    g172(.A(G104), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(G107), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n356), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT3), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(KEYINPUT71), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n362), .A2(KEYINPUT71), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n355), .A2(G104), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n354), .B1(new_n367), .B2(KEYINPUT72), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT72), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n361), .A2(new_n369), .A3(new_n366), .ZN(new_n370));
  XNOR2_X1  g184(.A(KEYINPUT73), .B(G101), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n361), .A2(new_n371), .A3(new_n366), .ZN(new_n372));
  AOI22_X1  g186(.A1(new_n368), .A2(new_n370), .B1(KEYINPUT4), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n357), .A2(KEYINPUT3), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n358), .B1(new_n360), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n359), .A2(G107), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n376), .B1(new_n363), .B2(new_n365), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT72), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n378), .A2(new_n370), .A3(KEYINPUT4), .A4(G101), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n297), .B1(new_n373), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n365), .B1(new_n356), .B2(KEYINPUT74), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT74), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n376), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(G101), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n372), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n294), .A2(new_n295), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n289), .A2(KEYINPUT5), .ZN(new_n388));
  OAI21_X1  g202(.A(G113), .B1(new_n291), .B2(KEYINPUT5), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n387), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(G110), .B(G122), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n381), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n393), .ZN(new_n395));
  INV_X1    g209(.A(new_n297), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n378), .A2(G101), .A3(new_n370), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n372), .A2(KEYINPUT4), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n396), .B1(new_n399), .B2(new_n379), .ZN(new_n400));
  INV_X1    g214(.A(new_n392), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n395), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT77), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n394), .A2(new_n402), .A3(new_n403), .A4(KEYINPUT6), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n394), .A2(new_n402), .A3(KEYINPUT6), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT6), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n406), .B(new_n395), .C1(new_n400), .C2(new_n401), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT77), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n404), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n262), .A2(new_n203), .A3(new_n270), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n283), .A2(G125), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G224), .ZN(new_n413));
  OR3_X1    g227(.A1(new_n413), .A2(KEYINPUT78), .A3(G953), .ZN(new_n414));
  OAI21_X1  g228(.A(KEYINPUT78), .B1(new_n413), .B2(G953), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  XOR2_X1   g230(.A(new_n416), .B(KEYINPUT79), .Z(new_n417));
  XNOR2_X1  g231(.A(new_n412), .B(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n409), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(G210), .B1(G237), .B2(G902), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n416), .A2(KEYINPUT81), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n422), .B1(new_n410), .B2(new_n411), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n414), .A2(KEYINPUT7), .A3(new_n415), .ZN(new_n424));
  OR2_X1    g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n424), .ZN(new_n426));
  XOR2_X1   g240(.A(new_n393), .B(KEYINPUT8), .Z(new_n427));
  NAND2_X1  g241(.A1(new_n372), .A2(new_n385), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n427), .B1(new_n428), .B2(new_n391), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n390), .A2(KEYINPUT80), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT80), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n389), .A2(new_n431), .B1(new_n289), .B2(KEYINPUT5), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n387), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n429), .B1(new_n428), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n425), .A2(new_n426), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n394), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n191), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n420), .A2(new_n421), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n421), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n394), .A2(new_n402), .A3(KEYINPUT6), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(KEYINPUT77), .A3(new_n407), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n418), .B1(new_n442), .B2(new_n404), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n440), .B1(new_n443), .B2(new_n437), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n353), .B1(new_n439), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G469), .ZN(new_n446));
  INV_X1    g260(.A(new_n283), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n447), .B1(new_n373), .B2(new_n380), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n266), .A2(new_n268), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n195), .B1(new_n258), .B2(KEYINPUT1), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n270), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n386), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT10), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n428), .A2(new_n453), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n306), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n448), .A2(new_n274), .A3(new_n454), .A4(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(G110), .B(G140), .ZN(new_n458));
  INV_X1    g272(.A(G227), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n459), .A2(G953), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n458), .B(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT75), .B1(new_n386), .B2(new_n306), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT75), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n428), .A2(new_n262), .A3(new_n465), .A4(new_n270), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n464), .A2(new_n452), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n303), .ZN(new_n468));
  AND2_X1   g282(.A1(KEYINPUT76), .A2(KEYINPUT12), .ZN(new_n469));
  NOR2_X1   g283(.A1(KEYINPUT76), .A2(KEYINPUT12), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n467), .B(new_n303), .C1(KEYINPUT76), .C2(KEYINPUT12), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n463), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n454), .A2(new_n456), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n283), .B1(new_n399), .B2(new_n379), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n303), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n462), .B1(new_n476), .B2(new_n457), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n446), .B(new_n191), .C1(new_n473), .C2(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n474), .A2(new_n475), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n461), .B1(new_n479), .B2(new_n274), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n476), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n471), .A2(new_n472), .B1(new_n274), .B2(new_n479), .ZN(new_n482));
  OAI211_X1 g296(.A(G469), .B(new_n481), .C1(new_n482), .C2(new_n462), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n446), .A2(new_n191), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n478), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  XNOR2_X1  g300(.A(KEYINPUT9), .B(G234), .ZN(new_n487));
  OAI21_X1  g301(.A(G221), .B1(new_n487), .B2(G902), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  XOR2_X1   g303(.A(G113), .B(G122), .Z(new_n490));
  XOR2_X1   g304(.A(KEYINPUT83), .B(G104), .Z(new_n491));
  XOR2_X1   g305(.A(new_n490), .B(new_n491), .Z(new_n492));
  AND3_X1   g306(.A1(new_n237), .A2(G143), .A3(G214), .ZN(new_n493));
  AOI21_X1  g307(.A(G143), .B1(new_n237), .B2(G214), .ZN(new_n494));
  OAI21_X1  g308(.A(G131), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n237), .A2(G214), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n267), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n237), .A2(G143), .A3(G214), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(new_n243), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT17), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n495), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT84), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n208), .A2(new_n209), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT84), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n495), .A2(new_n499), .A3(new_n504), .A4(new_n500), .ZN(new_n505));
  OR2_X1    g319(.A1(new_n495), .A2(new_n500), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n502), .A2(new_n503), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n214), .B1(new_n257), .B2(new_n212), .ZN(new_n508));
  OAI211_X1 g322(.A(KEYINPUT18), .B(G131), .C1(new_n493), .C2(new_n494), .ZN(new_n509));
  NAND2_X1  g323(.A1(KEYINPUT18), .A2(G131), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n497), .A2(new_n498), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n508), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n492), .B1(new_n507), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n507), .A2(new_n512), .A3(new_n492), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT85), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n507), .A2(KEYINPUT85), .A3(new_n512), .A4(new_n492), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n513), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(G475), .B1(new_n518), .B2(G902), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT20), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n516), .A2(new_n517), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n495), .A2(new_n499), .ZN(new_n522));
  AND2_X1   g336(.A1(KEYINPUT82), .A2(KEYINPUT19), .ZN(new_n523));
  NOR2_X1   g337(.A1(KEYINPUT82), .A2(KEYINPUT19), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n212), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n525), .B1(new_n212), .B2(new_n524), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n207), .B(new_n522), .C1(new_n526), .C2(new_n278), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n527), .A2(new_n512), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n528), .A2(new_n492), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n521), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(G475), .A2(G902), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n520), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n529), .B1(new_n516), .B2(new_n517), .ZN(new_n534));
  INV_X1    g348(.A(new_n532), .ZN(new_n535));
  NOR3_X1   g349(.A1(new_n534), .A2(KEYINPUT20), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n519), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n267), .A2(G128), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n195), .A2(G143), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(new_n539), .A3(new_n246), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n292), .A2(G122), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n292), .A2(G122), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n543), .A2(new_n355), .ZN(new_n544));
  NOR3_X1   g358(.A1(new_n541), .A2(new_n542), .A3(G107), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n540), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(KEYINPUT13), .B1(new_n267), .B2(G128), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n547), .B(KEYINPUT86), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT13), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n548), .B(new_n539), .C1(new_n549), .C2(new_n538), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n546), .B1(new_n550), .B2(G134), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(G217), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n487), .A2(new_n553), .A3(G953), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(KEYINPUT89), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT14), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n542), .B1(new_n541), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n292), .A2(G122), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n558), .A2(KEYINPUT87), .A3(KEYINPUT14), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(KEYINPUT87), .B1(new_n558), .B2(KEYINPUT14), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n557), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n562), .A2(KEYINPUT88), .A3(G107), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(KEYINPUT88), .B1(new_n562), .B2(G107), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n538), .A2(new_n539), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G134), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n540), .ZN(new_n569));
  INV_X1    g383(.A(new_n545), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n552), .B(new_n555), .C1(new_n566), .C2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n555), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n562), .A2(G107), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT88), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n571), .B1(new_n576), .B2(new_n563), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n573), .B1(new_n577), .B2(new_n551), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n572), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n579), .A2(KEYINPUT91), .A3(new_n191), .ZN(new_n580));
  INV_X1    g394(.A(G478), .ZN(new_n581));
  NOR2_X1   g395(.A1(KEYINPUT90), .A2(KEYINPUT15), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(KEYINPUT90), .A2(KEYINPUT15), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n581), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n580), .B(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(G234), .A2(G237), .ZN(new_n587));
  INV_X1    g401(.A(G953), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(G952), .A3(new_n588), .ZN(new_n589));
  XOR2_X1   g403(.A(KEYINPUT21), .B(G898), .Z(new_n590));
  NAND3_X1  g404(.A1(new_n587), .A2(G902), .A3(G953), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(KEYINPUT92), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n537), .A2(new_n586), .A3(new_n594), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n351), .A2(new_n445), .A3(new_n489), .A4(new_n595), .ZN(new_n596));
  XOR2_X1   g410(.A(new_n596), .B(new_n371), .Z(G3));
  NAND3_X1  g411(.A1(new_n579), .A2(new_n581), .A3(new_n191), .ZN(new_n598));
  NAND2_X1  g412(.A1(G478), .A2(G902), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT33), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n579), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n572), .A2(new_n578), .A3(KEYINPUT33), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n600), .B1(G478), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n537), .A2(new_n593), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n421), .B1(new_n420), .B2(new_n438), .ZN(new_n607));
  AOI211_X1 g421(.A(new_n440), .B(new_n437), .C1(new_n409), .C2(new_n419), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n352), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(KEYINPUT93), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT93), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n445), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n606), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n486), .A2(new_n488), .ZN(new_n614));
  OAI21_X1  g428(.A(G472), .B1(new_n328), .B2(G902), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n337), .A2(new_n329), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n614), .A2(new_n235), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT34), .B(G104), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G6));
  XNOR2_X1  g435(.A(new_n519), .B(KEYINPUT94), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n531), .A2(new_n520), .A3(new_n532), .ZN(new_n623));
  OAI21_X1  g437(.A(KEYINPUT20), .B1(new_n534), .B2(new_n535), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n627), .A2(new_n586), .A3(new_n593), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n610), .B2(new_n612), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n618), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT35), .B(G107), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G9));
  NAND2_X1  g446(.A1(new_n229), .A2(new_n230), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n189), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT95), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n216), .B1(KEYINPUT36), .B2(new_n223), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n223), .A2(KEYINPUT36), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n637), .A2(new_n210), .A3(new_n215), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n233), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n635), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n636), .A2(KEYINPUT95), .A3(new_n233), .A4(new_n638), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT96), .B1(new_n634), .B2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT96), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n231), .A2(new_n643), .A3(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n648), .A2(new_n615), .A3(new_n616), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n649), .A2(new_n489), .A3(new_n445), .A4(new_n595), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT37), .B(G110), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G12));
  NAND2_X1  g466(.A1(new_n610), .A2(new_n612), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n331), .A2(new_n339), .B1(G472), .B2(new_n349), .ZN(new_n654));
  INV_X1    g468(.A(new_n648), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n654), .A2(new_n614), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n580), .B(new_n585), .Z(new_n657));
  OR2_X1    g471(.A1(new_n591), .A2(G900), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n589), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n626), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n653), .A2(new_n656), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G128), .ZN(G30));
  XNOR2_X1  g477(.A(new_n659), .B(KEYINPUT39), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n489), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(KEYINPUT40), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT40), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n439), .A2(new_n444), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n537), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n657), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n634), .A2(new_n644), .ZN(new_n676));
  INV_X1    g490(.A(G472), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n333), .B1(new_n345), .B2(new_n322), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n319), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n677), .B1(new_n679), .B2(new_n191), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n680), .B1(new_n331), .B2(new_n339), .ZN(new_n681));
  NOR4_X1   g495(.A1(new_n675), .A2(new_n353), .A3(new_n676), .A4(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n667), .A2(new_n669), .A3(new_n672), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G143), .ZN(G45));
  NAND3_X1  g498(.A1(new_n537), .A2(new_n605), .A3(new_n659), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n653), .A2(new_n656), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G146), .ZN(G48));
  NAND2_X1  g502(.A1(new_n340), .A2(new_n350), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n467), .A2(new_n303), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n469), .A2(new_n470), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n472), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n476), .A2(new_n457), .ZN(new_n693));
  AOI22_X1  g507(.A1(new_n692), .A2(new_n480), .B1(new_n693), .B2(new_n461), .ZN(new_n694));
  OAI21_X1  g508(.A(G469), .B1(new_n694), .B2(G902), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(new_n488), .A3(new_n478), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(KEYINPUT98), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT98), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n695), .A2(new_n478), .A3(new_n698), .A4(new_n488), .ZN(new_n699));
  AND4_X1   g513(.A1(new_n689), .A2(new_n697), .A3(new_n234), .A4(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n613), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT41), .B(G113), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G15));
  NOR3_X1   g517(.A1(new_n626), .A2(new_n657), .A3(new_n594), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n700), .A2(new_n653), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G116), .ZN(G18));
  INV_X1    g520(.A(new_n696), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n689), .A2(new_n595), .A3(new_n648), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n653), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G119), .ZN(G21));
  AOI21_X1  g524(.A(new_n611), .B1(new_n670), .B2(new_n352), .ZN(new_n711));
  AOI211_X1 g525(.A(KEYINPUT93), .B(new_n353), .C1(new_n439), .C2(new_n444), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n674), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  XOR2_X1   g527(.A(KEYINPUT99), .B(G472), .Z(new_n714));
  OAI21_X1  g528(.A(new_n714), .B1(new_n328), .B2(G902), .ZN(new_n715));
  OAI22_X1  g529(.A1(new_n335), .A2(new_n336), .B1(new_n346), .B2(new_n241), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n329), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n235), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n719), .A2(new_n593), .A3(new_n697), .A4(new_n699), .ZN(new_n720));
  OAI21_X1  g534(.A(KEYINPUT100), .B1(new_n713), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n675), .B1(new_n610), .B2(new_n612), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT100), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n697), .A2(new_n699), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n715), .A2(new_n717), .A3(new_n234), .A4(new_n593), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n722), .A2(new_n723), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n721), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G122), .ZN(G24));
  AOI21_X1  g543(.A(new_n696), .B1(new_n610), .B2(new_n612), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n715), .A2(new_n676), .A3(new_n717), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n685), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G125), .ZN(G27));
  NAND3_X1  g548(.A1(new_n439), .A2(new_n444), .A3(new_n352), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(KEYINPUT101), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT101), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n439), .A2(new_n444), .A3(new_n737), .A4(new_n352), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n736), .A2(new_n489), .A3(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT102), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(KEYINPUT42), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n739), .A2(new_n351), .A3(new_n686), .A4(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n736), .A2(new_n351), .A3(new_n489), .A4(new_n738), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n741), .B1(new_n744), .B2(new_n685), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G131), .ZN(G33));
  INV_X1    g561(.A(new_n661), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n246), .ZN(G36));
  INV_X1    g564(.A(KEYINPUT105), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n673), .A2(new_n605), .ZN(new_n752));
  XOR2_X1   g566(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n753));
  AND2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT104), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(KEYINPUT43), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n751), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n752), .A2(new_n753), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n759), .B(KEYINPUT105), .C1(new_n752), .C2(new_n756), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n617), .A2(new_n676), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n758), .A2(KEYINPUT44), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT106), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n736), .A2(new_n738), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n762), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n763), .B1(new_n762), .B2(new_n765), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT103), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n481), .B1(new_n482), .B2(new_n462), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT45), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n446), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n772), .B1(new_n771), .B2(new_n770), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n485), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT46), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n773), .A2(KEYINPUT46), .A3(new_n485), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(new_n478), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n488), .ZN(new_n779));
  INV_X1    g593(.A(new_n664), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n769), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n758), .A2(new_n760), .A3(new_n761), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT44), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n778), .A2(KEYINPUT103), .A3(new_n488), .A4(new_n664), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n781), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n768), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(new_n248), .ZN(G39));
  NOR4_X1   g602(.A1(new_n764), .A2(new_n689), .A3(new_n234), .A4(new_n685), .ZN(new_n789));
  XNOR2_X1  g603(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n778), .A2(new_n488), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n790), .B1(new_n778), .B2(new_n488), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n789), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G140), .ZN(G42));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n795));
  AND4_X1   g609(.A1(new_n657), .A2(new_n622), .A3(new_n625), .A4(new_n659), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n796), .A2(new_n736), .A3(new_n738), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT110), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT110), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n796), .A2(new_n736), .A3(new_n799), .A4(new_n738), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n798), .A2(new_n656), .A3(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n736), .A2(new_n732), .A3(new_n489), .A4(new_n738), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n802), .B1(new_n744), .B2(new_n748), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n746), .A2(new_n801), .A3(new_n804), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n713), .A2(KEYINPUT100), .A3(new_n720), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n723), .B1(new_n722), .B2(new_n726), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n657), .A2(new_n537), .A3(new_n594), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n615), .A2(new_n616), .A3(new_n234), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n489), .A2(new_n445), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n650), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n701), .A2(new_n705), .A3(new_n812), .A4(new_n709), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n808), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT108), .B1(new_n609), .B2(new_n606), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT108), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n537), .A2(new_n605), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n445), .A2(new_n816), .A3(new_n817), .A4(new_n593), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n815), .A2(new_n618), .A3(new_n818), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n819), .A2(KEYINPUT109), .A3(new_n596), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT109), .B1(new_n819), .B2(new_n596), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n653), .B(new_n656), .C1(new_n661), .C2(new_n686), .ZN(new_n823));
  XOR2_X1   g637(.A(new_n659), .B(KEYINPUT111), .Z(new_n824));
  OR2_X1    g638(.A1(new_n676), .A2(new_n824), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n614), .A2(new_n681), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n653), .A2(new_n674), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n823), .A2(new_n733), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(KEYINPUT112), .A3(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n805), .A2(new_n814), .A3(new_n822), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n828), .A2(new_n829), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n828), .A2(KEYINPUT112), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n823), .A2(new_n733), .A3(KEYINPUT52), .A4(new_n827), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n795), .B1(new_n831), .B2(new_n835), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n629), .A2(new_n700), .B1(new_n730), .B2(new_n708), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n650), .A2(new_n811), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n838), .B1(new_n613), .B2(new_n700), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n728), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  AND4_X1   g654(.A1(new_n351), .A2(new_n736), .A3(new_n489), .A4(new_n738), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n742), .B1(new_n841), .B2(new_n686), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n744), .A2(new_n685), .A3(new_n741), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n804), .B(new_n801), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n820), .A2(new_n821), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n840), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n832), .A2(new_n834), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(KEYINPUT53), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n836), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT113), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n849), .A2(new_n850), .A3(KEYINPUT54), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n846), .A2(KEYINPUT53), .A3(new_n852), .A4(new_n830), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n847), .A2(new_n805), .A3(new_n814), .A4(new_n822), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n795), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n853), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n851), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n856), .B1(new_n836), .B2(new_n848), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n859), .A2(new_n850), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT114), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n853), .A2(new_n855), .A3(new_n856), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n862), .B1(new_n850), .B2(new_n859), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT114), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n849), .A2(KEYINPUT54), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT113), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n764), .A2(new_n696), .ZN(new_n868));
  INV_X1    g682(.A(new_n681), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n869), .A2(new_n235), .A3(new_n589), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT116), .Z(new_n872));
  INV_X1    g686(.A(new_n604), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n873), .A2(new_n581), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n872), .B(new_n673), .C1(new_n874), .C2(new_n600), .ZN(new_n875));
  INV_X1    g689(.A(new_n757), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n589), .B1(new_n876), .B2(new_n759), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n868), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n878), .A2(new_n731), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n877), .A2(new_n719), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n672), .A2(new_n352), .A3(new_n696), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT50), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n880), .A2(KEYINPUT50), .A3(new_n881), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n879), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n875), .A2(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n880), .A2(new_n765), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n791), .A2(new_n792), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n695), .A2(new_n478), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n891), .A2(new_n488), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n888), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n887), .A2(KEYINPUT51), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n872), .A2(new_n817), .ZN(new_n895));
  INV_X1    g709(.A(new_n351), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n878), .A2(new_n896), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT48), .Z(new_n898));
  INV_X1    g712(.A(G952), .ZN(new_n899));
  AOI211_X1 g713(.A(new_n899), .B(G953), .C1(new_n880), .C2(new_n730), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n894), .A2(new_n895), .A3(new_n898), .A4(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n892), .B1(new_n889), .B2(KEYINPUT115), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n902), .B1(KEYINPUT115), .B2(new_n889), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n888), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT51), .B1(new_n887), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n901), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n861), .A2(new_n867), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n899), .A2(new_n588), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n752), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n910), .A2(new_n234), .A3(new_n352), .A4(new_n488), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n891), .B(KEYINPUT49), .ZN(new_n912));
  OR4_X1    g726(.A1(new_n672), .A2(new_n911), .A3(new_n869), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n909), .A2(new_n913), .ZN(G75));
  NAND2_X1  g728(.A1(new_n853), .A2(new_n855), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n916), .A2(new_n191), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(G210), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n409), .B(new_n419), .ZN(new_n919));
  XNOR2_X1  g733(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n919), .B(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT118), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n922), .A2(KEYINPUT56), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n918), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n921), .B1(new_n918), .B2(new_n923), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n588), .A2(G952), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(G51));
  XNOR2_X1  g741(.A(new_n484), .B(KEYINPUT57), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n916), .A2(new_n856), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n928), .B1(new_n929), .B2(new_n862), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(new_n477), .B2(new_n473), .ZN(new_n931));
  OR3_X1    g745(.A1(new_n916), .A2(new_n191), .A3(new_n773), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n926), .B1(new_n931), .B2(new_n932), .ZN(G54));
  NAND3_X1  g747(.A1(new_n917), .A2(KEYINPUT58), .A3(G475), .ZN(new_n934));
  OR3_X1    g748(.A1(new_n934), .A2(KEYINPUT119), .A3(new_n534), .ZN(new_n935));
  OAI21_X1  g749(.A(KEYINPUT119), .B1(new_n934), .B2(new_n534), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n926), .B1(new_n934), .B2(new_n534), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(G60));
  XNOR2_X1  g752(.A(new_n599), .B(KEYINPUT59), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n873), .B(new_n939), .C1(new_n929), .C2(new_n862), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n940), .B1(G952), .B2(new_n588), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n858), .A2(new_n860), .A3(KEYINPUT114), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n864), .B1(new_n863), .B2(new_n866), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n939), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n941), .B1(new_n944), .B2(new_n604), .ZN(G63));
  NAND2_X1  g759(.A1(G217), .A2(G902), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT120), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT60), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n915), .A2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n232), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n926), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n949), .A2(new_n639), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT121), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n949), .A2(KEYINPUT121), .A3(new_n639), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n951), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT61), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI211_X1 g772(.A(KEYINPUT61), .B(new_n951), .C1(new_n954), .C2(new_n955), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(G66));
  AOI21_X1  g774(.A(new_n588), .B1(new_n590), .B2(G224), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n814), .A2(new_n822), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n961), .B1(new_n962), .B2(new_n588), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n442), .B(new_n404), .C1(G898), .C2(new_n588), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n963), .B(new_n964), .Z(G69));
  XOR2_X1   g779(.A(new_n325), .B(KEYINPUT122), .Z(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(new_n526), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n793), .B1(new_n768), .B2(new_n786), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n781), .A2(new_n351), .A3(new_n722), .A4(new_n785), .ZN(new_n969));
  INV_X1    g783(.A(new_n749), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n823), .A2(new_n733), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n969), .A2(new_n746), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n588), .B1(new_n968), .B2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(G900), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(G953), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n973), .A2(KEYINPUT125), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(KEYINPUT125), .B1(new_n973), .B2(new_n975), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n967), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(G953), .B1(new_n459), .B2(new_n974), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT124), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n971), .A2(new_n683), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT62), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n817), .B1(new_n586), .B2(new_n673), .ZN(new_n983));
  NOR4_X1   g797(.A1(new_n666), .A2(new_n764), .A3(new_n896), .A4(new_n983), .ZN(new_n984));
  OR3_X1    g798(.A1(new_n982), .A2(new_n968), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n588), .ZN(new_n986));
  INV_X1    g800(.A(new_n967), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT123), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(KEYINPUT123), .B1(new_n986), .B2(new_n987), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n978), .B(new_n980), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n980), .B1(new_n978), .B2(new_n988), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT126), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  AOI211_X1 g809(.A(KEYINPUT126), .B(new_n980), .C1(new_n978), .C2(new_n988), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n992), .B1(new_n995), .B2(new_n996), .ZN(G72));
  NAND2_X1  g811(.A1(G472), .A2(G902), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT63), .Z(new_n999));
  INV_X1    g813(.A(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(new_n849), .ZN(new_n1001));
  AOI211_X1 g815(.A(new_n1000), .B(new_n1001), .C1(new_n319), .C2(new_n342), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n999), .B1(new_n985), .B2(new_n962), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n326), .B(KEYINPUT127), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n1003), .A2(new_n241), .A3(new_n1004), .ZN(new_n1005));
  OR3_X1    g819(.A1(new_n968), .A2(new_n972), .A3(new_n962), .ZN(new_n1006));
  AOI211_X1 g820(.A(new_n241), .B(new_n1004), .C1(new_n1006), .C2(new_n999), .ZN(new_n1007));
  NOR4_X1   g821(.A1(new_n1002), .A2(new_n1005), .A3(new_n926), .A4(new_n1007), .ZN(G57));
endmodule


