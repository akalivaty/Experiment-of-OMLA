//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 1 1 1 1 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n568, new_n570, new_n571, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT66), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT67), .ZN(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G125), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n462), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(new_n469), .A3(G125), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g048(.A(G2105), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n475), .A2(G137), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  AND2_X1   g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n476), .B(KEYINPUT69), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n465), .A2(G2105), .ZN(new_n483));
  AOI22_X1  g058(.A1(new_n479), .A2(new_n482), .B1(G101), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n474), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G160));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n481), .A2(new_n480), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n471), .A2(KEYINPUT70), .ZN(new_n492));
  OAI21_X1  g067(.A(G2105), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G124), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n488), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n475), .B1(new_n491), .B2(new_n492), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n495), .B1(G136), .B2(new_n497), .ZN(new_n498));
  XNOR2_X1  g073(.A(new_n498), .B(KEYINPUT71), .ZN(G162));
  OAI21_X1  g074(.A(G2104), .B1(new_n475), .B2(G114), .ZN(new_n500));
  NOR2_X1   g075(.A1(G102), .A2(G2105), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(G126), .A2(G2105), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n503), .B1(new_n466), .B2(new_n467), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n475), .A2(G138), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n506), .B1(new_n489), .B2(new_n507), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n471), .A2(KEYINPUT4), .A3(G138), .A4(new_n475), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n505), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  NAND2_X1  g086(.A1(KEYINPUT72), .A2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(KEYINPUT73), .A3(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n515), .B1(KEYINPUT72), .B2(KEYINPUT5), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT5), .ZN(new_n517));
  OAI21_X1  g092(.A(G543), .B1(new_n517), .B2(KEYINPUT73), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n514), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n519), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(KEYINPUT6), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT6), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n526), .A2(new_n513), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G50), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT6), .B(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n519), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G88), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n522), .A2(new_n532), .ZN(G303));
  INV_X1    g108(.A(G303), .ZN(G166));
  NAND3_X1  g109(.A1(new_n519), .A2(G63), .A3(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(KEYINPUT74), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT74), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n519), .A2(new_n537), .A3(G63), .A4(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n529), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G51), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n512), .A2(KEYINPUT73), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n515), .A2(KEYINPUT5), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n545), .A2(G543), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n526), .B1(new_n547), .B2(new_n514), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n544), .B1(G89), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n539), .A2(new_n549), .ZN(G286));
  INV_X1    g125(.A(G286), .ZN(G168));
  AOI22_X1  g126(.A1(new_n548), .A2(G90), .B1(G52), .B2(new_n527), .ZN(new_n552));
  AND2_X1   g127(.A1(G77), .A2(G543), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n553), .B1(new_n519), .B2(G64), .ZN(new_n554));
  OAI21_X1  g129(.A(G651), .B1(new_n554), .B2(KEYINPUT75), .ZN(new_n555));
  INV_X1    g130(.A(G64), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n556), .B1(new_n547), .B2(new_n514), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT75), .ZN(new_n558));
  NOR3_X1   g133(.A1(new_n557), .A2(new_n558), .A3(new_n553), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n552), .B1(new_n555), .B2(new_n559), .ZN(G301));
  INV_X1    g135(.A(G301), .ZN(G171));
  AOI22_X1  g136(.A1(new_n548), .A2(G81), .B1(G43), .B2(new_n527), .ZN(new_n562));
  AND2_X1   g137(.A1(G68), .A2(G543), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n563), .B1(new_n519), .B2(G56), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n562), .B1(new_n521), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n568));
  XOR2_X1   g143(.A(new_n568), .B(KEYINPUT76), .Z(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n573), .B1(new_n547), .B2(new_n514), .ZN(new_n574));
  AND2_X1   g149(.A1(G78), .A2(G543), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n548), .A2(G91), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n523), .A2(new_n525), .A3(G53), .A4(G543), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT77), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT9), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n578), .A2(new_n579), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n529), .A2(KEYINPUT77), .A3(G53), .A4(G543), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n582), .A2(new_n583), .A3(KEYINPUT9), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n576), .A2(new_n577), .A3(new_n581), .A4(new_n584), .ZN(G299));
  INV_X1    g160(.A(G74), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n547), .A2(new_n586), .A3(new_n514), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n587), .A2(G651), .B1(new_n527), .B2(G49), .ZN(new_n588));
  AOI21_X1  g163(.A(KEYINPUT78), .B1(new_n548), .B2(G87), .ZN(new_n589));
  AND4_X1   g164(.A1(KEYINPUT78), .A2(new_n519), .A3(G87), .A4(new_n529), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(G288));
  NAND2_X1  g166(.A1(new_n527), .A2(G48), .ZN(new_n592));
  INV_X1    g167(.A(G86), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n519), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n594));
  OAI221_X1 g169(.A(new_n592), .B1(new_n530), .B2(new_n593), .C1(new_n594), .C2(new_n521), .ZN(G305));
  AOI22_X1  g170(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(new_n521), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n527), .A2(G47), .ZN(new_n598));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n530), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n527), .A2(G54), .ZN(new_n604));
  INV_X1    g179(.A(G66), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n605), .B1(new_n547), .B2(new_n514), .ZN(new_n606));
  AND2_X1   g181(.A1(G79), .A2(G543), .ZN(new_n607));
  OAI21_X1  g182(.A(G651), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g183(.A(KEYINPUT10), .B1(new_n548), .B2(G92), .ZN(new_n609));
  AND4_X1   g184(.A1(KEYINPUT10), .A2(new_n519), .A3(G92), .A4(new_n529), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n604), .B(new_n608), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n603), .B1(new_n612), .B2(G868), .ZN(G284));
  OAI21_X1  g188(.A(new_n603), .B1(new_n612), .B2(G868), .ZN(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  INV_X1    g190(.A(G299), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(G868), .B2(new_n616), .ZN(G297));
  OAI21_X1  g192(.A(new_n615), .B1(G868), .B2(new_n616), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n612), .B1(new_n619), .B2(G860), .ZN(G148));
  NAND2_X1  g195(.A1(new_n612), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n566), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n471), .A2(new_n483), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT12), .Z(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT13), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2100), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n497), .A2(G135), .ZN(new_n629));
  INV_X1    g204(.A(new_n493), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G123), .ZN(new_n631));
  OR2_X1    g206(.A1(G99), .A2(G2105), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n632), .B(G2104), .C1(G111), .C2(new_n475), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n629), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(G2096), .Z(new_n635));
  NAND2_X1  g210(.A1(new_n628), .A2(new_n635), .ZN(G156));
  XNOR2_X1  g211(.A(G2451), .B(G2454), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2443), .B(G2446), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(KEYINPUT15), .B(G2435), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2430), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  AND2_X1   g221(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n644), .A2(new_n646), .ZN(new_n648));
  XOR2_X1   g223(.A(KEYINPUT79), .B(KEYINPUT14), .Z(new_n649));
  NOR3_X1   g224(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n642), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n642), .A2(new_n650), .ZN(new_n652));
  AND3_X1   g227(.A1(new_n651), .A2(G14), .A3(new_n652), .ZN(G401));
  XOR2_X1   g228(.A(G2067), .B(G2678), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT80), .ZN(new_n655));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  XNOR2_X1  g231(.A(G2084), .B(G2090), .ZN(new_n657));
  NOR3_X1   g232(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT18), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n655), .A2(new_n656), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n656), .B(KEYINPUT17), .ZN(new_n661));
  OAI211_X1 g236(.A(new_n660), .B(new_n657), .C1(new_n655), .C2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n657), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n661), .A2(new_n655), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n659), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2096), .B(G2100), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT81), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n665), .B(new_n667), .ZN(G227));
  XOR2_X1   g243(.A(G1971), .B(G1976), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  XOR2_X1   g245(.A(G1956), .B(G2474), .Z(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n671), .A2(new_n672), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n675), .A2(new_n673), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n670), .A2(new_n675), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n678));
  OAI221_X1 g253(.A(new_n674), .B1(new_n676), .B2(new_n670), .C1(new_n677), .C2(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n677), .B2(new_n678), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT83), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G1981), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n680), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT84), .B(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(G229));
  INV_X1    g264(.A(KEYINPUT90), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(KEYINPUT36), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT91), .Z(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(G288), .A2(KEYINPUT88), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT88), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n695), .B(new_n588), .C1(new_n589), .C2(new_n590), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  MUX2_X1   g272(.A(G23), .B(new_n697), .S(G16), .Z(new_n698));
  OR2_X1    g273(.A1(new_n698), .A2(KEYINPUT33), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(KEYINPUT33), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G1976), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G6), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n594), .A2(new_n521), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n592), .B1(new_n530), .B2(new_n593), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n705), .B1(new_n708), .B2(new_n704), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT32), .B(G1981), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT87), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n704), .A2(G22), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G166), .B2(new_n704), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G1971), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n711), .A2(new_n712), .ZN(new_n717));
  NOR3_X1   g292(.A1(new_n713), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n699), .A2(G1976), .A3(new_n700), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n703), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT89), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n703), .A2(new_n718), .A3(KEYINPUT89), .A4(new_n719), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n722), .A2(KEYINPUT34), .A3(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G25), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n497), .A2(G131), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n630), .A2(G119), .ZN(new_n728));
  OR2_X1    g303(.A1(G95), .A2(G2105), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n729), .B(G2104), .C1(G107), .C2(new_n475), .ZN(new_n730));
  AND3_X1   g305(.A1(new_n727), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n726), .B1(new_n731), .B2(new_n725), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT85), .Z(new_n733));
  XOR2_X1   g308(.A(KEYINPUT35), .B(G1991), .Z(new_n734));
  OR2_X1    g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  AND3_X1   g311(.A1(new_n735), .A2(KEYINPUT86), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(KEYINPUT86), .B1(new_n735), .B2(new_n736), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n704), .A2(G24), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n601), .B2(new_n704), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G1986), .ZN(new_n741));
  NOR3_X1   g316(.A1(new_n737), .A2(new_n738), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n724), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(KEYINPUT34), .B1(new_n722), .B2(new_n723), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n693), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(new_n744), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n746), .A2(new_n692), .A3(new_n724), .A4(new_n742), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n497), .A2(G141), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n630), .A2(G129), .ZN(new_n749));
  NAND3_X1  g324(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT26), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n752), .A2(new_n753), .B1(G105), .B2(new_n483), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n748), .A2(new_n749), .A3(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n756), .A2(new_n725), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n725), .B2(G32), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT27), .B(G1996), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G28), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n761), .A2(KEYINPUT30), .ZN(new_n762));
  AOI21_X1  g337(.A(G29), .B1(new_n761), .B2(KEYINPUT30), .ZN(new_n763));
  OR2_X1    g338(.A1(KEYINPUT31), .A2(G11), .ZN(new_n764));
  NAND2_X1  g339(.A1(KEYINPUT31), .A2(G11), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n762), .A2(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n634), .B2(new_n725), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n725), .A2(G27), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G164), .B2(new_n725), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G2078), .ZN(new_n770));
  NOR3_X1   g345(.A1(new_n760), .A2(new_n767), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n704), .A2(G21), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G168), .B2(new_n704), .ZN(new_n773));
  INV_X1    g348(.A(G1966), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(KEYINPUT24), .A2(G34), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT24), .ZN(new_n777));
  INV_X1    g352(.A(G34), .ZN(new_n778));
  AOI21_X1  g353(.A(G29), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n485), .A2(G29), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(G2084), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT94), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n771), .A2(new_n775), .A3(new_n783), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n725), .A2(G33), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n497), .A2(G139), .ZN(new_n786));
  NAND2_X1  g361(.A1(G115), .A2(G2104), .ZN(new_n787));
  INV_X1    g362(.A(G127), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n489), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n475), .B1(new_n789), .B2(KEYINPUT93), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(KEYINPUT93), .B2(new_n789), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT25), .Z(new_n793));
  NAND3_X1  g368(.A1(new_n786), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n785), .B1(new_n794), .B2(G29), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n795), .A2(new_n442), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n795), .A2(new_n442), .ZN(new_n797));
  AOI211_X1 g372(.A(new_n796), .B(new_n797), .C1(new_n758), .C2(new_n759), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n780), .A2(new_n781), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT95), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n704), .A2(G5), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G171), .B2(new_n704), .ZN(new_n802));
  INV_X1    g377(.A(G1961), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n798), .A2(new_n800), .A3(new_n804), .ZN(new_n805));
  OR3_X1    g380(.A1(new_n784), .A2(KEYINPUT96), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(KEYINPUT96), .B1(new_n784), .B2(new_n805), .ZN(new_n807));
  OR2_X1    g382(.A1(G104), .A2(G2105), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n808), .B(G2104), .C1(G116), .C2(new_n475), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n630), .B2(G128), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n497), .A2(G140), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(G29), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT92), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n725), .A2(G26), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT28), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(G2067), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n725), .A2(G35), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G162), .B2(new_n725), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT29), .B(G2090), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n612), .A2(new_n704), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(G4), .B2(new_n704), .ZN(new_n825));
  INV_X1    g400(.A(G1348), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n704), .A2(G20), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT23), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n616), .B2(new_n704), .ZN(new_n830));
  INV_X1    g405(.A(G1956), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n825), .A2(new_n826), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n704), .A2(G19), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n566), .B2(new_n704), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(G1341), .Z(new_n836));
  NAND4_X1  g411(.A1(new_n827), .A2(new_n832), .A3(new_n833), .A4(new_n836), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n819), .A2(new_n823), .A3(new_n837), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n806), .A2(new_n807), .A3(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n745), .A2(new_n747), .A3(new_n839), .ZN(G150));
  INV_X1    g415(.A(G150), .ZN(G311));
  XNOR2_X1  g416(.A(KEYINPUT97), .B(G93), .ZN(new_n842));
  AOI22_X1  g417(.A1(new_n548), .A2(new_n842), .B1(G55), .B2(new_n527), .ZN(new_n843));
  INV_X1    g418(.A(G67), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(new_n547), .B2(new_n514), .ZN(new_n845));
  AND2_X1   g420(.A1(G80), .A2(G543), .ZN(new_n846));
  OAI21_X1  g421(.A(G651), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(G860), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT37), .Z(new_n850));
  NAND2_X1  g425(.A1(new_n565), .A2(new_n848), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n564), .A2(new_n521), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n852), .A2(new_n562), .A3(new_n847), .A4(new_n843), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT38), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n612), .A2(G559), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT39), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT98), .ZN(new_n860));
  INV_X1    g435(.A(G860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(new_n857), .B2(new_n858), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n850), .B1(new_n860), .B2(new_n862), .ZN(G145));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT99), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n865), .B1(new_n502), .B2(new_n504), .ZN(new_n866));
  INV_X1    g441(.A(new_n503), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(new_n481), .B2(new_n480), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n868), .B(KEYINPUT99), .C1(new_n501), .C2(new_n500), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n866), .A2(new_n869), .A3(new_n508), .A4(new_n509), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n811), .A2(new_n812), .A3(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n871), .B1(new_n811), .B2(new_n812), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n756), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n874), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n876), .A2(new_n872), .A3(new_n755), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n794), .B(KEYINPUT100), .Z(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n794), .A2(KEYINPUT100), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n875), .A2(new_n877), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n497), .A2(G142), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n630), .A2(G130), .ZN(new_n885));
  OR2_X1    g460(.A1(G106), .A2(G2105), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n886), .B(G2104), .C1(G118), .C2(new_n475), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(new_n626), .ZN(new_n889));
  INV_X1    g464(.A(new_n626), .ZN(new_n890));
  NAND4_X1  g465(.A1(new_n890), .A2(new_n884), .A3(new_n885), .A4(new_n887), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n889), .A2(new_n731), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n731), .B1(new_n889), .B2(new_n891), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n864), .B1(new_n883), .B2(new_n895), .ZN(new_n896));
  AOI211_X1 g471(.A(KEYINPUT101), .B(new_n894), .C1(new_n880), .C2(new_n882), .ZN(new_n897));
  OAI22_X1  g472(.A1(new_n896), .A2(new_n897), .B1(new_n895), .B2(new_n883), .ZN(new_n898));
  OR2_X1    g473(.A1(G162), .A2(new_n485), .ZN(new_n899));
  NAND2_X1  g474(.A1(G162), .A2(new_n485), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n634), .ZN(new_n902));
  INV_X1    g477(.A(new_n634), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n899), .A2(new_n903), .A3(new_n900), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(G37), .B1(new_n898), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n883), .A2(new_n895), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n907), .A2(KEYINPUT102), .ZN(new_n908));
  AOI22_X1  g483(.A1(new_n907), .A2(KEYINPUT102), .B1(new_n902), .B2(new_n904), .ZN(new_n909));
  OAI211_X1 g484(.A(new_n908), .B(new_n909), .C1(new_n896), .C2(new_n897), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT40), .ZN(G395));
  NAND3_X1  g487(.A1(new_n694), .A2(new_n601), .A3(new_n696), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n601), .B1(new_n694), .B2(new_n696), .ZN(new_n915));
  OAI21_X1  g490(.A(KEYINPUT104), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n915), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT104), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(new_n918), .A3(new_n913), .ZN(new_n919));
  XNOR2_X1  g494(.A(G303), .B(new_n708), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n916), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n920), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n922), .A2(new_n917), .A3(new_n918), .A4(new_n913), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT105), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(KEYINPUT106), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT42), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n925), .B(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT42), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT41), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n616), .A2(new_n611), .ZN(new_n933));
  INV_X1    g508(.A(new_n609), .ZN(new_n934));
  INV_X1    g509(.A(new_n610), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n608), .A2(new_n604), .ZN(new_n937));
  AOI21_X1  g512(.A(G299), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n932), .B1(new_n933), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n616), .A2(new_n611), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n936), .A2(new_n937), .A3(G299), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(new_n941), .A3(KEYINPUT41), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n941), .ZN(new_n944));
  XOR2_X1   g519(.A(new_n944), .B(KEYINPUT103), .Z(new_n945));
  XNOR2_X1  g520(.A(new_n621), .B(new_n854), .ZN(new_n946));
  MUX2_X1   g521(.A(new_n943), .B(new_n945), .S(new_n946), .Z(new_n947));
  AND3_X1   g522(.A1(new_n927), .A2(new_n931), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n947), .B1(new_n927), .B2(new_n931), .ZN(new_n949));
  OAI21_X1  g524(.A(G868), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n848), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n950), .B1(G868), .B2(new_n951), .ZN(G295));
  OAI21_X1  g527(.A(new_n950), .B1(G868), .B2(new_n951), .ZN(G331));
  INV_X1    g528(.A(G37), .ZN(new_n954));
  NOR2_X1   g529(.A1(G301), .A2(G286), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n558), .B1(new_n557), .B2(new_n553), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n519), .A2(G64), .ZN(new_n957));
  INV_X1    g532(.A(new_n553), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n957), .A2(KEYINPUT75), .A3(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n956), .A2(new_n959), .A3(G651), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n960), .A2(new_n552), .B1(new_n539), .B2(new_n549), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n854), .B1(new_n955), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT107), .ZN(new_n963));
  NAND2_X1  g538(.A1(G301), .A2(G286), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n960), .A2(new_n539), .A3(new_n549), .A4(new_n552), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n964), .A2(new_n851), .A3(new_n965), .A4(new_n853), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n962), .A2(new_n963), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n854), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n968), .A2(KEYINPUT107), .A3(new_n964), .A4(new_n965), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n967), .A2(new_n943), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT108), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n967), .A2(new_n943), .A3(new_n972), .A4(new_n969), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n962), .A2(new_n966), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n944), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n971), .A2(new_n973), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n954), .B1(new_n977), .B2(new_n924), .ZN(new_n978));
  AOI22_X1  g553(.A1(new_n970), .A2(KEYINPUT108), .B1(new_n944), .B2(new_n975), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n979), .A2(new_n973), .B1(new_n923), .B2(new_n921), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT43), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT109), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n983), .B(KEYINPUT43), .C1(new_n978), .C2(new_n980), .ZN(new_n984));
  INV_X1    g559(.A(new_n978), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT43), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n967), .A2(new_n969), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n945), .A2(new_n987), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n943), .A2(new_n974), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n924), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT110), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n992), .B(new_n924), .C1(new_n988), .C2(new_n989), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n985), .A2(new_n986), .A3(new_n991), .A4(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n982), .A2(new_n984), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT44), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AND4_X1   g572(.A1(KEYINPUT43), .A2(new_n985), .A3(new_n991), .A4(new_n993), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n978), .A2(new_n980), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(KEYINPUT43), .ZN(new_n1000));
  OAI21_X1  g575(.A(KEYINPUT44), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n997), .A2(new_n1001), .ZN(G397));
  INV_X1    g577(.A(G1384), .ZN(new_n1003));
  XOR2_X1   g578(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n1004));
  NAND3_X1  g579(.A1(new_n870), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT112), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n870), .A2(KEYINPUT112), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n474), .A2(new_n484), .A3(G40), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n510), .A2(new_n1003), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1010), .B1(KEYINPUT50), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT113), .B1(new_n1013), .B2(G2090), .ZN(new_n1014));
  OAI21_X1  g589(.A(G125), .B1(new_n481), .B2(new_n480), .ZN(new_n1015));
  AOI22_X1  g590(.A1(new_n1015), .A2(KEYINPUT68), .B1(G113), .B2(G2104), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n475), .B1(new_n1016), .B2(new_n472), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n483), .A2(G101), .ZN(new_n1018));
  INV_X1    g593(.A(new_n482), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT69), .B1(new_n471), .B2(new_n476), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1018), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G40), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n1017), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT45), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1011), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n870), .A2(KEYINPUT45), .A3(new_n1003), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1023), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G1971), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n1030));
  INV_X1    g605(.A(G2090), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1009), .A2(new_n1012), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1014), .A2(new_n1029), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(G303), .A2(G8), .ZN(new_n1036));
  XOR2_X1   g611(.A(new_n1036), .B(KEYINPUT55), .Z(new_n1037));
  NAND4_X1  g612(.A1(new_n1014), .A2(KEYINPUT114), .A3(new_n1029), .A4(new_n1032), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1035), .A2(G8), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1037), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1023), .B1(KEYINPUT50), .B2(new_n1011), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n870), .A2(new_n1003), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1043), .A2(new_n1004), .ZN(new_n1044));
  NOR3_X1   g619(.A1(new_n1041), .A2(new_n1044), .A3(G2090), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1045), .B1(new_n1028), .B2(new_n1027), .ZN(new_n1046));
  INV_X1    g621(.A(G8), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1040), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT115), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1043), .A2(new_n1023), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1049), .B1(new_n1050), .B2(G8), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1049), .B(G8), .C1(new_n1010), .C2(new_n1042), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  OR2_X1    g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT49), .ZN(new_n1055));
  NOR3_X1   g630(.A1(G305), .A2(KEYINPUT117), .A3(G1981), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n1057));
  INV_X1    g632(.A(G1981), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1057), .B1(new_n708), .B2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n708), .A2(new_n1058), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1055), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  OAI221_X1 g637(.A(KEYINPUT49), .B1(new_n1058), .B2(new_n708), .C1(new_n1056), .C2(new_n1059), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1054), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  XOR2_X1   g639(.A(KEYINPUT116), .B(G1976), .Z(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT52), .B1(G288), .B2(new_n1065), .ZN(new_n1066));
  OAI221_X1 g641(.A(new_n1066), .B1(new_n697), .B2(new_n702), .C1(new_n1051), .C2(new_n1053), .ZN(new_n1067));
  OAI22_X1  g642(.A1(new_n1051), .A2(new_n1053), .B1(new_n697), .B2(new_n702), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT52), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1064), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1039), .A2(new_n1048), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1009), .A2(new_n781), .A3(new_n1012), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT118), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1009), .A2(new_n1012), .A3(KEYINPUT118), .A4(new_n781), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT45), .B1(new_n870), .B2(new_n1003), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1076), .A2(new_n1010), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n510), .A2(KEYINPUT45), .A3(new_n1003), .ZN(new_n1078));
  AOI21_X1  g653(.A(G1966), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1074), .A2(G168), .A3(new_n1075), .A4(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1079), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1082));
  AOI21_X1  g657(.A(G168), .B1(new_n1082), .B2(new_n1075), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT51), .ZN(new_n1084));
  OAI211_X1 g659(.A(G8), .B(new_n1081), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1081), .A2(G8), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(KEYINPUT51), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1009), .A2(new_n1089), .A3(new_n1012), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1089), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n803), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1077), .A2(KEYINPUT53), .A3(new_n443), .A4(new_n1078), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1023), .A2(new_n1025), .A3(new_n443), .A4(new_n1026), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1094), .A2(KEYINPUT122), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1092), .A2(new_n1093), .A3(new_n1096), .A4(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g675(.A(G301), .B(KEYINPUT54), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1096), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1091), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1009), .A2(new_n1089), .A3(new_n1012), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1102), .B1(new_n1105), .B2(new_n803), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1026), .A2(KEYINPUT53), .A3(new_n443), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1101), .B1(new_n1077), .B2(new_n1107), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1100), .A2(new_n1101), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1071), .A2(KEYINPUT123), .A3(new_n1088), .A4(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT123), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1088), .A2(new_n1109), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1039), .A2(new_n1048), .A3(new_n1070), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n831), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1115));
  XNOR2_X1  g690(.A(G299), .B(KEYINPUT57), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g692(.A(KEYINPUT56), .B(G2072), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1023), .A2(new_n1026), .A3(new_n1025), .A4(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1115), .A2(new_n1117), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n826), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1121));
  INV_X1    g696(.A(G2067), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1043), .A2(new_n1023), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n611), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1117), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1120), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1121), .A2(KEYINPUT60), .A3(new_n1123), .ZN(new_n1127));
  AOI21_X1  g702(.A(KEYINPUT60), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1127), .A2(new_n1128), .A3(new_n611), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT61), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1120), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1130), .B1(new_n1131), .B2(new_n1125), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1121), .A2(KEYINPUT60), .A3(new_n611), .A4(new_n1123), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(new_n1116), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1135), .A2(KEYINPUT61), .A3(new_n1120), .ZN(new_n1136));
  XOR2_X1   g711(.A(KEYINPUT58), .B(G1341), .Z(new_n1137));
  NAND2_X1  g712(.A1(new_n1050), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(G1996), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1023), .A2(new_n1025), .A3(new_n1139), .A4(new_n1026), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n565), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT59), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1141), .B(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1132), .A2(new_n1133), .A3(new_n1136), .A4(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1126), .B1(new_n1129), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g722(.A(KEYINPUT121), .B(new_n1126), .C1(new_n1129), .C2(new_n1144), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1110), .A2(new_n1114), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  AOI211_X1 g724(.A(new_n1047), .B(G286), .C1(new_n1082), .C2(new_n1075), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1039), .A2(new_n1048), .A3(new_n1070), .A4(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT63), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT119), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1151), .A2(KEYINPUT119), .A3(new_n1152), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1035), .A2(G8), .A3(new_n1038), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(new_n1040), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1150), .A2(KEYINPUT63), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1158), .A2(new_n1039), .A3(new_n1159), .A4(new_n1070), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1155), .A2(new_n1156), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(G288), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n1064), .A2(new_n702), .A3(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1054), .B1(new_n1163), .B2(new_n1060), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1070), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1164), .B1(new_n1039), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT62), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1085), .A2(new_n1167), .A3(new_n1087), .ZN(new_n1168));
  AOI21_X1  g743(.A(G301), .B1(new_n1106), .B2(new_n1093), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1167), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1166), .B1(new_n1172), .B2(new_n1071), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1149), .A2(new_n1161), .A3(new_n1173), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n1023), .A2(new_n1076), .ZN(new_n1175));
  XOR2_X1   g750(.A(new_n731), .B(new_n734), .Z(new_n1176));
  XNOR2_X1  g751(.A(new_n813), .B(new_n1122), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n755), .B(new_n1139), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(G1986), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n601), .B(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1175), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1174), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1175), .A2(KEYINPUT46), .A3(new_n1139), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT46), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1175), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1185), .B1(new_n1186), .B2(G1996), .ZN(new_n1187));
  AND2_X1   g762(.A1(new_n1177), .A2(new_n756), .ZN(new_n1188));
  OAI211_X1 g763(.A(new_n1184), .B(new_n1187), .C1(new_n1188), .C2(new_n1186), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n1189), .B(KEYINPUT124), .ZN(new_n1190));
  OR2_X1    g765(.A1(new_n1190), .A2(KEYINPUT47), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(KEYINPUT47), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1177), .A2(new_n1178), .A3(new_n734), .A4(new_n731), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n811), .A2(new_n1122), .A3(new_n812), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1186), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1179), .A2(new_n1175), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1175), .A2(new_n1180), .A3(new_n601), .ZN(new_n1197));
  XNOR2_X1  g772(.A(new_n1197), .B(KEYINPUT48), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1195), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1191), .A2(new_n1192), .A3(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n1200), .B(KEYINPUT125), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1183), .A2(new_n1201), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g777(.A1(G401), .A2(G227), .A3(new_n460), .ZN(new_n1204));
  AND2_X1   g778(.A1(new_n1204), .A2(KEYINPUT126), .ZN(new_n1205));
  NOR2_X1   g779(.A1(new_n1204), .A2(KEYINPUT126), .ZN(new_n1206));
  OAI21_X1  g780(.A(new_n688), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g781(.A(new_n1207), .B1(new_n906), .B2(new_n910), .ZN(new_n1208));
  AND3_X1   g782(.A1(new_n995), .A2(KEYINPUT127), .A3(new_n1208), .ZN(new_n1209));
  AOI21_X1  g783(.A(KEYINPUT127), .B1(new_n995), .B2(new_n1208), .ZN(new_n1210));
  NOR2_X1   g784(.A1(new_n1209), .A2(new_n1210), .ZN(G308));
  NAND2_X1  g785(.A1(new_n995), .A2(new_n1208), .ZN(G225));
endmodule


