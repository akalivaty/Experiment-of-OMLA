

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587;

  XOR2_X1 U322 ( .A(KEYINPUT36), .B(n554), .Z(n495) );
  NOR2_X1 U323 ( .A1(n559), .A2(n493), .ZN(n586) );
  XNOR2_X1 U324 ( .A(n484), .B(n483), .ZN(n575) );
  NOR2_X1 U325 ( .A1(n482), .A2(n545), .ZN(n484) );
  XNOR2_X1 U326 ( .A(n453), .B(n452), .ZN(n517) );
  XOR2_X1 U327 ( .A(n442), .B(n297), .Z(n290) );
  XOR2_X1 U328 ( .A(KEYINPUT112), .B(n460), .Z(n291) );
  XOR2_X1 U329 ( .A(n446), .B(n352), .Z(n292) );
  XNOR2_X1 U330 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U331 ( .A(n438), .B(n437), .ZN(n440) );
  NOR2_X1 U332 ( .A1(n382), .A2(n381), .ZN(n383) );
  XNOR2_X1 U333 ( .A(KEYINPUT119), .B(KEYINPUT54), .ZN(n477) );
  INV_X1 U334 ( .A(G134GAT), .ZN(n315) );
  XNOR2_X1 U335 ( .A(n446), .B(n445), .ZN(n447) );
  INV_X1 U336 ( .A(KEYINPUT96), .ZN(n354) );
  XNOR2_X1 U337 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U338 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U339 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U340 ( .A(n418), .B(n317), .ZN(n318) );
  NOR2_X1 U341 ( .A1(n495), .A2(n410), .ZN(n412) );
  XNOR2_X1 U342 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U343 ( .A(n380), .B(n379), .ZN(n559) );
  XNOR2_X1 U344 ( .A(n451), .B(KEYINPUT105), .ZN(n452) );
  XOR2_X1 U345 ( .A(KEYINPUT81), .B(n566), .Z(n554) );
  XOR2_X1 U346 ( .A(n309), .B(n308), .Z(n538) );
  INV_X1 U347 ( .A(KEYINPUT108), .ZN(n489) );
  XNOR2_X1 U348 ( .A(n496), .B(G218GAT), .ZN(n497) );
  XNOR2_X1 U349 ( .A(n485), .B(G190GAT), .ZN(n486) );
  XNOR2_X1 U350 ( .A(n489), .B(G50GAT), .ZN(n490) );
  XNOR2_X1 U351 ( .A(n454), .B(G43GAT), .ZN(n455) );
  XNOR2_X1 U352 ( .A(n498), .B(n497), .ZN(G1355GAT) );
  XNOR2_X1 U353 ( .A(n487), .B(n486), .ZN(G1351GAT) );
  XNOR2_X1 U354 ( .A(n491), .B(n490), .ZN(G1331GAT) );
  XOR2_X1 U355 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n294) );
  XNOR2_X1 U356 ( .A(KEYINPUT87), .B(KEYINPUT66), .ZN(n293) );
  XNOR2_X1 U357 ( .A(n294), .B(n293), .ZN(n309) );
  XOR2_X1 U358 ( .A(G120GAT), .B(G71GAT), .Z(n442) );
  XOR2_X1 U359 ( .A(KEYINPUT88), .B(G99GAT), .Z(n296) );
  XNOR2_X1 U360 ( .A(G43GAT), .B(G190GAT), .ZN(n295) );
  XNOR2_X1 U361 ( .A(n296), .B(n295), .ZN(n297) );
  NAND2_X1 U362 ( .A1(G227GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U363 ( .A(n290), .B(n298), .ZN(n302) );
  XOR2_X1 U364 ( .A(G176GAT), .B(G15GAT), .Z(n300) );
  XNOR2_X1 U365 ( .A(G169GAT), .B(G113GAT), .ZN(n299) );
  XNOR2_X1 U366 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U367 ( .A(n302), .B(n301), .Z(n307) );
  XOR2_X1 U368 ( .A(G183GAT), .B(KEYINPUT18), .Z(n304) );
  XNOR2_X1 U369 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n303) );
  XNOR2_X1 U370 ( .A(n304), .B(n303), .ZN(n352) );
  XNOR2_X1 U371 ( .A(G134GAT), .B(G127GAT), .ZN(n305) );
  XNOR2_X1 U372 ( .A(n305), .B(KEYINPUT0), .ZN(n388) );
  XNOR2_X1 U373 ( .A(n352), .B(n388), .ZN(n306) );
  XNOR2_X1 U374 ( .A(n307), .B(n306), .ZN(n308) );
  INV_X1 U375 ( .A(n538), .ZN(n545) );
  XOR2_X1 U376 ( .A(KEYINPUT9), .B(KEYINPUT78), .Z(n312) );
  XOR2_X1 U377 ( .A(G50GAT), .B(G162GAT), .Z(n363) );
  XNOR2_X1 U378 ( .A(G99GAT), .B(G106GAT), .ZN(n310) );
  XNOR2_X1 U379 ( .A(n310), .B(G85GAT), .ZN(n438) );
  XNOR2_X1 U380 ( .A(n363), .B(n438), .ZN(n311) );
  XNOR2_X1 U381 ( .A(n312), .B(n311), .ZN(n319) );
  XOR2_X1 U382 ( .A(G29GAT), .B(G43GAT), .Z(n314) );
  XNOR2_X1 U383 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n313) );
  XNOR2_X1 U384 ( .A(n314), .B(n313), .ZN(n418) );
  NAND2_X1 U385 ( .A1(G232GAT), .A2(G233GAT), .ZN(n316) );
  XOR2_X1 U386 ( .A(n319), .B(n318), .Z(n327) );
  XOR2_X1 U387 ( .A(KEYINPUT80), .B(G92GAT), .Z(n321) );
  XNOR2_X1 U388 ( .A(G190GAT), .B(G218GAT), .ZN(n320) );
  XNOR2_X1 U389 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U390 ( .A(G36GAT), .B(n322), .Z(n351) );
  XOR2_X1 U391 ( .A(KEYINPUT79), .B(KEYINPUT10), .Z(n324) );
  XNOR2_X1 U392 ( .A(KEYINPUT67), .B(KEYINPUT11), .ZN(n323) );
  XNOR2_X1 U393 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U394 ( .A(n351), .B(n325), .ZN(n326) );
  XNOR2_X1 U395 ( .A(n327), .B(n326), .ZN(n566) );
  XOR2_X1 U396 ( .A(G78GAT), .B(G211GAT), .Z(n329) );
  XNOR2_X1 U397 ( .A(G183GAT), .B(G127GAT), .ZN(n328) );
  XNOR2_X1 U398 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U399 ( .A(G155GAT), .B(G1GAT), .Z(n331) );
  XNOR2_X1 U400 ( .A(G22GAT), .B(G8GAT), .ZN(n330) );
  XNOR2_X1 U401 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U402 ( .A(n333), .B(n332), .Z(n339) );
  XNOR2_X1 U403 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n334) );
  XNOR2_X1 U404 ( .A(n334), .B(KEYINPUT75), .ZN(n439) );
  XOR2_X1 U405 ( .A(n439), .B(G71GAT), .Z(n336) );
  NAND2_X1 U406 ( .A1(G231GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U407 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U408 ( .A(G15GAT), .B(n337), .ZN(n338) );
  XNOR2_X1 U409 ( .A(n339), .B(n338), .ZN(n347) );
  XOR2_X1 U410 ( .A(KEYINPUT84), .B(KEYINPUT82), .Z(n341) );
  XNOR2_X1 U411 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n340) );
  XNOR2_X1 U412 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U413 ( .A(KEYINPUT83), .B(KEYINPUT85), .Z(n343) );
  XNOR2_X1 U414 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n342) );
  XNOR2_X1 U415 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U416 ( .A(n345), .B(n344), .Z(n346) );
  XOR2_X1 U417 ( .A(n347), .B(n346), .Z(n585) );
  INV_X1 U418 ( .A(n585), .ZN(n499) );
  XOR2_X1 U419 ( .A(KEYINPUT21), .B(G211GAT), .Z(n349) );
  XNOR2_X1 U420 ( .A(KEYINPUT90), .B(G204GAT), .ZN(n348) );
  XNOR2_X1 U421 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U422 ( .A(G197GAT), .B(n350), .Z(n371) );
  XNOR2_X1 U423 ( .A(n371), .B(n351), .ZN(n359) );
  XOR2_X1 U424 ( .A(G176GAT), .B(G64GAT), .Z(n446) );
  NAND2_X1 U425 ( .A1(G226GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U426 ( .A(n292), .B(n353), .ZN(n357) );
  XOR2_X1 U427 ( .A(G169GAT), .B(G8GAT), .Z(n421) );
  XNOR2_X1 U428 ( .A(n421), .B(KEYINPUT95), .ZN(n355) );
  XOR2_X1 U429 ( .A(n359), .B(n358), .Z(n360) );
  INV_X1 U430 ( .A(n360), .ZN(n535) );
  NAND2_X1 U431 ( .A1(n535), .A2(n538), .ZN(n376) );
  XOR2_X1 U432 ( .A(KEYINPUT91), .B(KEYINPUT23), .Z(n362) );
  XNOR2_X1 U433 ( .A(KEYINPUT22), .B(KEYINPUT24), .ZN(n361) );
  XNOR2_X1 U434 ( .A(n362), .B(n361), .ZN(n375) );
  XOR2_X1 U435 ( .A(G106GAT), .B(G218GAT), .Z(n365) );
  XOR2_X1 U436 ( .A(G148GAT), .B(G78GAT), .Z(n441) );
  XNOR2_X1 U437 ( .A(n363), .B(n441), .ZN(n364) );
  XNOR2_X1 U438 ( .A(n365), .B(n364), .ZN(n370) );
  XNOR2_X1 U439 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n366) );
  XNOR2_X1 U440 ( .A(n366), .B(KEYINPUT2), .ZN(n384) );
  XOR2_X1 U441 ( .A(KEYINPUT89), .B(n384), .Z(n368) );
  NAND2_X1 U442 ( .A1(G228GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U443 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U444 ( .A(n370), .B(n369), .Z(n373) );
  XOR2_X1 U445 ( .A(G141GAT), .B(G22GAT), .Z(n417) );
  XNOR2_X1 U446 ( .A(n417), .B(n371), .ZN(n372) );
  XNOR2_X1 U447 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U448 ( .A(n375), .B(n374), .ZN(n457) );
  NAND2_X1 U449 ( .A1(n376), .A2(n457), .ZN(n377) );
  XNOR2_X1 U450 ( .A(n377), .B(KEYINPUT25), .ZN(n378) );
  XNOR2_X1 U451 ( .A(n378), .B(KEYINPUT98), .ZN(n382) );
  XNOR2_X1 U452 ( .A(n360), .B(KEYINPUT27), .ZN(n404) );
  NOR2_X1 U453 ( .A1(n538), .A2(n457), .ZN(n380) );
  XNOR2_X1 U454 ( .A(KEYINPUT26), .B(KEYINPUT97), .ZN(n379) );
  NOR2_X1 U455 ( .A1(n404), .A2(n559), .ZN(n381) );
  XNOR2_X1 U456 ( .A(n383), .B(KEYINPUT99), .ZN(n403) );
  XOR2_X1 U457 ( .A(G113GAT), .B(G1GAT), .Z(n415) );
  XOR2_X1 U458 ( .A(n384), .B(n415), .Z(n386) );
  NAND2_X1 U459 ( .A1(G225GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U460 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U461 ( .A(n387), .B(KEYINPUT92), .Z(n390) );
  XNOR2_X1 U462 ( .A(n388), .B(KEYINPUT94), .ZN(n389) );
  XNOR2_X1 U463 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U464 ( .A(G85GAT), .B(G162GAT), .Z(n392) );
  XNOR2_X1 U465 ( .A(G29GAT), .B(G120GAT), .ZN(n391) );
  XNOR2_X1 U466 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U467 ( .A(n394), .B(n393), .Z(n402) );
  XOR2_X1 U468 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n396) );
  XNOR2_X1 U469 ( .A(KEYINPUT6), .B(KEYINPUT93), .ZN(n395) );
  XNOR2_X1 U470 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U471 ( .A(KEYINPUT1), .B(G57GAT), .Z(n398) );
  XNOR2_X1 U472 ( .A(G141GAT), .B(G148GAT), .ZN(n397) );
  XNOR2_X1 U473 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U474 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U475 ( .A(n402), .B(n401), .Z(n514) );
  NAND2_X1 U476 ( .A1(n403), .A2(n514), .ZN(n408) );
  NOR2_X1 U477 ( .A1(n404), .A2(n514), .ZN(n544) );
  XOR2_X1 U478 ( .A(KEYINPUT28), .B(KEYINPUT68), .Z(n405) );
  XOR2_X1 U479 ( .A(n457), .B(n405), .Z(n488) );
  INV_X1 U480 ( .A(n488), .ZN(n548) );
  NOR2_X1 U481 ( .A1(n538), .A2(n548), .ZN(n406) );
  NAND2_X1 U482 ( .A1(n544), .A2(n406), .ZN(n407) );
  NAND2_X1 U483 ( .A1(n408), .A2(n407), .ZN(n501) );
  NAND2_X1 U484 ( .A1(n499), .A2(n501), .ZN(n409) );
  XOR2_X1 U485 ( .A(KEYINPUT103), .B(n409), .Z(n410) );
  XNOR2_X1 U486 ( .A(KEYINPUT37), .B(KEYINPUT104), .ZN(n411) );
  XNOR2_X1 U487 ( .A(n412), .B(n411), .ZN(n532) );
  XOR2_X1 U488 ( .A(G197GAT), .B(G15GAT), .Z(n414) );
  XNOR2_X1 U489 ( .A(G50GAT), .B(G36GAT), .ZN(n413) );
  XNOR2_X1 U490 ( .A(n414), .B(n413), .ZN(n416) );
  XOR2_X1 U491 ( .A(n416), .B(n415), .Z(n424) );
  XOR2_X1 U492 ( .A(n418), .B(n417), .Z(n420) );
  NAND2_X1 U493 ( .A1(G229GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U494 ( .A(n420), .B(n419), .ZN(n422) );
  XNOR2_X1 U495 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U496 ( .A(n424), .B(n423), .ZN(n432) );
  XOR2_X1 U497 ( .A(KEYINPUT72), .B(KEYINPUT74), .Z(n426) );
  XNOR2_X1 U498 ( .A(KEYINPUT73), .B(KEYINPUT71), .ZN(n425) );
  XNOR2_X1 U499 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U500 ( .A(KEYINPUT29), .B(KEYINPUT70), .Z(n428) );
  XNOR2_X1 U501 ( .A(KEYINPUT30), .B(KEYINPUT69), .ZN(n427) );
  XNOR2_X1 U502 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U503 ( .A(n430), .B(n429), .Z(n431) );
  XOR2_X1 U504 ( .A(n432), .B(n431), .Z(n520) );
  INV_X1 U505 ( .A(n520), .ZN(n578) );
  XOR2_X1 U506 ( .A(KEYINPUT77), .B(KEYINPUT32), .Z(n434) );
  XNOR2_X1 U507 ( .A(KEYINPUT33), .B(KEYINPUT76), .ZN(n433) );
  XOR2_X1 U508 ( .A(n434), .B(n433), .Z(n450) );
  NAND2_X1 U509 ( .A1(G230GAT), .A2(G233GAT), .ZN(n436) );
  INV_X1 U510 ( .A(KEYINPUT31), .ZN(n435) );
  XNOR2_X1 U511 ( .A(n440), .B(n439), .ZN(n444) );
  XNOR2_X1 U512 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U513 ( .A(n444), .B(n443), .ZN(n448) );
  XNOR2_X1 U514 ( .A(G204GAT), .B(G92GAT), .ZN(n445) );
  XNOR2_X1 U515 ( .A(n450), .B(n449), .ZN(n459) );
  INV_X1 U516 ( .A(n459), .ZN(n468) );
  NAND2_X1 U517 ( .A1(n578), .A2(n468), .ZN(n503) );
  NOR2_X1 U518 ( .A1(n532), .A2(n503), .ZN(n453) );
  XNOR2_X1 U519 ( .A(KEYINPUT106), .B(KEYINPUT38), .ZN(n451) );
  NOR2_X1 U520 ( .A1(n545), .A2(n517), .ZN(n456) );
  XNOR2_X1 U521 ( .A(KEYINPUT40), .B(KEYINPUT107), .ZN(n454) );
  XNOR2_X1 U522 ( .A(n456), .B(n455), .ZN(G1330GAT) );
  AND2_X1 U523 ( .A1(n514), .A2(n457), .ZN(n479) );
  XOR2_X1 U524 ( .A(KEYINPUT118), .B(n360), .Z(n476) );
  XNOR2_X1 U525 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n475) );
  INV_X1 U526 ( .A(KEYINPUT114), .ZN(n464) );
  XNOR2_X1 U527 ( .A(KEYINPUT41), .B(KEYINPUT65), .ZN(n458) );
  XNOR2_X1 U528 ( .A(n459), .B(n458), .ZN(n519) );
  NAND2_X1 U529 ( .A1(n519), .A2(n578), .ZN(n461) );
  XOR2_X1 U530 ( .A(KEYINPUT113), .B(KEYINPUT46), .Z(n460) );
  XNOR2_X1 U531 ( .A(n461), .B(n291), .ZN(n462) );
  NOR2_X1 U532 ( .A1(n585), .A2(n462), .ZN(n463) );
  XNOR2_X1 U533 ( .A(n464), .B(n463), .ZN(n465) );
  NOR2_X1 U534 ( .A1(n465), .A2(n566), .ZN(n466) );
  XNOR2_X1 U535 ( .A(n466), .B(KEYINPUT47), .ZN(n473) );
  NOR2_X1 U536 ( .A1(n495), .A2(n499), .ZN(n467) );
  XNOR2_X1 U537 ( .A(n467), .B(KEYINPUT45), .ZN(n469) );
  NAND2_X1 U538 ( .A1(n469), .A2(n468), .ZN(n470) );
  NOR2_X1 U539 ( .A1(n578), .A2(n470), .ZN(n471) );
  XNOR2_X1 U540 ( .A(KEYINPUT115), .B(n471), .ZN(n472) );
  NAND2_X1 U541 ( .A1(n473), .A2(n472), .ZN(n474) );
  XNOR2_X1 U542 ( .A(n475), .B(n474), .ZN(n543) );
  NAND2_X1 U543 ( .A1(n476), .A2(n543), .ZN(n478) );
  XNOR2_X1 U544 ( .A(n478), .B(n477), .ZN(n492) );
  NAND2_X1 U545 ( .A1(n479), .A2(n492), .ZN(n481) );
  XOR2_X1 U546 ( .A(KEYINPUT120), .B(KEYINPUT55), .Z(n480) );
  XNOR2_X1 U547 ( .A(n481), .B(n480), .ZN(n482) );
  INV_X1 U548 ( .A(KEYINPUT121), .ZN(n483) );
  NAND2_X1 U549 ( .A1(n575), .A2(n554), .ZN(n487) );
  XOR2_X1 U550 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n485) );
  NOR2_X1 U551 ( .A1(n488), .A2(n517), .ZN(n491) );
  NAND2_X1 U552 ( .A1(n514), .A2(n492), .ZN(n493) );
  INV_X1 U553 ( .A(n586), .ZN(n494) );
  NOR2_X1 U554 ( .A1(n495), .A2(n494), .ZN(n498) );
  XNOR2_X1 U555 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n496) );
  NOR2_X1 U556 ( .A1(n554), .A2(n499), .ZN(n500) );
  XNOR2_X1 U557 ( .A(n500), .B(KEYINPUT16), .ZN(n502) );
  NAND2_X1 U558 ( .A1(n502), .A2(n501), .ZN(n521) );
  NOR2_X1 U559 ( .A1(n503), .A2(n521), .ZN(n511) );
  INV_X1 U560 ( .A(n514), .ZN(n533) );
  NAND2_X1 U561 ( .A1(n511), .A2(n533), .ZN(n504) );
  XNOR2_X1 U562 ( .A(n504), .B(KEYINPUT34), .ZN(n505) );
  XNOR2_X1 U563 ( .A(G1GAT), .B(n505), .ZN(G1324GAT) );
  NAND2_X1 U564 ( .A1(n511), .A2(n535), .ZN(n506) );
  XNOR2_X1 U565 ( .A(n506), .B(KEYINPUT100), .ZN(n507) );
  XNOR2_X1 U566 ( .A(G8GAT), .B(n507), .ZN(G1325GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n509) );
  NAND2_X1 U568 ( .A1(n511), .A2(n538), .ZN(n508) );
  XNOR2_X1 U569 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U570 ( .A(G15GAT), .B(n510), .Z(G1326GAT) );
  NAND2_X1 U571 ( .A1(n511), .A2(n548), .ZN(n512) );
  XNOR2_X1 U572 ( .A(n512), .B(KEYINPUT102), .ZN(n513) );
  XNOR2_X1 U573 ( .A(G22GAT), .B(n513), .ZN(G1327GAT) );
  NOR2_X1 U574 ( .A1(n514), .A2(n517), .ZN(n516) );
  XNOR2_X1 U575 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n515) );
  XNOR2_X1 U576 ( .A(n516), .B(n515), .ZN(G1328GAT) );
  NOR2_X1 U577 ( .A1(n360), .A2(n517), .ZN(n518) );
  XOR2_X1 U578 ( .A(G36GAT), .B(n518), .Z(G1329GAT) );
  XNOR2_X1 U579 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n523) );
  NAND2_X1 U580 ( .A1(n520), .A2(n519), .ZN(n531) );
  NOR2_X1 U581 ( .A1(n531), .A2(n521), .ZN(n528) );
  NAND2_X1 U582 ( .A1(n533), .A2(n528), .ZN(n522) );
  XNOR2_X1 U583 ( .A(n523), .B(n522), .ZN(G1332GAT) );
  XOR2_X1 U584 ( .A(G64GAT), .B(KEYINPUT109), .Z(n525) );
  NAND2_X1 U585 ( .A1(n528), .A2(n535), .ZN(n524) );
  XNOR2_X1 U586 ( .A(n525), .B(n524), .ZN(G1333GAT) );
  NAND2_X1 U587 ( .A1(n528), .A2(n538), .ZN(n526) );
  XNOR2_X1 U588 ( .A(n526), .B(KEYINPUT110), .ZN(n527) );
  XNOR2_X1 U589 ( .A(G71GAT), .B(n527), .ZN(G1334GAT) );
  XOR2_X1 U590 ( .A(G78GAT), .B(KEYINPUT43), .Z(n530) );
  NAND2_X1 U591 ( .A1(n528), .A2(n548), .ZN(n529) );
  XNOR2_X1 U592 ( .A(n530), .B(n529), .ZN(G1335GAT) );
  NOR2_X1 U593 ( .A1(n532), .A2(n531), .ZN(n540) );
  NAND2_X1 U594 ( .A1(n533), .A2(n540), .ZN(n534) );
  XNOR2_X1 U595 ( .A(G85GAT), .B(n534), .ZN(G1336GAT) );
  XOR2_X1 U596 ( .A(G92GAT), .B(KEYINPUT111), .Z(n537) );
  NAND2_X1 U597 ( .A1(n540), .A2(n535), .ZN(n536) );
  XNOR2_X1 U598 ( .A(n537), .B(n536), .ZN(G1337GAT) );
  NAND2_X1 U599 ( .A1(n540), .A2(n538), .ZN(n539) );
  XNOR2_X1 U600 ( .A(n539), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U601 ( .A1(n540), .A2(n548), .ZN(n541) );
  XNOR2_X1 U602 ( .A(n541), .B(KEYINPUT44), .ZN(n542) );
  XNOR2_X1 U603 ( .A(G106GAT), .B(n542), .ZN(G1339GAT) );
  NAND2_X1 U604 ( .A1(n544), .A2(n543), .ZN(n558) );
  NOR2_X1 U605 ( .A1(n545), .A2(n558), .ZN(n546) );
  XOR2_X1 U606 ( .A(KEYINPUT116), .B(n546), .Z(n547) );
  NOR2_X1 U607 ( .A1(n548), .A2(n547), .ZN(n555) );
  NAND2_X1 U608 ( .A1(n578), .A2(n555), .ZN(n549) );
  XNOR2_X1 U609 ( .A(n549), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U610 ( .A(G120GAT), .B(KEYINPUT49), .Z(n551) );
  NAND2_X1 U611 ( .A1(n555), .A2(n519), .ZN(n550) );
  XNOR2_X1 U612 ( .A(n551), .B(n550), .ZN(G1341GAT) );
  NAND2_X1 U613 ( .A1(n555), .A2(n585), .ZN(n552) );
  XNOR2_X1 U614 ( .A(n552), .B(KEYINPUT50), .ZN(n553) );
  XNOR2_X1 U615 ( .A(G127GAT), .B(n553), .ZN(G1342GAT) );
  XOR2_X1 U616 ( .A(G134GAT), .B(KEYINPUT51), .Z(n557) );
  NAND2_X1 U617 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U618 ( .A(n557), .B(n556), .ZN(G1343GAT) );
  NOR2_X1 U619 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U620 ( .A(KEYINPUT117), .B(n560), .Z(n567) );
  NAND2_X1 U621 ( .A1(n567), .A2(n578), .ZN(n561) );
  XNOR2_X1 U622 ( .A(G141GAT), .B(n561), .ZN(G1344GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n563) );
  NAND2_X1 U624 ( .A1(n567), .A2(n519), .ZN(n562) );
  XNOR2_X1 U625 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(n564), .ZN(G1345GAT) );
  NAND2_X1 U627 ( .A1(n567), .A2(n585), .ZN(n565) );
  XNOR2_X1 U628 ( .A(n565), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U629 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U630 ( .A(n568), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U631 ( .A1(n578), .A2(n575), .ZN(n569) );
  XNOR2_X1 U632 ( .A(n569), .B(KEYINPUT122), .ZN(n570) );
  XNOR2_X1 U633 ( .A(n570), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U634 ( .A1(n575), .A2(n519), .ZN(n572) );
  XOR2_X1 U635 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n571) );
  XNOR2_X1 U636 ( .A(n572), .B(n571), .ZN(n574) );
  XOR2_X1 U637 ( .A(G176GAT), .B(KEYINPUT56), .Z(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(G1349GAT) );
  NAND2_X1 U639 ( .A1(n575), .A2(n585), .ZN(n576) );
  XNOR2_X1 U640 ( .A(n576), .B(KEYINPUT124), .ZN(n577) );
  XNOR2_X1 U641 ( .A(n577), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n580) );
  NAND2_X1 U643 ( .A1(n586), .A2(n578), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n583) );
  NAND2_X1 U647 ( .A1(n586), .A2(n459), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(G204GAT), .B(n584), .ZN(G1353GAT) );
  NAND2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U651 ( .A(n587), .B(G211GAT), .ZN(G1354GAT) );
endmodule

