//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 0 1 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 1 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925;
  INV_X1    g000(.A(KEYINPUT90), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G43gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G71gat), .B(G99gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G127gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT70), .B1(new_n207), .B2(G134gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(G113gat), .B(G120gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n208), .B1(new_n209), .B2(KEYINPUT1), .ZN(new_n210));
  XNOR2_X1  g009(.A(G127gat), .B(G134gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n213), .B(KEYINPUT24), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n214), .B1(G183gat), .B2(G190gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT23), .ZN(new_n217));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(G169gat), .B2(G176gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n217), .A2(new_n218), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT65), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n217), .A2(KEYINPUT65), .A3(new_n220), .A4(new_n218), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n215), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n225), .A2(KEYINPUT66), .A3(new_n226), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT67), .B1(G183gat), .B2(G190gat), .ZN(new_n231));
  OR3_X1    g030(.A1(KEYINPUT67), .A2(G183gat), .A3(G190gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n214), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n221), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(KEYINPUT25), .A3(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n229), .A2(new_n230), .A3(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(KEYINPUT27), .B(G183gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n238), .A2(G190gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  OR2_X1    g039(.A1(new_n240), .A2(KEYINPUT69), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(KEYINPUT69), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n216), .A2(KEYINPUT26), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT26), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n218), .A2(new_n247), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n246), .B(new_n213), .C1(new_n248), .C2(new_n216), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n241), .A2(KEYINPUT68), .A3(KEYINPUT28), .A4(new_n242), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n245), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n212), .B1(new_n236), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G227gat), .ZN(new_n255));
  INV_X1    g054(.A(G233gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n236), .A2(new_n212), .A3(new_n252), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n254), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT33), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n206), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n258), .ZN(new_n262));
  OAI22_X1  g061(.A1(new_n262), .A2(new_n253), .B1(new_n255), .B2(new_n256), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT34), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT71), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n259), .A2(KEYINPUT32), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(new_n270), .A3(KEYINPUT34), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n259), .B(KEYINPUT32), .C1(KEYINPUT71), .C2(new_n264), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n261), .A2(new_n266), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n268), .A2(new_n271), .A3(new_n272), .A4(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n271), .A2(new_n272), .ZN(new_n275));
  INV_X1    g074(.A(new_n273), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n275), .B1(new_n276), .B2(new_n267), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT36), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT29), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n225), .A2(KEYINPUT66), .A3(new_n226), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT66), .B1(new_n225), .B2(new_n226), .ZN(new_n282));
  INV_X1    g081(.A(new_n235), .ZN(new_n283));
  NOR3_X1   g082(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n252), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n280), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(G226gat), .A2(G233gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(KEYINPUT74), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n287), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n290), .B1(new_n284), .B2(new_n285), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT75), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n236), .A2(new_n252), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n294), .A2(KEYINPUT75), .A3(new_n290), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n289), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT76), .ZN(new_n297));
  XNOR2_X1  g096(.A(G211gat), .B(G218gat), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n298), .A2(KEYINPUT73), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(KEYINPUT73), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT22), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT72), .B(G211gat), .ZN(new_n303));
  INV_X1    g102(.A(G218gat), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G197gat), .B(G204gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n301), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n306), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n308), .A2(new_n300), .A3(new_n299), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n296), .A2(new_n297), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(KEYINPUT75), .B1(new_n294), .B2(new_n290), .ZN(new_n313));
  AOI211_X1 g112(.A(new_n292), .B(new_n287), .C1(new_n236), .C2(new_n252), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n310), .B1(new_n315), .B2(new_n289), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n286), .A2(new_n287), .ZN(new_n317));
  INV_X1    g116(.A(new_n288), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n294), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n317), .A2(new_n310), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT76), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n312), .B1(new_n316), .B2(new_n321), .ZN(new_n322));
  XOR2_X1   g121(.A(KEYINPUT77), .B(G64gat), .Z(new_n323));
  XNOR2_X1  g122(.A(KEYINPUT78), .B(G92gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n323), .B(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G8gat), .B(G36gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n325), .B(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n322), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT30), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT85), .ZN(new_n331));
  XOR2_X1   g130(.A(G141gat), .B(G148gat), .Z(new_n332));
  INV_X1    g131(.A(G155gat), .ZN(new_n333));
  INV_X1    g132(.A(G162gat), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT2), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G155gat), .B(G162gat), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n332), .A2(new_n337), .A3(new_n335), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n339), .A2(KEYINPUT79), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT79), .B1(new_n339), .B2(new_n340), .ZN(new_n343));
  OAI211_X1 g142(.A(KEYINPUT80), .B(KEYINPUT3), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT3), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n339), .A2(new_n340), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT79), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n345), .B1(new_n348), .B2(new_n341), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n346), .A2(KEYINPUT3), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT80), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n212), .B(new_n344), .C1(new_n349), .C2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(G225gat), .A2(G233gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(KEYINPUT81), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n212), .A2(new_n346), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT4), .ZN(new_n358));
  INV_X1    g157(.A(new_n357), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT82), .B(KEYINPUT4), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n353), .A2(new_n356), .A3(new_n358), .A4(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n212), .B1(new_n342), .B2(new_n343), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(new_n359), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n355), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n362), .A2(KEYINPUT5), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n359), .A2(KEYINPUT84), .A3(KEYINPUT4), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT84), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT4), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n368), .B1(new_n357), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n357), .A2(new_n360), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n367), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n355), .A2(KEYINPUT5), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n372), .A2(new_n353), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n366), .A2(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(KEYINPUT83), .B(KEYINPUT0), .Z(new_n376));
  XNOR2_X1  g175(.A(G1gat), .B(G29gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G57gat), .B(G85gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT6), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n331), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n366), .A2(new_n374), .A3(new_n380), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n382), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n375), .A2(KEYINPUT85), .A3(KEYINPUT6), .A4(new_n381), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n384), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  OR2_X1    g187(.A1(new_n316), .A2(new_n321), .ZN(new_n389));
  INV_X1    g188(.A(new_n327), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(new_n312), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n322), .A2(KEYINPUT30), .A3(new_n327), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n330), .A2(new_n388), .A3(new_n391), .A4(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT86), .ZN(new_n394));
  AND3_X1   g193(.A1(new_n322), .A2(KEYINPUT30), .A3(new_n327), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT30), .B1(new_n322), .B2(new_n327), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT86), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n397), .A2(new_n398), .A3(new_n388), .A4(new_n391), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n394), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT88), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT87), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n307), .A2(new_n309), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n301), .A2(KEYINPUT87), .A3(new_n305), .A4(new_n306), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n280), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n401), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n403), .A2(KEYINPUT88), .A3(new_n280), .A4(new_n405), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n407), .A2(new_n345), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n346), .ZN(new_n410));
  NAND2_X1  g209(.A1(G228gat), .A2(G233gat), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n311), .B1(KEYINPUT29), .B2(new_n350), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n345), .B1(new_n311), .B2(KEYINPUT29), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n414), .B1(new_n342), .B2(new_n343), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n411), .B1(new_n415), .B2(new_n412), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(G22gat), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n413), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n418), .B1(new_n413), .B2(new_n417), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT89), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n421), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT89), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n423), .A2(new_n419), .A3(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(G78gat), .B(G106gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT31), .B(G50gat), .ZN(new_n427));
  XOR2_X1   g226(.A(new_n426), .B(new_n427), .Z(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n422), .A2(new_n425), .A3(new_n429), .ZN(new_n430));
  OAI211_X1 g229(.A(KEYINPUT89), .B(new_n428), .C1(new_n420), .C2(new_n421), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n202), .B(new_n279), .C1(new_n400), .C2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n433), .B1(new_n394), .B2(new_n399), .ZN(new_n435));
  XOR2_X1   g234(.A(new_n278), .B(KEYINPUT36), .Z(new_n436));
  OAI21_X1  g235(.A(KEYINPUT90), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT37), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n322), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n296), .A2(new_n310), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n317), .A2(new_n319), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n440), .B(KEYINPUT37), .C1(new_n310), .C2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT38), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n439), .A2(new_n442), .A3(new_n443), .A4(new_n390), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n328), .A2(new_n387), .A3(new_n384), .A4(new_n386), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT91), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n389), .A2(KEYINPUT37), .A3(new_n312), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n448), .A2(new_n390), .A3(new_n439), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT38), .ZN(new_n450));
  INV_X1    g249(.A(new_n388), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT91), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n451), .A2(new_n444), .A3(new_n452), .A4(new_n328), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n447), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n397), .A2(new_n391), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n356), .B1(new_n372), .B2(new_n353), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT39), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n381), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n364), .A2(new_n355), .ZN(new_n459));
  OR2_X1    g258(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n458), .B1(new_n460), .B2(new_n457), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n461), .B(KEYINPUT40), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n455), .A2(new_n382), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n454), .A2(new_n433), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n434), .A2(new_n437), .A3(new_n464), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n394), .A2(new_n399), .A3(KEYINPUT35), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n278), .A2(new_n430), .A3(new_n431), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n393), .A2(KEYINPUT92), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT92), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n397), .A2(new_n469), .A3(new_n388), .A4(new_n391), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n470), .A3(new_n467), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT35), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n466), .A2(new_n467), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n465), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT101), .ZN(new_n475));
  AND2_X1   g274(.A1(G15gat), .A2(G22gat), .ZN(new_n476));
  NOR2_X1   g275(.A1(G15gat), .A2(G22gat), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT100), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(G15gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n418), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT100), .ZN(new_n481));
  NAND2_X1  g280(.A1(G15gat), .A2(G22gat), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(G1gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT16), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(G8gat), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n478), .A2(new_n483), .A3(new_n485), .ZN(new_n489));
  AND4_X1   g288(.A1(new_n475), .A2(new_n487), .A3(new_n488), .A4(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT101), .B1(new_n484), .B2(new_n486), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n488), .B1(new_n491), .B2(new_n489), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT102), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT17), .ZN(new_n495));
  INV_X1    g294(.A(G50gat), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n496), .A2(G43gat), .ZN(new_n497));
  INV_X1    g296(.A(G43gat), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n498), .A2(G50gat), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT94), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(G50gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n496), .A2(G43gat), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT94), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n500), .A2(KEYINPUT15), .A3(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(G29gat), .A2(G36gat), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT95), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT14), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(KEYINPUT95), .A2(KEYINPUT14), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n506), .A2(new_n510), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT99), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(G29gat), .A2(G36gat), .ZN(new_n514));
  AND3_X1   g313(.A1(new_n505), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  OR3_X1    g314(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT99), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT15), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n501), .A2(KEYINPUT97), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT97), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n519), .A2(new_n498), .A3(G50gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n498), .A2(KEYINPUT96), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT96), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(G43gat), .ZN(new_n524));
  AND3_X1   g323(.A1(new_n522), .A2(new_n524), .A3(new_n496), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n517), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT98), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI211_X1 g327(.A(KEYINPUT98), .B(new_n517), .C1(new_n521), .C2(new_n525), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n515), .A2(new_n516), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n514), .B1(new_n511), .B2(new_n512), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n531), .A2(KEYINPUT15), .A3(new_n504), .A4(new_n500), .ZN(new_n532));
  AOI211_X1 g331(.A(new_n494), .B(new_n495), .C1(new_n530), .C2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n494), .A2(new_n495), .ZN(new_n534));
  NAND2_X1  g333(.A1(KEYINPUT102), .A2(KEYINPUT17), .ZN(new_n535));
  AND4_X1   g334(.A1(new_n532), .A2(new_n530), .A3(new_n534), .A4(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n493), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(G229gat), .A2(G233gat), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n493), .B1(new_n532), .B2(new_n530), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n537), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT18), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n537), .A2(KEYINPUT18), .A3(new_n538), .A4(new_n540), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n538), .B(KEYINPUT13), .Z(new_n545));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n532), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n487), .A2(new_n475), .A3(new_n489), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(G8gat), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n545), .B1(new_n549), .B2(new_n539), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT103), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n546), .B(new_n548), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n553), .A2(KEYINPUT103), .A3(new_n545), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n543), .A2(new_n544), .A3(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(G169gat), .B(G197gat), .Z(new_n557));
  XNOR2_X1  g356(.A(G113gat), .B(G141gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XOR2_X1   g358(.A(KEYINPUT93), .B(KEYINPUT11), .Z(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT12), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n556), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n543), .A2(new_n555), .A3(new_n544), .A4(new_n562), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n568));
  XOR2_X1   g367(.A(G57gat), .B(G64gat), .Z(new_n569));
  NAND2_X1  g368(.A1(G71gat), .A2(G78gat), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT9), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G71gat), .B(G78gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n548), .B1(KEYINPUT21), .B2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(G183gat), .ZN(new_n577));
  INV_X1    g376(.A(G231gat), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n578), .A2(new_n256), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n577), .A2(new_n579), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n568), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n582), .ZN(new_n584));
  INV_X1    g383(.A(new_n568), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n584), .A2(new_n580), .A3(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n575), .A2(KEYINPUT21), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(G211gat), .ZN(new_n588));
  XOR2_X1   g387(.A(G127gat), .B(G155gat), .Z(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  AND3_X1   g391(.A1(new_n583), .A2(new_n586), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n592), .B1(new_n583), .B2(new_n586), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT8), .ZN(new_n597));
  INV_X1    g396(.A(G85gat), .ZN(new_n598));
  INV_X1    g397(.A(G92gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AND3_X1   g399(.A1(new_n597), .A2(KEYINPUT106), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(KEYINPUT106), .B1(new_n597), .B2(new_n600), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT107), .ZN(new_n604));
  XOR2_X1   g403(.A(G99gat), .B(G106gat), .Z(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(G85gat), .A2(G92gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT7), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n603), .A2(new_n604), .A3(new_n606), .A4(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n608), .B1(new_n601), .B2(new_n602), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(new_n605), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n606), .B(new_n608), .C1(new_n601), .C2(new_n602), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(KEYINPUT107), .A3(new_n612), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n609), .B(new_n613), .C1(new_n533), .C2(new_n536), .ZN(new_n614));
  XNOR2_X1  g413(.A(G190gat), .B(G218gat), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n615), .B(KEYINPUT108), .Z(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(new_n609), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n546), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n614), .A2(new_n616), .A3(new_n618), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(KEYINPUT109), .ZN(new_n621));
  XNOR2_X1  g420(.A(G134gat), .B(G162gat), .ZN(new_n622));
  AOI21_X1  g421(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n614), .A2(new_n618), .A3(new_n619), .ZN(new_n626));
  INV_X1    g425(.A(new_n616), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n620), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n625), .A2(new_n629), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(G230gat), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n635), .A2(new_n256), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n573), .B(new_n574), .Z(new_n637));
  NAND3_X1  g436(.A1(new_n613), .A2(new_n609), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT110), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n613), .A2(new_n637), .A3(KEYINPUT110), .A4(new_n609), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT10), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n575), .A2(new_n612), .A3(new_n611), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n617), .A2(KEYINPUT10), .A3(new_n575), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n636), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AOI211_X1 g446(.A(new_n635), .B(new_n256), .C1(new_n642), .C2(new_n644), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(G120gat), .B(G148gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(G176gat), .B(G204gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n649), .B(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n595), .A2(new_n634), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n474), .A2(new_n567), .A3(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n658), .A2(new_n388), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(new_n485), .ZN(G1324gat));
  INV_X1    g459(.A(new_n455), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(KEYINPUT112), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT112), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n664), .B1(new_n658), .B2(new_n661), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(G8gat), .ZN(new_n667));
  XOR2_X1   g466(.A(KEYINPUT16), .B(G8gat), .Z(new_n668));
  NAND3_X1  g467(.A1(new_n662), .A2(KEYINPUT42), .A3(new_n668), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n663), .A2(new_n665), .A3(new_n668), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT111), .B(KEYINPUT42), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n667), .B(new_n669), .C1(new_n670), .C2(new_n671), .ZN(G1325gat));
  NOR3_X1   g471(.A1(new_n658), .A2(new_n479), .A3(new_n279), .ZN(new_n673));
  INV_X1    g472(.A(new_n658), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(new_n278), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n673), .B1(new_n479), .B2(new_n675), .ZN(G1326gat));
  NOR2_X1   g475(.A1(new_n658), .A2(new_n433), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT43), .B(G22gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  NOR3_X1   g478(.A1(new_n595), .A2(new_n566), .A3(new_n654), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n474), .A2(new_n633), .A3(new_n680), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n681), .A2(G29gat), .A3(new_n388), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(KEYINPUT45), .Z(new_n683));
  NAND3_X1  g482(.A1(new_n474), .A2(KEYINPUT44), .A3(new_n633), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n471), .A2(new_n472), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n394), .A2(new_n399), .A3(new_n467), .A4(KEYINPUT35), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n435), .A2(new_n436), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n688), .B1(new_n689), .B2(new_n464), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n685), .B1(new_n690), .B2(new_n634), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n684), .A2(new_n691), .A3(new_n680), .ZN(new_n692));
  OAI21_X1  g491(.A(G29gat), .B1(new_n692), .B2(new_n388), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n683), .A2(new_n693), .ZN(G1328gat));
  NOR3_X1   g493(.A1(new_n681), .A2(G36gat), .A3(new_n661), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT46), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n696), .ZN(new_n698));
  OAI21_X1  g497(.A(G36gat), .B1(new_n692), .B2(new_n661), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(G1329gat));
  NAND2_X1  g499(.A1(new_n522), .A2(new_n524), .ZN(new_n701));
  INV_X1    g500(.A(new_n278), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n701), .B1(new_n681), .B2(new_n702), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n279), .A2(new_n701), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n703), .B1(new_n692), .B2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g505(.A1(new_n684), .A2(new_n691), .A3(new_n432), .A4(new_n680), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(G50gat), .ZN(new_n708));
  AOI21_X1  g507(.A(KEYINPUT48), .B1(new_n708), .B2(KEYINPUT113), .ZN(new_n709));
  OR3_X1    g508(.A1(new_n681), .A2(G50gat), .A3(new_n433), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n708), .B(new_n710), .C1(KEYINPUT113), .C2(KEYINPUT48), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(G1331gat));
  NAND2_X1  g513(.A1(new_n689), .A2(new_n464), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n473), .ZN(new_n716));
  INV_X1    g515(.A(new_n595), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n717), .A2(new_n633), .A3(new_n655), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n716), .A2(new_n566), .A3(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n719), .A2(new_n388), .ZN(new_n720));
  XOR2_X1   g519(.A(KEYINPUT114), .B(G57gat), .Z(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1332gat));
  NOR2_X1   g521(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n661), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n724));
  XOR2_X1   g523(.A(new_n724), .B(KEYINPUT115), .Z(new_n725));
  OR3_X1    g524(.A1(new_n719), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n723), .B1(new_n719), .B2(new_n725), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(KEYINPUT116), .B(KEYINPUT117), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1333gat));
  OR3_X1    g529(.A1(new_n719), .A2(G71gat), .A3(new_n702), .ZN(new_n731));
  OAI21_X1  g530(.A(G71gat), .B1(new_n719), .B2(new_n279), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n733), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n433), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g535(.A1(new_n595), .A2(new_n567), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n684), .A2(new_n691), .A3(new_n654), .A4(new_n737), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n738), .A2(new_n598), .A3(new_n388), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT51), .ZN(new_n740));
  AND4_X1   g539(.A1(new_n740), .A2(new_n716), .A3(new_n633), .A4(new_n737), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n634), .B1(new_n715), .B2(new_n473), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n740), .B1(new_n742), .B2(new_n737), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n744), .A2(new_n451), .A3(new_n654), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n739), .B1(new_n598), .B2(new_n745), .ZN(G1336gat));
  OAI21_X1  g545(.A(G92gat), .B1(new_n738), .B2(new_n661), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n744), .A2(new_n599), .A3(new_n455), .A4(new_n654), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT52), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n747), .A2(new_n748), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(G1337gat));
  OAI21_X1  g552(.A(G99gat), .B1(new_n738), .B2(new_n279), .ZN(new_n754));
  INV_X1    g553(.A(G99gat), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n744), .A2(new_n755), .A3(new_n654), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n756), .B2(new_n702), .ZN(G1338gat));
  OAI21_X1  g556(.A(G106gat), .B1(new_n738), .B2(new_n433), .ZN(new_n758));
  INV_X1    g557(.A(G106gat), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n744), .A2(new_n759), .A3(new_n432), .A4(new_n654), .ZN(new_n760));
  XNOR2_X1  g559(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n761));
  AND3_X1   g560(.A1(new_n758), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n761), .B1(new_n758), .B2(new_n760), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(G1339gat));
  AOI21_X1  g563(.A(new_n538), .B1(new_n537), .B2(new_n540), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n553), .A2(new_n545), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n561), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n565), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n654), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT54), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n653), .B1(new_n647), .B2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n644), .ZN(new_n772));
  AOI211_X1 g571(.A(KEYINPUT10), .B(new_n772), .C1(new_n640), .C2(new_n641), .ZN(new_n773));
  INV_X1    g572(.A(new_n646), .ZN(new_n774));
  OAI22_X1  g573(.A1(new_n773), .A2(new_n774), .B1(new_n635), .B2(new_n256), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n645), .A2(new_n636), .A3(new_n646), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n775), .A2(new_n776), .A3(KEYINPUT54), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n771), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT55), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n649), .A2(new_n653), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n771), .A2(new_n777), .A3(KEYINPUT55), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n769), .B1(new_n783), .B2(new_n566), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT119), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT119), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n769), .B(new_n786), .C1(new_n783), .C2(new_n566), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n785), .A2(new_n634), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n633), .A2(new_n768), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n789), .A2(new_n783), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n595), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n656), .A2(new_n567), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n794), .A2(new_n388), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n467), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n796), .A2(new_n455), .ZN(new_n797));
  INV_X1    g596(.A(G113gat), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n797), .A2(new_n798), .A3(new_n567), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n661), .A2(new_n451), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n800), .A2(new_n702), .ZN(new_n801));
  OAI211_X1 g600(.A(KEYINPUT120), .B(new_n433), .C1(new_n792), .C2(new_n793), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n793), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n633), .B1(new_n784), .B2(KEYINPUT119), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n790), .B1(new_n805), .B2(new_n787), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n806), .B2(new_n595), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT120), .B1(new_n807), .B2(new_n433), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n801), .B1(new_n803), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT121), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT121), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n811), .B(new_n801), .C1(new_n803), .C2(new_n808), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n813), .A2(new_n567), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n799), .B1(new_n814), .B2(new_n798), .ZN(G1340gat));
  INV_X1    g614(.A(KEYINPUT122), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n810), .A2(new_n654), .A3(new_n812), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(G120gat), .ZN(new_n818));
  NOR4_X1   g617(.A1(new_n796), .A2(G120gat), .A3(new_n455), .A4(new_n655), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n816), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  AOI211_X1 g620(.A(KEYINPUT122), .B(new_n819), .C1(new_n817), .C2(G120gat), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n821), .A2(new_n822), .ZN(G1341gat));
  AOI21_X1  g622(.A(G127gat), .B1(new_n797), .B2(new_n595), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n717), .A2(new_n207), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n824), .B1(new_n813), .B2(new_n825), .ZN(G1342gat));
  NOR4_X1   g625(.A1(new_n796), .A2(G134gat), .A3(new_n455), .A4(new_n634), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(KEYINPUT56), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n813), .A2(new_n633), .ZN(new_n829));
  INV_X1    g628(.A(G134gat), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(G1343gat));
  NAND2_X1  g630(.A1(new_n784), .A2(new_n634), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n595), .B1(new_n791), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n432), .B1(new_n833), .B2(new_n793), .ZN(new_n834));
  AOI211_X1 g633(.A(new_n436), .B(new_n800), .C1(new_n834), .C2(KEYINPUT57), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n794), .A2(new_n433), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n835), .A2(new_n838), .A3(new_n567), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(G141gat), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT58), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n436), .A2(new_n433), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n795), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT124), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n795), .A2(KEYINPUT124), .A3(new_n842), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n845), .A2(new_n661), .A3(new_n846), .ZN(new_n847));
  OR2_X1    g646(.A1(new_n566), .A2(G141gat), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n840), .B(new_n841), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n839), .A2(KEYINPUT123), .A3(G141gat), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT123), .B1(new_n839), .B2(G141gat), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n843), .A2(new_n455), .A3(new_n848), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n849), .B1(new_n853), .B2(new_n841), .ZN(G1344gat));
  INV_X1    g653(.A(new_n847), .ZN(new_n855));
  INV_X1    g654(.A(G148gat), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n855), .A2(new_n856), .A3(new_n654), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n836), .A2(KEYINPUT57), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n834), .A2(new_n837), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n436), .A2(new_n800), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n861), .A2(new_n654), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n858), .B1(new_n863), .B2(G148gat), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n835), .A2(new_n838), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n858), .B1(new_n865), .B2(new_n655), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n856), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n857), .B1(new_n864), .B2(new_n867), .ZN(G1345gat));
  NOR3_X1   g667(.A1(new_n865), .A2(new_n333), .A3(new_n717), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n855), .A2(new_n595), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n869), .B1(new_n870), .B2(new_n333), .ZN(G1346gat));
  NOR3_X1   g670(.A1(new_n865), .A2(new_n334), .A3(new_n634), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n855), .A2(new_n633), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n872), .B1(new_n873), .B2(new_n334), .ZN(G1347gat));
  NOR2_X1   g673(.A1(new_n661), .A2(new_n451), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n278), .B(new_n875), .C1(new_n803), .C2(new_n808), .ZN(new_n876));
  OAI21_X1  g675(.A(G169gat), .B1(new_n876), .B2(new_n566), .ZN(new_n877));
  AND4_X1   g676(.A1(new_n388), .A2(new_n807), .A3(new_n455), .A4(new_n467), .ZN(new_n878));
  INV_X1    g677(.A(G169gat), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n878), .A2(new_n879), .A3(new_n567), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n877), .A2(new_n880), .ZN(G1348gat));
  AOI21_X1  g680(.A(G176gat), .B1(new_n878), .B2(new_n654), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n876), .A2(new_n655), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n882), .B1(new_n883), .B2(G176gat), .ZN(G1349gat));
  NAND3_X1  g683(.A1(new_n878), .A2(new_n237), .A3(new_n595), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT125), .ZN(new_n886));
  OAI21_X1  g685(.A(G183gat), .B1(new_n876), .B2(new_n717), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT60), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT60), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n886), .A2(new_n890), .A3(new_n887), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(G1350gat));
  INV_X1    g691(.A(G190gat), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n878), .A2(new_n893), .A3(new_n633), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n876), .A2(new_n634), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT61), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n895), .A2(new_n896), .A3(G190gat), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n896), .B1(new_n895), .B2(G190gat), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(G1351gat));
  INV_X1    g698(.A(KEYINPUT126), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n875), .A2(new_n279), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n901), .B1(new_n859), .B2(new_n860), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n900), .B1(new_n903), .B2(new_n566), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n902), .A2(KEYINPUT126), .A3(new_n567), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n904), .A2(G197gat), .A3(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n794), .A2(new_n451), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n455), .A3(new_n842), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n566), .A2(G197gat), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(G1352gat));
  NOR3_X1   g709(.A1(new_n908), .A2(G204gat), .A3(new_n655), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT62), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n861), .A2(new_n654), .ZN(new_n913));
  OAI21_X1  g712(.A(G204gat), .B1(new_n913), .B2(new_n901), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(G1353gat));
  INV_X1    g714(.A(new_n908), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n303), .A3(new_n595), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n595), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n918), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n919));
  AOI21_X1  g718(.A(KEYINPUT63), .B1(new_n918), .B2(G211gat), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n917), .B1(new_n919), .B2(new_n920), .ZN(G1354gat));
  OAI21_X1  g720(.A(new_n304), .B1(new_n908), .B2(new_n634), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT127), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n922), .B(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n634), .A2(new_n304), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n924), .B1(new_n902), .B2(new_n925), .ZN(G1355gat));
endmodule


