//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 0 0 1 1 0 0 0 0 1 0 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 1 1 0 0 1 0 1 1 1 0 0 0 1 1 1 1 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n568, new_n569, new_n570, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n632,
    new_n633, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1207;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n455), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  AOI22_X1  g036(.A1(new_n461), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT66), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n463), .A2(G2104), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n466), .B1(new_n470), .B2(G137), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n464), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n473), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n475), .A2(new_n476), .A3(G2105), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n472), .A2(new_n478), .ZN(G160));
  OR2_X1    g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n463), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n463), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n486), .B1(G136), .B2(new_n470), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT67), .ZN(G162));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n490), .B1(new_n467), .B2(new_n468), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT69), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n461), .A2(new_n493), .A3(new_n490), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n492), .A2(KEYINPUT4), .A3(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n463), .A2(G114), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(G114), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n500), .A2(new_n502), .A3(KEYINPUT68), .A4(G2104), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n499), .A2(new_n503), .B1(new_n482), .B2(G126), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n491), .A2(KEYINPUT69), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n495), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  OR2_X1    g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OR2_X1    g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(new_n511), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  INV_X1    g094(.A(G50), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  OAI21_X1  g097(.A(G543), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n514), .A2(new_n524), .ZN(G166));
  NAND3_X1  g100(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  INV_X1    g103(.A(G89), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n526), .B(new_n528), .C1(new_n518), .C2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G51), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT70), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n517), .A2(new_n532), .A3(G543), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n523), .A2(KEYINPUT70), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n530), .A2(new_n535), .ZN(G168));
  INV_X1    g111(.A(KEYINPUT71), .ZN(new_n537));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n509), .A2(new_n510), .ZN(new_n539));
  INV_X1    g114(.A(G64), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n515), .A2(new_n516), .B1(new_n509), .B2(new_n510), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n541), .A2(G651), .B1(G90), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n533), .A2(new_n534), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G52), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n537), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n547), .A2(new_n513), .B1(new_n518), .B2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(G52), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n550), .B1(new_n533), .B2(new_n534), .ZN(new_n551));
  NOR3_X1   g126(.A1(new_n549), .A2(new_n551), .A3(KEYINPUT71), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n546), .A2(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  AOI22_X1  g129(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G81), .ZN(new_n556));
  OAI22_X1  g131(.A1(new_n555), .A2(new_n513), .B1(new_n518), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT72), .ZN(new_n559));
  INV_X1    g134(.A(G43), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n560), .B1(new_n533), .B2(new_n534), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n558), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT72), .B1(new_n557), .B2(new_n561), .ZN(new_n564));
  AND2_X1   g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  NAND4_X1  g141(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT73), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(G188));
  INV_X1    g146(.A(G543), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n572), .B1(new_n515), .B2(new_n516), .ZN(new_n573));
  INV_X1    g148(.A(G53), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(KEYINPUT74), .B2(KEYINPUT9), .ZN(new_n575));
  OAI211_X1 g150(.A(new_n573), .B(new_n575), .C1(KEYINPUT74), .C2(KEYINPUT9), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n542), .A2(G91), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT74), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT9), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n578), .B(new_n579), .C1(new_n523), .C2(new_n574), .ZN(new_n580));
  AND3_X1   g155(.A1(new_n576), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(G65), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n582), .B1(new_n509), .B2(new_n510), .ZN(new_n583));
  AND2_X1   g158(.A1(G78), .A2(G543), .ZN(new_n584));
  OR3_X1    g159(.A1(new_n583), .A2(KEYINPUT75), .A3(new_n584), .ZN(new_n585));
  OAI21_X1  g160(.A(KEYINPUT75), .B1(new_n583), .B2(new_n584), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n585), .A2(G651), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n581), .A2(new_n587), .ZN(G299));
  INV_X1    g163(.A(G168), .ZN(G286));
  INV_X1    g164(.A(G166), .ZN(G303));
  OAI21_X1  g165(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n573), .A2(G49), .ZN(new_n592));
  AND2_X1   g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n542), .A2(G87), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(G288));
  AOI22_X1  g170(.A1(new_n511), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(new_n513), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT76), .ZN(new_n598));
  INV_X1    g173(.A(G48), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n523), .B2(new_n599), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n517), .A2(KEYINPUT76), .A3(G48), .A4(G543), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n542), .A2(G86), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n597), .A2(new_n602), .A3(new_n603), .ZN(G305));
  AOI22_X1  g179(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n605), .A2(new_n513), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT77), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n606), .A2(new_n607), .B1(G85), .B2(new_n542), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n544), .A2(G47), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n608), .B(new_n609), .C1(new_n607), .C2(new_n606), .ZN(G290));
  NAND2_X1  g185(.A1(G301), .A2(G868), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n611), .A2(KEYINPUT78), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT10), .ZN(new_n613));
  INV_X1    g188(.A(G92), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n518), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n542), .A2(KEYINPUT10), .A3(G92), .ZN(new_n616));
  NAND2_X1  g191(.A1(G79), .A2(G543), .ZN(new_n617));
  INV_X1    g192(.A(G66), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n539), .B2(new_n618), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n615), .A2(new_n616), .B1(new_n619), .B2(G651), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n544), .A2(G54), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT79), .Z(new_n623));
  INV_X1    g198(.A(G868), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AND2_X1   g200(.A1(new_n611), .A2(KEYINPUT78), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n612), .B1(new_n625), .B2(new_n626), .ZN(G284));
  AOI21_X1  g202(.A(new_n612), .B1(new_n625), .B2(new_n626), .ZN(G321));
  NAND2_X1  g203(.A1(G299), .A2(new_n624), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(new_n624), .B2(G168), .ZN(G297));
  OAI21_X1  g205(.A(new_n629), .B1(new_n624), .B2(G168), .ZN(G280));
  NOR2_X1   g206(.A1(new_n623), .A2(G559), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n622), .B(KEYINPUT79), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n632), .B1(G860), .B2(new_n633), .ZN(G148));
  NAND2_X1  g209(.A1(new_n563), .A2(new_n564), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(new_n624), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(new_n632), .B2(new_n624), .ZN(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g213(.A1(new_n482), .A2(G123), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n463), .A2(G111), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(G135), .B2(new_n470), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT81), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n644), .A2(G2096), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(G2096), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n461), .A2(new_n465), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT12), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2100), .ZN(new_n649));
  XOR2_X1   g224(.A(KEYINPUT80), .B(KEYINPUT13), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n645), .A2(new_n646), .A3(new_n651), .ZN(G156));
  INV_X1    g227(.A(KEYINPUT14), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2427), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2430), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2435), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n657), .B1(new_n656), .B2(new_n655), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1341), .B(G1348), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n658), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2443), .B(G2446), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  AND3_X1   g241(.A1(new_n665), .A2(G14), .A3(new_n666), .ZN(G401));
  INV_X1    g242(.A(KEYINPUT18), .ZN(new_n668));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(KEYINPUT17), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n669), .A2(new_n670), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n668), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G2100), .ZN(new_n675));
  XOR2_X1   g250(.A(G2072), .B(G2078), .Z(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n671), .B2(KEYINPUT18), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2096), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n675), .B(new_n678), .ZN(G227));
  XOR2_X1   g254(.A(G1971), .B(G1976), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  XOR2_X1   g256(.A(G1956), .B(G2474), .Z(new_n682));
  XOR2_X1   g257(.A(G1961), .B(G1966), .Z(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n682), .A2(new_n683), .ZN(new_n686));
  NOR3_X1   g261(.A1(new_n681), .A2(new_n686), .A3(new_n684), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n681), .A2(new_n686), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n689));
  AOI211_X1 g264(.A(new_n685), .B(new_n687), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(new_n688), .B2(new_n689), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G1981), .B(G1986), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G229));
  MUX2_X1   g272(.A(G6), .B(G305), .S(G16), .Z(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT32), .B(G1981), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G23), .ZN(new_n702));
  INV_X1    g277(.A(G288), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(new_n701), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT33), .B(G1976), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n704), .B(new_n705), .Z(new_n706));
  NAND2_X1  g281(.A1(new_n701), .A2(G22), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G166), .B2(new_n701), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n708), .A2(G1971), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(G1971), .ZN(new_n710));
  NOR4_X1   g285(.A1(new_n700), .A2(new_n706), .A3(new_n709), .A4(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT34), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n482), .A2(G119), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n463), .A2(G107), .ZN(new_n716));
  OAI21_X1  g291(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n717));
  INV_X1    g292(.A(G131), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n461), .A2(new_n463), .ZN(new_n719));
  OAI221_X1 g294(.A(new_n715), .B1(new_n716), .B2(new_n717), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  MUX2_X1   g295(.A(G25), .B(new_n720), .S(G29), .Z(new_n721));
  XOR2_X1   g296(.A(KEYINPUT35), .B(G1991), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G1986), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n701), .A2(G24), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G290), .B2(G16), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n723), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n724), .B2(new_n726), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n713), .A2(new_n714), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(KEYINPUT83), .A2(KEYINPUT36), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n729), .B(new_n730), .Z(new_n731));
  NOR2_X1   g306(.A1(G29), .A2(G35), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G162), .B2(G29), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT29), .Z(new_n734));
  INV_X1    g309(.A(G2090), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n736), .A2(KEYINPUT89), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n736), .A2(KEYINPUT89), .ZN(new_n738));
  INV_X1    g313(.A(G29), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G33), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT25), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n461), .A2(G127), .ZN(new_n743));
  NAND2_X1  g318(.A1(G115), .A2(G2104), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n463), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AOI211_X1 g320(.A(new_n742), .B(new_n745), .C1(G139), .C2(new_n470), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n740), .B1(new_n746), .B2(new_n739), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G2072), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n739), .A2(G26), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT28), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n482), .A2(G128), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n463), .A2(G116), .ZN(new_n752));
  OAI21_X1  g327(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n753));
  INV_X1    g328(.A(G140), .ZN(new_n754));
  OAI221_X1 g329(.A(new_n751), .B1(new_n752), .B2(new_n753), .C1(new_n754), .C2(new_n719), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n750), .B1(new_n755), .B2(G29), .ZN(new_n756));
  INV_X1    g331(.A(G2067), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n748), .A2(new_n758), .ZN(new_n759));
  AND2_X1   g334(.A1(KEYINPUT24), .A2(G34), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n739), .B1(KEYINPUT24), .B2(G34), .ZN(new_n761));
  OAI22_X1  g336(.A1(G160), .A2(new_n739), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(G2084), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n701), .A2(G20), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT23), .Z(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G299), .B2(G16), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1956), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT85), .B(KEYINPUT31), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G11), .ZN(new_n770));
  INV_X1    g345(.A(G28), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n771), .A2(KEYINPUT30), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT86), .Z(new_n773));
  AOI21_X1  g348(.A(G29), .B1(new_n771), .B2(KEYINPUT30), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n770), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n644), .B2(new_n739), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n776), .A2(KEYINPUT87), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n759), .A2(new_n764), .A3(new_n768), .A4(new_n777), .ZN(new_n778));
  NOR3_X1   g353(.A1(new_n737), .A2(new_n738), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g354(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT26), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G129), .B2(new_n482), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n470), .A2(G141), .B1(G105), .B2(new_n465), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  MUX2_X1   g359(.A(G32), .B(new_n784), .S(G29), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT27), .ZN(new_n786));
  INV_X1    g361(.A(G1996), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n701), .A2(G21), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G168), .B2(new_n701), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(G1966), .Z(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n776), .B2(KEYINPUT87), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n739), .A2(G27), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G164), .B2(new_n739), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT88), .Z(new_n796));
  INV_X1    g371(.A(G2078), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n633), .A2(new_n701), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G4), .B2(new_n701), .ZN(new_n801));
  INV_X1    g376(.A(G1348), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n793), .A2(new_n798), .A3(new_n799), .A4(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(G5), .A2(G16), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G171), .B2(G16), .ZN(new_n806));
  INV_X1    g381(.A(G1961), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n802), .B2(new_n801), .ZN(new_n809));
  INV_X1    g384(.A(G19), .ZN(new_n810));
  OR3_X1    g385(.A1(new_n810), .A2(KEYINPUT84), .A3(G16), .ZN(new_n811));
  OAI21_X1  g386(.A(KEYINPUT84), .B1(new_n810), .B2(G16), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n811), .B(new_n812), .C1(new_n565), .C2(new_n701), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G1341), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n734), .A2(new_n735), .ZN(new_n815));
  NOR4_X1   g390(.A1(new_n804), .A2(new_n809), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n731), .A2(new_n779), .A3(new_n816), .ZN(G150));
  INV_X1    g392(.A(G150), .ZN(G311));
  NAND2_X1  g393(.A1(new_n633), .A2(G559), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT92), .B(KEYINPUT38), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n819), .B(new_n820), .Z(new_n821));
  NOR2_X1   g396(.A1(new_n557), .A2(new_n561), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n823), .A2(new_n513), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT91), .ZN(new_n826));
  INV_X1    g401(.A(G55), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(new_n533), .B2(new_n534), .ZN(new_n828));
  XOR2_X1   g403(.A(KEYINPUT90), .B(G93), .Z(new_n829));
  AND2_X1   g404(.A1(new_n542), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n826), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  NOR3_X1   g407(.A1(new_n828), .A2(new_n830), .A3(new_n826), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n822), .B(new_n825), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n544), .A2(G55), .B1(new_n542), .B2(new_n829), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(KEYINPUT91), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n824), .B1(new_n836), .B2(new_n831), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n834), .B1(new_n565), .B2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n821), .B(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT39), .ZN(new_n841));
  AOI21_X1  g416(.A(G860), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n841), .B2(new_n840), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n825), .B1(new_n832), .B2(new_n833), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(G860), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT37), .Z(new_n846));
  NAND2_X1  g421(.A1(new_n843), .A2(new_n846), .ZN(G145));
  INV_X1    g422(.A(KEYINPUT93), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n644), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(G162), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n850), .A2(G160), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(G160), .ZN(new_n852));
  OAI21_X1  g427(.A(KEYINPUT98), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n850), .A2(G160), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT98), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n850), .A2(G160), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT96), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n720), .B(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n648), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n482), .A2(G130), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n463), .A2(G118), .ZN(new_n862));
  OAI21_X1  g437(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT95), .ZN(new_n864));
  AND3_X1   g439(.A1(new_n470), .A2(new_n864), .A3(G142), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n864), .B1(new_n470), .B2(G142), .ZN(new_n866));
  OAI221_X1 g441(.A(new_n861), .B1(new_n862), .B2(new_n863), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n860), .B(new_n867), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n868), .A2(KEYINPUT97), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(KEYINPUT97), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n746), .B(new_n784), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n755), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n492), .A2(KEYINPUT4), .A3(new_n494), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n499), .A2(new_n503), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n482), .A2(G126), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n506), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(KEYINPUT94), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT94), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n495), .A2(new_n504), .A3(new_n879), .A4(new_n506), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n873), .B(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n871), .A2(new_n883), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n860), .B(new_n867), .Z(new_n885));
  NAND2_X1  g460(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n853), .A2(new_n857), .A3(new_n884), .A4(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n851), .A2(new_n852), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n871), .A2(new_n883), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n882), .B1(new_n869), .B2(new_n870), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(G37), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n887), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g469(.A(KEYINPUT101), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n895), .B1(new_n837), .B2(G868), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n632), .B(new_n839), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n622), .A2(G299), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n620), .A2(new_n581), .A3(new_n587), .A4(new_n621), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT99), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n897), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT41), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n905), .B1(new_n898), .B2(new_n899), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n898), .A2(new_n905), .A3(new_n899), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n897), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(KEYINPUT42), .B1(new_n904), .B2(new_n910), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n897), .A2(new_n909), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT42), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(new_n913), .A3(new_n903), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(G290), .B(G305), .ZN(new_n916));
  XOR2_X1   g491(.A(G166), .B(G288), .Z(new_n917));
  XNOR2_X1  g492(.A(new_n916), .B(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT100), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n624), .B1(new_n915), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n911), .A2(new_n914), .A3(new_n920), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n896), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n904), .A2(new_n910), .A3(KEYINPUT42), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n913), .B1(new_n912), .B2(new_n903), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n921), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AND4_X1   g502(.A1(KEYINPUT101), .A2(new_n927), .A3(G868), .A4(new_n923), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n924), .A2(new_n928), .ZN(G295));
  NOR2_X1   g504(.A1(new_n924), .A2(new_n928), .ZN(G331));
  INV_X1    g505(.A(KEYINPUT104), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n908), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n906), .B1(new_n931), .B2(new_n908), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n543), .A2(new_n537), .A3(new_n545), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT71), .B1(new_n549), .B2(new_n551), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(new_n935), .A3(G168), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(G168), .B1(new_n934), .B2(new_n935), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n838), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(G286), .B1(new_n546), .B2(new_n552), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n936), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n844), .A2(new_n635), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n942), .A2(new_n943), .A3(new_n834), .ZN(new_n944));
  AOI22_X1  g519(.A1(new_n932), .A2(new_n933), .B1(new_n940), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT103), .B1(new_n838), .B2(new_n939), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n940), .A2(new_n944), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n946), .B1(new_n947), .B2(KEYINPUT103), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n945), .B1(new_n948), .B2(new_n901), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT105), .B1(new_n949), .B2(new_n918), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT103), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n952), .B1(new_n940), .B2(new_n944), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n953), .A2(new_n902), .A3(new_n946), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n951), .B(new_n919), .C1(new_n954), .C2(new_n945), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n909), .B1(new_n953), .B2(new_n946), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n947), .A2(new_n900), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n956), .A2(new_n918), .A3(new_n957), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n950), .A2(new_n892), .A3(new_n955), .A4(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT107), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n958), .A2(new_n892), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n961), .A2(new_n962), .A3(new_n950), .A4(new_n955), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n960), .A2(KEYINPUT43), .A3(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n958), .A2(new_n892), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n918), .B1(new_n956), .B2(new_n957), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XOR2_X1   g543(.A(KEYINPUT102), .B(KEYINPUT43), .Z(new_n969));
  AOI21_X1  g544(.A(new_n965), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n964), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n961), .A2(new_n955), .A3(new_n950), .A4(new_n969), .ZN(new_n972));
  INV_X1    g547(.A(new_n969), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n973), .B1(new_n966), .B2(new_n967), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT106), .B1(new_n975), .B2(new_n965), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT106), .ZN(new_n977));
  AOI211_X1 g552(.A(new_n977), .B(KEYINPUT44), .C1(new_n972), .C2(new_n974), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n971), .B1(new_n976), .B2(new_n978), .ZN(G397));
  XNOR2_X1  g554(.A(KEYINPUT108), .B(G1384), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n878), .A2(new_n880), .A3(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n464), .A2(new_n471), .A3(new_n477), .A4(G40), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n784), .B(new_n787), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n755), .B(new_n757), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n722), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n720), .B(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n988), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(G290), .B(new_n724), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n994), .B1(new_n987), .B2(new_n995), .ZN(new_n996));
  XOR2_X1   g571(.A(new_n996), .B(KEYINPUT109), .Z(new_n997));
  XOR2_X1   g572(.A(G299), .B(KEYINPUT57), .Z(new_n998));
  INV_X1    g573(.A(G1384), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n999), .B1(new_n874), .B2(new_n877), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n1000), .A2(KEYINPUT110), .A3(new_n983), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n986), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT45), .B1(new_n507), .B2(new_n999), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1003), .A2(KEYINPUT110), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n980), .A2(new_n983), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n878), .A2(new_n880), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT111), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT111), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n878), .A2(new_n1009), .A3(new_n880), .A4(new_n1006), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(KEYINPUT56), .B(G2072), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1005), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1000), .A2(KEYINPUT50), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT50), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n507), .A2(new_n1015), .A3(new_n999), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1014), .A2(new_n986), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G1956), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n998), .B1(new_n1013), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1013), .A2(new_n998), .A3(new_n1019), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1000), .A2(new_n985), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n1017), .A2(new_n802), .B1(new_n757), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1023), .A2(new_n623), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1020), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT61), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1021), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1026), .B1(new_n1027), .B2(new_n1020), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1013), .A2(new_n1019), .ZN(new_n1029));
  INV_X1    g604(.A(new_n998), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1031), .A2(KEYINPUT61), .A3(new_n1021), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1028), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1005), .A2(new_n787), .A3(new_n1011), .ZN(new_n1034));
  XOR2_X1   g609(.A(KEYINPUT58), .B(G1341), .Z(new_n1035));
  OAI21_X1  g610(.A(new_n1035), .B1(new_n1000), .B2(new_n985), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n565), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT59), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n633), .A2(KEYINPUT60), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1041), .A2(new_n1023), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1041), .A2(new_n1023), .ZN(new_n1043));
  OAI22_X1  g618(.A1(new_n1042), .A2(new_n1043), .B1(KEYINPUT60), .B2(new_n633), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1037), .A2(KEYINPUT59), .A3(new_n565), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1040), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1025), .B1(new_n1033), .B2(new_n1046), .ZN(new_n1047));
  XOR2_X1   g622(.A(KEYINPUT121), .B(KEYINPUT54), .Z(new_n1048));
  INV_X1    g623(.A(new_n1004), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n985), .B1(new_n1003), .B2(KEYINPUT110), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1011), .A2(new_n797), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1017), .A2(new_n807), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n999), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n1055), .A2(new_n1003), .A3(new_n985), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(KEYINPUT53), .A3(new_n797), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1053), .A2(new_n1054), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(G171), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n1051), .A2(new_n1052), .B1(new_n807), .B2(new_n1017), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n463), .B1(new_n475), .B2(KEYINPUT122), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(KEYINPUT122), .B2(new_n475), .ZN(new_n1062));
  NAND2_X1  g637(.A1(KEYINPUT53), .A2(G40), .ZN(new_n1063));
  OR2_X1    g638(.A1(KEYINPUT123), .A2(G2078), .ZN(new_n1064));
  NAND2_X1  g639(.A1(KEYINPUT123), .A2(G2078), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1063), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1062), .A2(new_n471), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1067), .B1(new_n982), .B2(new_n983), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1011), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT124), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT124), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1011), .A2(new_n1071), .A3(new_n1068), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1060), .A2(new_n1073), .A3(G301), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1048), .B1(new_n1059), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G8), .ZN(new_n1076));
  NOR2_X1   g651(.A1(G166), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT55), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT112), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OR2_X1    g655(.A1(new_n1077), .A2(KEYINPUT55), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1077), .A2(KEYINPUT112), .A3(KEYINPUT55), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1005), .A2(new_n1011), .ZN(new_n1085));
  INV_X1    g660(.A(G1971), .ZN(new_n1086));
  OR2_X1    g661(.A1(new_n1017), .A2(KEYINPUT118), .ZN(new_n1087));
  AOI21_X1  g662(.A(G2090), .B1(new_n1017), .B2(KEYINPUT118), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1085), .A2(new_n1086), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1084), .B1(new_n1089), .B2(new_n1076), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1014), .A2(new_n986), .A3(new_n763), .A4(new_n1016), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n985), .B1(new_n1000), .B2(new_n983), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n999), .ZN(new_n1094));
  AOI21_X1  g669(.A(G1966), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(G8), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(G168), .A2(new_n1076), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT51), .B1(new_n1098), .B2(KEYINPUT120), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1096), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1091), .B1(new_n1056), .B2(G1966), .ZN(new_n1102));
  OAI211_X1 g677(.A(G8), .B(new_n1099), .C1(new_n1102), .C2(G286), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1097), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1101), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(G1971), .B1(new_n1005), .B2(new_n1011), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1017), .A2(G2090), .ZN(new_n1107));
  OAI211_X1 g682(.A(G8), .B(new_n1083), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT114), .B(G86), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n600), .A2(new_n601), .B1(new_n542), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n597), .B1(new_n1110), .B2(KEYINPUT115), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n542), .A2(new_n1109), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n602), .A2(KEYINPUT115), .A3(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(G1981), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(G1981), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n597), .A2(new_n1115), .A3(new_n602), .A4(new_n603), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1114), .A2(KEYINPUT49), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT116), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT116), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1114), .A2(new_n1119), .A3(KEYINPUT49), .A4(new_n1116), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1022), .A2(new_n1076), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT49), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n596), .A2(new_n513), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n602), .A2(new_n1112), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT115), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1123), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1110), .A2(KEYINPUT115), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1115), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1116), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1122), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1118), .A2(new_n1120), .A3(new_n1121), .A4(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n593), .A2(G1976), .A3(new_n594), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT113), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(G1976), .B1(new_n593), .B2(new_n594), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1121), .B(new_n1134), .C1(KEYINPUT52), .C2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1134), .B(G8), .C1(new_n1000), .C2(new_n985), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1135), .B(G8), .C1(new_n1000), .C2(new_n985), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT52), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1136), .A2(new_n1140), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1131), .A2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1090), .A2(new_n1105), .A3(new_n1108), .A4(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1075), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1060), .A2(G301), .A3(new_n1057), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n1060), .A2(new_n1073), .ZN(new_n1146));
  OAI211_X1 g721(.A(KEYINPUT54), .B(new_n1145), .C1(new_n1146), .C2(G301), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1047), .A2(new_n1144), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(G1976), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1131), .A2(new_n1149), .A3(new_n703), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n1116), .ZN(new_n1151));
  XOR2_X1   g726(.A(new_n1121), .B(KEYINPUT117), .Z(new_n1152));
  INV_X1    g727(.A(new_n1108), .ZN(new_n1153));
  AOI22_X1  g728(.A1(new_n1151), .A2(new_n1152), .B1(new_n1153), .B2(new_n1142), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT126), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1105), .A2(KEYINPUT62), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(KEYINPUT125), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT125), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1105), .A2(new_n1158), .A3(KEYINPUT62), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  AND2_X1   g735(.A1(new_n1142), .A2(new_n1108), .ZN(new_n1161));
  AOI21_X1  g736(.A(G301), .B1(new_n1060), .B2(new_n1057), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT62), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1101), .A2(new_n1103), .A3(new_n1163), .A4(new_n1104), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1161), .A2(new_n1090), .A3(new_n1162), .A4(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1155), .B1(new_n1160), .B2(new_n1165), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1086), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1076), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1142), .B(new_n1108), .C1(new_n1171), .C2(new_n1083), .ZN(new_n1172));
  AND4_X1   g747(.A1(new_n1163), .A2(new_n1101), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1173));
  NOR3_X1   g748(.A1(new_n1172), .A2(new_n1173), .A3(new_n1059), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1174), .A2(KEYINPUT126), .A3(new_n1159), .A4(new_n1157), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1148), .A2(new_n1154), .A3(new_n1166), .A4(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT63), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1102), .A2(G8), .A3(G168), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1177), .B1(new_n1172), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT119), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g756(.A(KEYINPUT119), .B(new_n1177), .C1(new_n1172), .C2(new_n1178), .ZN(new_n1182));
  OAI21_X1  g757(.A(G8), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1183));
  AOI211_X1 g758(.A(new_n1177), .B(new_n1178), .C1(new_n1183), .C2(new_n1084), .ZN(new_n1184));
  AOI22_X1  g759(.A1(new_n1181), .A2(new_n1182), .B1(new_n1161), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n997), .B1(new_n1176), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(new_n990), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n988), .B1(new_n784), .B2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n987), .A2(G1996), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1189), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n1190), .A2(KEYINPUT46), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1190), .A2(KEYINPUT46), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1188), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  XOR2_X1   g768(.A(new_n1193), .B(KEYINPUT47), .Z(new_n1194));
  NOR2_X1   g769(.A1(new_n720), .A2(new_n992), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n1195), .B(KEYINPUT127), .ZN(new_n1196));
  OAI22_X1  g771(.A1(new_n991), .A2(new_n1196), .B1(G2067), .B2(new_n755), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n988), .A2(new_n1197), .ZN(new_n1198));
  OR3_X1    g773(.A1(new_n987), .A2(G1986), .A3(G290), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1199), .ZN(new_n1200));
  AND2_X1   g775(.A1(new_n1200), .A2(KEYINPUT48), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n994), .B1(new_n1200), .B2(KEYINPUT48), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1198), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n1194), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1186), .A2(new_n1204), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g780(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1207));
  NAND3_X1  g781(.A1(new_n1207), .A2(new_n893), .A3(new_n975), .ZN(G225));
  INV_X1    g782(.A(G225), .ZN(G308));
endmodule


