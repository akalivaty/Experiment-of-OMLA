

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793;

  XNOR2_X1 U380 ( .A(n663), .B(n662), .ZN(n664) );
  AND2_X1 U381 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U382 ( .A(n457), .B(KEYINPUT96), .ZN(n561) );
  BUF_X1 U383 ( .A(G128), .Z(n359) );
  XOR2_X2 U384 ( .A(n562), .B(KEYINPUT34), .Z(n563) );
  XNOR2_X2 U385 ( .A(n367), .B(n491), .ZN(n687) );
  XNOR2_X2 U386 ( .A(n427), .B(KEYINPUT105), .ZN(n736) );
  XNOR2_X1 U387 ( .A(n534), .B(n533), .ZN(n558) );
  XNOR2_X2 U388 ( .A(n578), .B(n577), .ZN(n677) );
  XNOR2_X2 U389 ( .A(n392), .B(G146), .ZN(n368) );
  XNOR2_X2 U390 ( .A(n367), .B(n482), .ZN(n741) );
  XNOR2_X1 U391 ( .A(KEYINPUT64), .B(G953), .ZN(n781) );
  NOR2_X1 U392 ( .A1(n729), .A2(n627), .ZN(n618) );
  AND2_X4 U393 ( .A1(n402), .A2(n401), .ZN(n685) );
  XNOR2_X2 U394 ( .A(n368), .B(n476), .ZN(n367) );
  XNOR2_X2 U395 ( .A(n611), .B(n407), .ZN(n790) );
  NOR2_X1 U396 ( .A1(n388), .A2(n387), .ZN(n643) );
  BUF_X1 U397 ( .A(n543), .Z(n615) );
  BUF_X1 U398 ( .A(n569), .Z(n704) );
  XNOR2_X1 U399 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U400 ( .A(n687), .B(n686), .ZN(n688) );
  XNOR2_X1 U401 ( .A(n489), .B(n413), .ZN(n770) );
  NAND2_X1 U402 ( .A1(n552), .A2(n431), .ZN(n554) );
  XNOR2_X1 U403 ( .A(n410), .B(n770), .ZN(n671) );
  INV_X1 U404 ( .A(n685), .ZN(n360) );
  INV_X1 U405 ( .A(n360), .ZN(n361) );
  XNOR2_X2 U406 ( .A(n776), .B(n436), .ZN(n476) );
  BUF_X1 U407 ( .A(n655), .Z(n656) );
  XNOR2_X1 U408 ( .A(n493), .B(n492), .ZN(n569) );
  XNOR2_X1 U409 ( .A(n459), .B(n458), .ZN(n524) );
  XOR2_X1 U410 ( .A(G137), .B(G140), .Z(n477) );
  XNOR2_X1 U411 ( .A(G902), .B(KEYINPUT15), .ZN(n651) );
  XNOR2_X1 U412 ( .A(n476), .B(n411), .ZN(n410) );
  XNOR2_X1 U413 ( .A(n435), .B(n412), .ZN(n411) );
  XNOR2_X1 U414 ( .A(n604), .B(n603), .ZN(n378) );
  INV_X1 U415 ( .A(KEYINPUT30), .ZN(n603) );
  NAND2_X1 U416 ( .A1(n386), .A2(n384), .ZN(n387) );
  OR2_X1 U417 ( .A1(n790), .A2(n619), .ZN(n386) );
  XNOR2_X1 U418 ( .A(n364), .B(n601), .ZN(n655) );
  XNOR2_X1 U419 ( .A(n472), .B(n471), .ZN(n543) );
  BUF_X1 U420 ( .A(n652), .Z(n779) );
  XNOR2_X1 U421 ( .A(G119), .B(G110), .ZN(n461) );
  INV_X1 U422 ( .A(KEYINPUT23), .ZN(n419) );
  XNOR2_X1 U423 ( .A(n524), .B(n460), .ZN(n775) );
  XNOR2_X1 U424 ( .A(G104), .B(G107), .ZN(n478) );
  AND2_X1 U425 ( .A1(n376), .A2(n373), .ZN(n372) );
  NOR2_X1 U426 ( .A1(n371), .A2(n609), .ZN(n370) );
  NAND2_X1 U427 ( .A1(n628), .A2(n453), .ZN(n456) );
  XNOR2_X1 U428 ( .A(n569), .B(n568), .ZN(n613) );
  AND2_X1 U429 ( .A1(n543), .A2(n550), .ZN(n416) );
  XNOR2_X1 U430 ( .A(n440), .B(n414), .ZN(n413) );
  XNOR2_X1 U431 ( .A(n518), .B(n501), .ZN(n414) );
  XNOR2_X1 U432 ( .A(n508), .B(n507), .ZN(n658) );
  NAND2_X1 U433 ( .A1(n403), .A2(n363), .ZN(n402) );
  NAND2_X1 U434 ( .A1(n734), .A2(n733), .ZN(n383) );
  INV_X1 U435 ( .A(KEYINPUT114), .ZN(n382) );
  OR2_X1 U436 ( .A1(n759), .A2(n746), .ZN(n588) );
  XNOR2_X1 U437 ( .A(n432), .B(G125), .ZN(n459) );
  INV_X1 U438 ( .A(G146), .ZN(n432) );
  NAND2_X1 U439 ( .A1(n389), .A2(n642), .ZN(n388) );
  NAND2_X1 U440 ( .A1(G234), .A2(G237), .ZN(n446) );
  INV_X1 U441 ( .A(G237), .ZN(n441) );
  XNOR2_X1 U442 ( .A(G143), .B(G122), .ZN(n519) );
  INV_X1 U443 ( .A(G134), .ZN(n428) );
  XNOR2_X1 U444 ( .A(n459), .B(n433), .ZN(n412) );
  XNOR2_X1 U445 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n433) );
  NAND2_X1 U446 ( .A1(n615), .A2(KEYINPUT28), .ZN(n396) );
  NOR2_X1 U447 ( .A1(n614), .A2(n398), .ZN(n397) );
  NAND2_X1 U448 ( .A1(n400), .A2(n399), .ZN(n398) );
  INV_X1 U449 ( .A(KEYINPUT28), .ZN(n399) );
  OR2_X1 U450 ( .A1(n584), .A2(n585), .ZN(n714) );
  NAND2_X1 U451 ( .A1(n375), .A2(n608), .ZN(n374) );
  INV_X1 U452 ( .A(n609), .ZN(n375) );
  NOR2_X1 U453 ( .A1(n445), .A2(n362), .ZN(n421) );
  BUF_X1 U454 ( .A(n534), .Z(n606) );
  INV_X1 U455 ( .A(G902), .ZN(n528) );
  NOR2_X1 U456 ( .A1(G953), .A2(G237), .ZN(n511) );
  XNOR2_X1 U457 ( .A(G137), .B(G113), .ZN(n485) );
  XNOR2_X1 U458 ( .A(n415), .B(n438), .ZN(n489) );
  XNOR2_X1 U459 ( .A(n437), .B(KEYINPUT77), .ZN(n415) );
  XNOR2_X1 U460 ( .A(KEYINPUT3), .B(G119), .ZN(n437) );
  XNOR2_X1 U461 ( .A(KEYINPUT79), .B(KEYINPUT16), .ZN(n439) );
  NAND2_X1 U462 ( .A1(n394), .A2(n393), .ZN(n627) );
  NAND2_X1 U463 ( .A1(n614), .A2(KEYINPUT28), .ZN(n393) );
  NOR2_X1 U464 ( .A1(n397), .A2(n395), .ZN(n394) );
  NAND2_X1 U465 ( .A1(n616), .A2(n396), .ZN(n395) );
  XNOR2_X1 U466 ( .A(n466), .B(n417), .ZN(n680) );
  XNOR2_X1 U467 ( .A(n775), .B(n418), .ZN(n417) );
  XNOR2_X1 U468 ( .A(n461), .B(n419), .ZN(n418) );
  XNOR2_X1 U469 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U470 ( .A(n660), .B(KEYINPUT92), .ZN(n690) );
  INV_X1 U471 ( .A(KEYINPUT40), .ZN(n407) );
  AND2_X1 U472 ( .A1(n644), .A2(n756), .ZN(n611) );
  BUF_X1 U473 ( .A(n597), .Z(n737) );
  NAND2_X1 U474 ( .A1(n378), .A2(n608), .ZN(n622) );
  AND2_X1 U475 ( .A1(n570), .A2(n573), .ZN(n426) );
  INV_X1 U476 ( .A(G110), .ZN(n735) );
  XNOR2_X1 U477 ( .A(n409), .B(n408), .ZN(n661) );
  INV_X1 U478 ( .A(n658), .ZN(n408) );
  INV_X1 U479 ( .A(KEYINPUT53), .ZN(n379) );
  XNOR2_X1 U480 ( .A(KEYINPUT68), .B(KEYINPUT19), .ZN(n362) );
  OR2_X1 U481 ( .A1(n651), .A2(n650), .ZN(n363) );
  NAND2_X1 U482 ( .A1(n365), .A2(n600), .ZN(n364) );
  XNOR2_X1 U483 ( .A(n366), .B(KEYINPUT89), .ZN(n365) );
  NAND2_X1 U484 ( .A1(n595), .A2(n596), .ZN(n366) );
  XNOR2_X2 U485 ( .A(n523), .B(n428), .ZN(n392) );
  NAND2_X1 U486 ( .A1(n372), .A2(n369), .ZN(n644) );
  NAND2_X1 U487 ( .A1(n378), .A2(n370), .ZN(n369) );
  NAND2_X1 U488 ( .A1(n608), .A2(n610), .ZN(n371) );
  NAND2_X1 U489 ( .A1(n374), .A2(KEYINPUT39), .ZN(n373) );
  NAND2_X1 U490 ( .A1(n377), .A2(KEYINPUT39), .ZN(n376) );
  INV_X1 U491 ( .A(n378), .ZN(n377) );
  XNOR2_X1 U492 ( .A(n380), .B(n379), .ZN(G75) );
  NAND2_X1 U493 ( .A1(n381), .A2(n764), .ZN(n380) );
  XNOR2_X1 U494 ( .A(n383), .B(n382), .ZN(n381) );
  NAND2_X1 U495 ( .A1(n790), .A2(n385), .ZN(n384) );
  AND2_X1 U496 ( .A1(n793), .A2(n619), .ZN(n385) );
  NAND2_X1 U497 ( .A1(n391), .A2(n390), .ZN(n389) );
  INV_X1 U498 ( .A(n619), .ZN(n390) );
  INV_X1 U499 ( .A(n793), .ZN(n391) );
  OR2_X2 U500 ( .A1(n677), .A2(n736), .ZN(n598) );
  BUF_X1 U501 ( .A(n552), .Z(n582) );
  INV_X1 U502 ( .A(n695), .ZN(n401) );
  NOR2_X2 U503 ( .A1(n655), .A2(n651), .ZN(n602) );
  XNOR2_X1 U504 ( .A(n392), .B(n776), .ZN(n777) );
  INV_X1 U505 ( .A(n615), .ZN(n400) );
  NAND2_X1 U506 ( .A1(n598), .A2(KEYINPUT44), .ZN(n592) );
  NAND2_X1 U507 ( .A1(n598), .A2(KEYINPUT66), .ZN(n579) );
  NAND2_X1 U508 ( .A1(n404), .A2(n653), .ZN(n403) );
  XNOR2_X1 U509 ( .A(n602), .B(n405), .ZN(n404) );
  INV_X1 U510 ( .A(KEYINPUT87), .ZN(n405) );
  NAND2_X1 U511 ( .A1(n575), .A2(n406), .ZN(n578) );
  NAND2_X1 U512 ( .A1(n406), .A2(n426), .ZN(n427) );
  AND2_X1 U513 ( .A1(n406), .A2(n573), .ZN(n571) );
  XNOR2_X2 U514 ( .A(n554), .B(n553), .ZN(n406) );
  NAND2_X1 U515 ( .A1(n361), .A2(G478), .ZN(n409) );
  NOR2_X2 U516 ( .A1(n657), .A2(n656), .ZN(n695) );
  NOR2_X2 U517 ( .A1(n581), .A2(n572), .ZN(n560) );
  XNOR2_X2 U518 ( .A(n559), .B(KEYINPUT80), .ZN(n581) );
  NOR2_X2 U519 ( .A1(n719), .A2(n561), .ZN(n564) );
  XNOR2_X2 U520 ( .A(n704), .B(n544), .ZN(n572) );
  XNOR2_X2 U521 ( .A(n498), .B(KEYINPUT4), .ZN(n776) );
  NAND2_X1 U522 ( .A1(n558), .A2(n416), .ZN(n559) );
  NAND2_X1 U523 ( .A1(n616), .A2(n416), .ZN(n495) );
  AND2_X1 U524 ( .A1(n607), .A2(n416), .ZN(n608) );
  NOR2_X1 U525 ( .A1(n697), .A2(n416), .ZN(n699) );
  NAND2_X2 U526 ( .A1(n423), .A2(n420), .ZN(n628) );
  NAND2_X1 U527 ( .A1(n422), .A2(n421), .ZN(n420) );
  INV_X1 U528 ( .A(n548), .ZN(n422) );
  AND2_X2 U529 ( .A1(n425), .A2(n424), .ZN(n423) );
  NAND2_X1 U530 ( .A1(n445), .A2(n362), .ZN(n424) );
  NAND2_X1 U531 ( .A1(n548), .A2(n362), .ZN(n425) );
  XNOR2_X2 U532 ( .A(n443), .B(n442), .ZN(n548) );
  XNOR2_X2 U533 ( .A(n429), .B(KEYINPUT72), .ZN(n523) );
  XNOR2_X2 U534 ( .A(G131), .B(KEYINPUT73), .ZN(n429) );
  BUF_X1 U535 ( .A(n548), .Z(n623) );
  OR2_X1 U536 ( .A1(n781), .A2(n480), .ZN(n430) );
  AND2_X1 U537 ( .A1(n551), .A2(n550), .ZN(n431) );
  XNOR2_X1 U538 ( .A(KEYINPUT65), .B(KEYINPUT46), .ZN(n619) );
  INV_X1 U539 ( .A(n477), .ZN(n460) );
  INV_X1 U540 ( .A(KEYINPUT10), .ZN(n458) );
  XNOR2_X1 U541 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U542 ( .A(n481), .B(n430), .ZN(n482) );
  INV_X1 U543 ( .A(KEYINPUT39), .ZN(n610) );
  XNOR2_X1 U544 ( .A(n505), .B(n504), .ZN(n508) );
  INV_X1 U545 ( .A(G224), .ZN(n434) );
  NOR2_X1 U546 ( .A1(n781), .A2(n434), .ZN(n435) );
  XNOR2_X2 U547 ( .A(G143), .B(G128), .ZN(n498) );
  XNOR2_X1 U548 ( .A(KEYINPUT70), .B(G101), .ZN(n436) );
  XNOR2_X1 U549 ( .A(G116), .B(KEYINPUT76), .ZN(n438) );
  XNOR2_X2 U550 ( .A(G113), .B(G104), .ZN(n518) );
  XNOR2_X2 U551 ( .A(G122), .B(G107), .ZN(n501) );
  XNOR2_X1 U552 ( .A(n439), .B(n735), .ZN(n440) );
  NAND2_X1 U553 ( .A1(n671), .A2(n651), .ZN(n443) );
  NAND2_X1 U554 ( .A1(n528), .A2(n441), .ZN(n444) );
  NAND2_X1 U555 ( .A1(n444), .A2(G210), .ZN(n442) );
  NAND2_X1 U556 ( .A1(n444), .A2(G214), .ZN(n711) );
  INV_X1 U557 ( .A(n711), .ZN(n445) );
  XNOR2_X1 U558 ( .A(n446), .B(KEYINPUT14), .ZN(n450) );
  NAND2_X1 U559 ( .A1(n450), .A2(G902), .ZN(n447) );
  XNOR2_X1 U560 ( .A(n447), .B(KEYINPUT94), .ZN(n536) );
  INV_X1 U561 ( .A(G953), .ZN(n764) );
  NOR2_X1 U562 ( .A1(n764), .A2(G898), .ZN(n448) );
  XNOR2_X1 U563 ( .A(n448), .B(KEYINPUT93), .ZN(n771) );
  NOR2_X1 U564 ( .A1(n536), .A2(n771), .ZN(n449) );
  XNOR2_X1 U565 ( .A(n449), .B(KEYINPUT95), .ZN(n452) );
  NAND2_X1 U566 ( .A1(G952), .A2(n450), .ZN(n726) );
  NOR2_X1 U567 ( .A1(n726), .A2(G953), .ZN(n539) );
  INV_X1 U568 ( .A(n539), .ZN(n451) );
  NAND2_X1 U569 ( .A1(n452), .A2(n451), .ZN(n453) );
  INV_X1 U570 ( .A(KEYINPUT90), .ZN(n454) );
  XNOR2_X1 U571 ( .A(n454), .B(KEYINPUT0), .ZN(n455) );
  XNOR2_X2 U572 ( .A(n456), .B(n455), .ZN(n552) );
  INV_X1 U573 ( .A(n552), .ZN(n457) );
  INV_X1 U574 ( .A(n561), .ZN(n497) );
  INV_X1 U575 ( .A(n781), .ZN(n535) );
  NAND2_X1 U576 ( .A1(n535), .A2(G234), .ZN(n463) );
  XNOR2_X1 U577 ( .A(KEYINPUT71), .B(KEYINPUT8), .ZN(n462) );
  XNOR2_X1 U578 ( .A(n463), .B(n462), .ZN(n506) );
  AND2_X1 U579 ( .A1(n506), .A2(G221), .ZN(n465) );
  XOR2_X1 U580 ( .A(n359), .B(KEYINPUT24), .Z(n464) );
  NAND2_X1 U581 ( .A1(n680), .A2(n528), .ZN(n472) );
  XOR2_X1 U582 ( .A(KEYINPUT82), .B(KEYINPUT25), .Z(n470) );
  XOR2_X1 U583 ( .A(KEYINPUT97), .B(KEYINPUT20), .Z(n468) );
  NAND2_X1 U584 ( .A1(G234), .A2(n651), .ZN(n467) );
  XNOR2_X1 U585 ( .A(n468), .B(n467), .ZN(n473) );
  NAND2_X1 U586 ( .A1(n473), .A2(G217), .ZN(n469) );
  XNOR2_X1 U587 ( .A(n470), .B(n469), .ZN(n471) );
  AND2_X1 U588 ( .A1(n473), .A2(G221), .ZN(n475) );
  INV_X1 U589 ( .A(KEYINPUT21), .ZN(n474) );
  XNOR2_X1 U590 ( .A(n475), .B(n474), .ZN(n701) );
  INV_X1 U591 ( .A(n701), .ZN(n550) );
  XOR2_X1 U592 ( .A(n477), .B(G110), .Z(n479) );
  XNOR2_X1 U593 ( .A(n479), .B(n478), .ZN(n481) );
  INV_X1 U594 ( .A(G227), .ZN(n480) );
  NAND2_X1 U595 ( .A1(n741), .A2(n528), .ZN(n484) );
  XNOR2_X1 U596 ( .A(KEYINPUT75), .B(G469), .ZN(n483) );
  XNOR2_X2 U597 ( .A(n484), .B(n483), .ZN(n534) );
  INV_X1 U598 ( .A(n606), .ZN(n616) );
  XOR2_X1 U599 ( .A(KEYINPUT5), .B(KEYINPUT81), .Z(n486) );
  XNOR2_X1 U600 ( .A(n486), .B(n485), .ZN(n488) );
  NAND2_X1 U601 ( .A1(n511), .A2(G210), .ZN(n487) );
  XNOR2_X1 U602 ( .A(n488), .B(n487), .ZN(n490) );
  XNOR2_X1 U603 ( .A(n490), .B(n489), .ZN(n491) );
  NAND2_X1 U604 ( .A1(n687), .A2(n528), .ZN(n493) );
  INV_X1 U605 ( .A(G472), .ZN(n492) );
  INV_X1 U606 ( .A(n704), .ZN(n494) );
  NOR2_X1 U607 ( .A1(n495), .A2(n494), .ZN(n496) );
  AND2_X1 U608 ( .A1(n497), .A2(n496), .ZN(n746) );
  XOR2_X1 U609 ( .A(n498), .B(G116), .Z(n499) );
  XNOR2_X1 U610 ( .A(n499), .B(KEYINPUT7), .ZN(n505) );
  INV_X1 U611 ( .A(KEYINPUT101), .ZN(n500) );
  XNOR2_X1 U612 ( .A(n501), .B(n500), .ZN(n503) );
  XNOR2_X1 U613 ( .A(G134), .B(KEYINPUT9), .ZN(n502) );
  XNOR2_X1 U614 ( .A(n503), .B(n502), .ZN(n504) );
  NAND2_X1 U615 ( .A1(n506), .A2(G217), .ZN(n507) );
  NAND2_X1 U616 ( .A1(n658), .A2(n528), .ZN(n510) );
  XNOR2_X1 U617 ( .A(KEYINPUT102), .B(G478), .ZN(n509) );
  XNOR2_X1 U618 ( .A(n510), .B(n509), .ZN(n585) );
  INV_X1 U619 ( .A(n585), .ZN(n531) );
  XOR2_X1 U620 ( .A(KEYINPUT100), .B(KEYINPUT98), .Z(n513) );
  NAND2_X1 U621 ( .A1(G214), .A2(n511), .ZN(n512) );
  XNOR2_X1 U622 ( .A(n513), .B(n512), .ZN(n517) );
  XOR2_X1 U623 ( .A(KEYINPUT12), .B(KEYINPUT99), .Z(n515) );
  XNOR2_X1 U624 ( .A(G140), .B(KEYINPUT11), .ZN(n514) );
  XNOR2_X1 U625 ( .A(n515), .B(n514), .ZN(n516) );
  XOR2_X1 U626 ( .A(n517), .B(n516), .Z(n522) );
  INV_X1 U627 ( .A(n518), .ZN(n520) );
  XNOR2_X1 U628 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U629 ( .A(n522), .B(n521), .ZN(n527) );
  INV_X1 U630 ( .A(n523), .ZN(n525) );
  XOR2_X1 U631 ( .A(n525), .B(n524), .Z(n526) );
  XNOR2_X1 U632 ( .A(n527), .B(n526), .ZN(n663) );
  NAND2_X1 U633 ( .A1(n663), .A2(n528), .ZN(n530) );
  XOR2_X1 U634 ( .A(KEYINPUT13), .B(G475), .Z(n529) );
  XNOR2_X1 U635 ( .A(n530), .B(n529), .ZN(n584) );
  AND2_X1 U636 ( .A1(n531), .A2(n584), .ZN(n756) );
  NAND2_X1 U637 ( .A1(n746), .A2(n756), .ZN(n532) );
  XNOR2_X1 U638 ( .A(n532), .B(G104), .ZN(G6) );
  XNOR2_X1 U639 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n533) );
  INV_X1 U640 ( .A(n558), .ZN(n573) );
  INV_X1 U641 ( .A(n573), .ZN(n697) );
  INV_X1 U642 ( .A(n756), .ZN(n542) );
  OR2_X1 U643 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U644 ( .A1(G900), .A2(n537), .ZN(n538) );
  NOR2_X1 U645 ( .A1(n539), .A2(n538), .ZN(n605) );
  NOR2_X1 U646 ( .A1(n605), .A2(n701), .ZN(n540) );
  XNOR2_X1 U647 ( .A(n540), .B(KEYINPUT74), .ZN(n612) );
  NAND2_X1 U648 ( .A1(n711), .A2(n612), .ZN(n541) );
  NOR2_X1 U649 ( .A1(n542), .A2(n541), .ZN(n546) );
  INV_X1 U650 ( .A(KEYINPUT6), .ZN(n544) );
  NOR2_X1 U651 ( .A1(n615), .A2(n572), .ZN(n545) );
  NAND2_X1 U652 ( .A1(n546), .A2(n545), .ZN(n624) );
  OR2_X1 U653 ( .A1(n697), .A2(n624), .ZN(n547) );
  XNOR2_X1 U654 ( .A(n547), .B(KEYINPUT43), .ZN(n549) );
  AND2_X1 U655 ( .A1(n549), .A2(n623), .ZN(n647) );
  XOR2_X1 U656 ( .A(n647), .B(G140), .Z(G42) );
  INV_X1 U657 ( .A(n714), .ZN(n551) );
  INV_X1 U658 ( .A(KEYINPUT22), .ZN(n553) );
  INV_X1 U659 ( .A(n571), .ZN(n557) );
  XNOR2_X1 U660 ( .A(n615), .B(KEYINPUT103), .ZN(n700) );
  INV_X1 U661 ( .A(n700), .ZN(n555) );
  NAND2_X1 U662 ( .A1(n555), .A2(n572), .ZN(n556) );
  OR2_X1 U663 ( .A1(n557), .A2(n556), .ZN(n589) );
  XNOR2_X1 U664 ( .A(n589), .B(G101), .ZN(G3) );
  XNOR2_X1 U665 ( .A(n560), .B(KEYINPUT33), .ZN(n719) );
  INV_X1 U666 ( .A(KEYINPUT78), .ZN(n562) );
  XNOR2_X1 U667 ( .A(n564), .B(n563), .ZN(n565) );
  AND2_X1 U668 ( .A1(n585), .A2(n584), .ZN(n620) );
  NAND2_X1 U669 ( .A1(n565), .A2(n620), .ZN(n567) );
  XNOR2_X1 U670 ( .A(KEYINPUT83), .B(KEYINPUT35), .ZN(n566) );
  XNOR2_X1 U671 ( .A(n567), .B(n566), .ZN(n597) );
  INV_X1 U672 ( .A(KEYINPUT104), .ZN(n568) );
  NOR2_X1 U673 ( .A1(n613), .A2(n615), .ZN(n570) );
  NAND2_X1 U674 ( .A1(n572), .A2(n700), .ZN(n574) );
  NOR2_X1 U675 ( .A1(n574), .A2(n573), .ZN(n575) );
  INV_X1 U676 ( .A(KEYINPUT84), .ZN(n576) );
  XNOR2_X1 U677 ( .A(n576), .B(KEYINPUT32), .ZN(n577) );
  NAND2_X1 U678 ( .A1(n597), .A2(n579), .ZN(n580) );
  NAND2_X1 U679 ( .A1(n580), .A2(KEYINPUT44), .ZN(n596) );
  NOR2_X1 U680 ( .A1(n581), .A2(n704), .ZN(n708) );
  NAND2_X1 U681 ( .A1(n708), .A2(n582), .ZN(n583) );
  XNOR2_X1 U682 ( .A(n583), .B(KEYINPUT31), .ZN(n759) );
  INV_X1 U683 ( .A(n584), .ZN(n586) );
  AND2_X1 U684 ( .A1(n586), .A2(n585), .ZN(n760) );
  OR2_X1 U685 ( .A1(n756), .A2(n760), .ZN(n633) );
  XNOR2_X1 U686 ( .A(n633), .B(KEYINPUT86), .ZN(n587) );
  NAND2_X1 U687 ( .A1(n588), .A2(n587), .ZN(n590) );
  NAND2_X1 U688 ( .A1(n590), .A2(n589), .ZN(n594) );
  INV_X1 U689 ( .A(KEYINPUT66), .ZN(n591) );
  NOR2_X1 U690 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U691 ( .A1(n598), .A2(KEYINPUT44), .ZN(n599) );
  NAND2_X1 U692 ( .A1(n737), .A2(n599), .ZN(n600) );
  INV_X1 U693 ( .A(KEYINPUT45), .ZN(n601) );
  NAND2_X1 U694 ( .A1(n711), .A2(n613), .ZN(n604) );
  NOR2_X1 U695 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U696 ( .A(n623), .B(KEYINPUT38), .ZN(n712) );
  INV_X1 U697 ( .A(n712), .ZN(n609) );
  NAND2_X1 U698 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U699 ( .A1(n712), .A2(n711), .ZN(n715) );
  NOR2_X1 U700 ( .A1(n715), .A2(n714), .ZN(n617) );
  XNOR2_X1 U701 ( .A(n617), .B(KEYINPUT41), .ZN(n729) );
  XOR2_X1 U702 ( .A(KEYINPUT42), .B(n618), .Z(n793) );
  NAND2_X1 U703 ( .A1(n422), .A2(n620), .ZN(n621) );
  NOR2_X1 U704 ( .A1(n622), .A2(n621), .ZN(n753) );
  NOR2_X1 U705 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U706 ( .A(n625), .B(KEYINPUT36), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n626), .A2(n697), .ZN(n763) );
  INV_X1 U708 ( .A(n627), .ZN(n629) );
  NAND2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n634) );
  INV_X1 U710 ( .A(n634), .ZN(n754) );
  NOR2_X1 U711 ( .A1(n633), .A2(KEYINPUT86), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n754), .A2(n630), .ZN(n631) );
  NAND2_X1 U713 ( .A1(n763), .A2(n631), .ZN(n632) );
  NOR2_X1 U714 ( .A1(n753), .A2(n632), .ZN(n641) );
  INV_X1 U715 ( .A(KEYINPUT47), .ZN(n636) );
  INV_X1 U716 ( .A(n633), .ZN(n716) );
  NOR2_X1 U717 ( .A1(n634), .A2(n716), .ZN(n637) );
  NAND2_X1 U718 ( .A1(n637), .A2(KEYINPUT86), .ZN(n635) );
  NAND2_X1 U719 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n637), .A2(KEYINPUT47), .ZN(n638) );
  NAND2_X1 U721 ( .A1(n639), .A2(n638), .ZN(n640) );
  AND2_X1 U722 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U723 ( .A(n643), .B(KEYINPUT48), .ZN(n649) );
  NAND2_X1 U724 ( .A1(n644), .A2(n760), .ZN(n646) );
  INV_X1 U725 ( .A(KEYINPUT106), .ZN(n645) );
  XNOR2_X1 U726 ( .A(n646), .B(n645), .ZN(n792) );
  NOR2_X1 U727 ( .A1(n792), .A2(n647), .ZN(n648) );
  NAND2_X1 U728 ( .A1(n649), .A2(n648), .ZN(n652) );
  INV_X1 U729 ( .A(KEYINPUT2), .ZN(n650) );
  INV_X1 U730 ( .A(n652), .ZN(n653) );
  NAND2_X1 U731 ( .A1(n653), .A2(KEYINPUT2), .ZN(n654) );
  XNOR2_X1 U732 ( .A(n654), .B(KEYINPUT88), .ZN(n657) );
  INV_X1 U733 ( .A(G952), .ZN(n659) );
  NAND2_X1 U734 ( .A1(n781), .A2(n659), .ZN(n660) );
  INV_X1 U735 ( .A(n690), .ZN(n744) );
  NOR2_X1 U736 ( .A1(n661), .A2(n744), .ZN(G63) );
  NAND2_X1 U737 ( .A1(n685), .A2(G475), .ZN(n665) );
  XNOR2_X1 U738 ( .A(KEYINPUT91), .B(KEYINPUT59), .ZN(n662) );
  XNOR2_X1 U739 ( .A(n665), .B(n664), .ZN(n666) );
  NAND2_X1 U740 ( .A1(n666), .A2(n690), .ZN(n668) );
  XNOR2_X1 U741 ( .A(KEYINPUT69), .B(KEYINPUT60), .ZN(n667) );
  XNOR2_X1 U742 ( .A(n668), .B(n667), .ZN(G60) );
  NAND2_X1 U743 ( .A1(n685), .A2(G210), .ZN(n673) );
  XNOR2_X1 U744 ( .A(KEYINPUT115), .B(KEYINPUT54), .ZN(n669) );
  XNOR2_X1 U745 ( .A(n669), .B(KEYINPUT55), .ZN(n670) );
  XNOR2_X1 U746 ( .A(n673), .B(n672), .ZN(n674) );
  NAND2_X1 U747 ( .A1(n674), .A2(n690), .ZN(n676) );
  XOR2_X1 U748 ( .A(KEYINPUT116), .B(KEYINPUT56), .Z(n675) );
  XNOR2_X1 U749 ( .A(n676), .B(n675), .ZN(G51) );
  XNOR2_X1 U750 ( .A(G119), .B(KEYINPUT126), .ZN(n678) );
  XOR2_X1 U751 ( .A(n678), .B(n677), .Z(G21) );
  NAND2_X1 U752 ( .A1(n685), .A2(G217), .ZN(n682) );
  XOR2_X1 U753 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n679) );
  XNOR2_X1 U754 ( .A(n682), .B(n681), .ZN(n683) );
  NAND2_X1 U755 ( .A1(n683), .A2(n690), .ZN(n684) );
  XNOR2_X1 U756 ( .A(n684), .B(KEYINPUT121), .ZN(G66) );
  NAND2_X1 U757 ( .A1(n685), .A2(G472), .ZN(n689) );
  XOR2_X1 U758 ( .A(KEYINPUT107), .B(KEYINPUT62), .Z(n686) );
  XNOR2_X1 U759 ( .A(n689), .B(n688), .ZN(n691) );
  NAND2_X1 U760 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U761 ( .A(n692), .B(KEYINPUT63), .ZN(G57) );
  NOR2_X1 U762 ( .A1(n656), .A2(n779), .ZN(n694) );
  XOR2_X1 U763 ( .A(KEYINPUT2), .B(KEYINPUT85), .Z(n693) );
  NOR2_X1 U764 ( .A1(n694), .A2(n693), .ZN(n696) );
  OR2_X1 U765 ( .A1(n696), .A2(n695), .ZN(n734) );
  XNOR2_X1 U766 ( .A(KEYINPUT50), .B(KEYINPUT110), .ZN(n698) );
  XNOR2_X1 U767 ( .A(n699), .B(n698), .ZN(n706) );
  NAND2_X1 U768 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U769 ( .A(KEYINPUT49), .B(n702), .Z(n703) );
  NAND2_X1 U770 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U771 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U772 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U773 ( .A(KEYINPUT51), .B(n709), .Z(n710) );
  NOR2_X1 U774 ( .A1(n729), .A2(n710), .ZN(n723) );
  NOR2_X1 U775 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U776 ( .A1(n714), .A2(n713), .ZN(n718) );
  NOR2_X1 U777 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U778 ( .A1(n718), .A2(n717), .ZN(n720) );
  BUF_X1 U779 ( .A(n719), .Z(n730) );
  NOR2_X1 U780 ( .A1(n720), .A2(n730), .ZN(n721) );
  XOR2_X1 U781 ( .A(KEYINPUT111), .B(n721), .Z(n722) );
  NOR2_X1 U782 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U783 ( .A(KEYINPUT112), .B(n724), .Z(n725) );
  XOR2_X1 U784 ( .A(KEYINPUT52), .B(n725), .Z(n727) );
  NOR2_X1 U785 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U786 ( .A(n728), .B(KEYINPUT113), .Z(n732) );
  NOR2_X1 U787 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U788 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U789 ( .A(n736), .B(n735), .ZN(G12) );
  XNOR2_X1 U790 ( .A(n737), .B(G122), .ZN(G24) );
  NAND2_X1 U791 ( .A1(n361), .A2(G469), .ZN(n743) );
  XOR2_X1 U792 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n739) );
  XNOR2_X1 U793 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n738) );
  XNOR2_X1 U794 ( .A(n739), .B(n738), .ZN(n740) );
  XNOR2_X1 U795 ( .A(n741), .B(n740), .ZN(n742) );
  XNOR2_X1 U796 ( .A(n743), .B(n742), .ZN(n745) );
  NOR2_X1 U797 ( .A1(n745), .A2(n744), .ZN(G54) );
  XNOR2_X1 U798 ( .A(G107), .B(KEYINPUT26), .ZN(n750) );
  NAND2_X1 U799 ( .A1(n746), .A2(n760), .ZN(n748) );
  XOR2_X1 U800 ( .A(KEYINPUT27), .B(KEYINPUT108), .Z(n747) );
  XNOR2_X1 U801 ( .A(n748), .B(n747), .ZN(n749) );
  XNOR2_X1 U802 ( .A(n750), .B(n749), .ZN(G9) );
  XOR2_X1 U803 ( .A(n359), .B(KEYINPUT29), .Z(n752) );
  NAND2_X1 U804 ( .A1(n754), .A2(n760), .ZN(n751) );
  XNOR2_X1 U805 ( .A(n752), .B(n751), .ZN(G30) );
  XOR2_X1 U806 ( .A(G143), .B(n753), .Z(G45) );
  NAND2_X1 U807 ( .A1(n754), .A2(n756), .ZN(n755) );
  XNOR2_X1 U808 ( .A(n755), .B(G146), .ZN(G48) );
  XOR2_X1 U809 ( .A(G113), .B(KEYINPUT109), .Z(n758) );
  NAND2_X1 U810 ( .A1(n756), .A2(n759), .ZN(n757) );
  XNOR2_X1 U811 ( .A(n758), .B(n757), .ZN(G15) );
  NAND2_X1 U812 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U813 ( .A(n761), .B(G116), .ZN(G18) );
  XOR2_X1 U814 ( .A(G125), .B(KEYINPUT37), .Z(n762) );
  XNOR2_X1 U815 ( .A(n763), .B(n762), .ZN(G27) );
  INV_X1 U816 ( .A(n656), .ZN(n765) );
  NAND2_X1 U817 ( .A1(n765), .A2(n764), .ZN(n769) );
  NAND2_X1 U818 ( .A1(G953), .A2(G224), .ZN(n766) );
  XNOR2_X1 U819 ( .A(KEYINPUT61), .B(n766), .ZN(n767) );
  NAND2_X1 U820 ( .A1(n767), .A2(G898), .ZN(n768) );
  NAND2_X1 U821 ( .A1(n769), .A2(n768), .ZN(n774) );
  XNOR2_X1 U822 ( .A(n770), .B(G101), .ZN(n772) );
  NAND2_X1 U823 ( .A1(n772), .A2(n771), .ZN(n773) );
  XOR2_X1 U824 ( .A(n774), .B(n773), .Z(G69) );
  XOR2_X1 U825 ( .A(KEYINPUT122), .B(n775), .Z(n778) );
  XNOR2_X1 U826 ( .A(n778), .B(n777), .ZN(n783) );
  XOR2_X1 U827 ( .A(n783), .B(n779), .Z(n780) );
  NOR2_X1 U828 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U829 ( .A(n782), .B(KEYINPUT123), .ZN(n789) );
  XNOR2_X1 U830 ( .A(n783), .B(G227), .ZN(n784) );
  XNOR2_X1 U831 ( .A(n784), .B(KEYINPUT124), .ZN(n785) );
  NAND2_X1 U832 ( .A1(n785), .A2(G900), .ZN(n786) );
  XOR2_X1 U833 ( .A(KEYINPUT125), .B(n786), .Z(n787) );
  NAND2_X1 U834 ( .A1(n787), .A2(G953), .ZN(n788) );
  NAND2_X1 U835 ( .A1(n789), .A2(n788), .ZN(G72) );
  XOR2_X1 U836 ( .A(G131), .B(n790), .Z(n791) );
  XNOR2_X1 U837 ( .A(KEYINPUT127), .B(n791), .ZN(G33) );
  XOR2_X1 U838 ( .A(G134), .B(n792), .Z(G36) );
  XNOR2_X1 U839 ( .A(G137), .B(n793), .ZN(G39) );
endmodule

