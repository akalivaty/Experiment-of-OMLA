//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 1 0 0 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931;
  INV_X1    g000(.A(KEYINPUT81), .ZN(new_n187));
  INV_X1    g001(.A(G469), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(KEYINPUT1), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n192), .A2(new_n194), .A3(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(KEYINPUT1), .A3(G146), .ZN(new_n198));
  XNOR2_X1  g012(.A(G143), .B(G146), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n197), .B(new_n198), .C1(G128), .C2(new_n199), .ZN(new_n200));
  OR2_X1    g014(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G104), .ZN(new_n203));
  AND2_X1   g017(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n201), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G101), .ZN(new_n206));
  INV_X1    g020(.A(G104), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G107), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(G107), .ZN(new_n209));
  NOR2_X1   g023(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n205), .A2(new_n206), .A3(new_n208), .A4(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n203), .A2(new_n208), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G101), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n200), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT76), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT10), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n208), .B1(new_n201), .B2(new_n203), .ZN(new_n219));
  NAND2_X1  g033(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n210), .B1(new_n209), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(G101), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(KEYINPUT4), .A3(new_n212), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n199), .A2(KEYINPUT0), .A3(G128), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT0), .B(G128), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n224), .B1(new_n199), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT4), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n228), .B(G101), .C1(new_n219), .C2(new_n221), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n223), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT10), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n215), .A2(new_n216), .A3(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n218), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT11), .ZN(new_n234));
  INV_X1    g048(.A(G134), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n234), .B1(new_n235), .B2(G137), .ZN(new_n236));
  INV_X1    g050(.A(G137), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(KEYINPUT11), .A3(G134), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT64), .ZN(new_n240));
  INV_X1    g054(.A(G131), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n235), .A2(G137), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n239), .A2(new_n240), .A3(new_n241), .A4(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n236), .A2(new_n238), .A3(new_n241), .A4(new_n242), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT64), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n236), .A2(new_n242), .A3(new_n238), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n241), .B1(new_n247), .B2(KEYINPUT65), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT65), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n236), .A2(new_n238), .A3(new_n249), .A4(new_n242), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n233), .A2(new_n252), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n243), .A2(new_n245), .B1(new_n248), .B2(new_n250), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n218), .A2(new_n254), .A3(new_n230), .A4(new_n232), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n253), .A2(KEYINPUT78), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT78), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n233), .A2(new_n257), .A3(new_n252), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(G110), .B(G140), .ZN(new_n260));
  INV_X1    g074(.A(G953), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n261), .A2(G227), .ZN(new_n262));
  XOR2_X1   g076(.A(new_n260), .B(new_n262), .Z(new_n263));
  NAND2_X1  g077(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n212), .A2(new_n214), .ZN(new_n265));
  INV_X1    g079(.A(new_n200), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n215), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n252), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT12), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(new_n254), .B2(KEYINPUT77), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n268), .A2(KEYINPUT77), .A3(new_n270), .A4(new_n252), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n272), .A2(new_n255), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n263), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n264), .A2(G469), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n256), .A2(new_n275), .A3(new_n258), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT80), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT80), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n256), .A2(new_n280), .A3(new_n275), .A4(new_n258), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n272), .A2(new_n255), .A3(new_n263), .A4(new_n273), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n283), .B(KEYINPUT79), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(G902), .B1(new_n282), .B2(new_n285), .ZN(new_n286));
  AOI211_X1 g100(.A(new_n190), .B(new_n277), .C1(new_n286), .C2(new_n188), .ZN(new_n287));
  INV_X1    g101(.A(G221), .ZN(new_n288));
  XOR2_X1   g102(.A(KEYINPUT9), .B(G234), .Z(new_n289));
  AOI21_X1  g103(.A(new_n288), .B1(new_n289), .B2(new_n189), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n187), .B1(new_n287), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n282), .A2(new_n285), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n292), .A2(new_n188), .A3(new_n189), .ZN(new_n293));
  INV_X1    g107(.A(new_n190), .ZN(new_n294));
  INV_X1    g108(.A(new_n277), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n290), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(KEYINPUT81), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n291), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(G472), .A2(G902), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT31), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n247), .A2(KEYINPUT65), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n302), .A2(G131), .A3(new_n250), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n244), .B(new_n240), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n227), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT66), .ZN(new_n306));
  INV_X1    g120(.A(new_n242), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n235), .A2(G137), .ZN(new_n308));
  OAI21_X1  g122(.A(G131), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n246), .A2(new_n306), .A3(new_n309), .A4(new_n200), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n200), .A2(new_n309), .ZN(new_n311));
  OAI21_X1  g125(.A(KEYINPUT66), .B1(new_n304), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n305), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT30), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(KEYINPUT2), .A2(G113), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT67), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT67), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(KEYINPUT2), .A3(G113), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT2), .ZN(new_n321));
  INV_X1    g135(.A(G113), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(G116), .B(G119), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n317), .A2(new_n319), .B1(new_n321), .B2(new_n322), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n325), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n244), .A2(KEYINPUT64), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n244), .A2(KEYINPUT64), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n309), .B(new_n200), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  OAI211_X1 g147(.A(KEYINPUT30), .B(new_n333), .C1(new_n254), .C2(new_n226), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n315), .A2(new_n330), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n327), .A2(new_n329), .A3(KEYINPUT68), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT68), .B1(new_n327), .B2(new_n329), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n305), .B(new_n333), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT26), .B(G101), .ZN(new_n340));
  INV_X1    g154(.A(G237), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(new_n261), .A3(G210), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n340), .B(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n343), .B(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n335), .A2(new_n339), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT70), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT70), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n335), .A2(new_n348), .A3(new_n339), .A4(new_n345), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n301), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT28), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n339), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n333), .B1(new_n254), .B2(new_n226), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n337), .A2(new_n338), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n355), .B1(new_n330), .B2(new_n313), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n352), .B1(new_n356), .B2(new_n351), .ZN(new_n357));
  INV_X1    g171(.A(new_n345), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n335), .A2(new_n301), .A3(new_n339), .A4(new_n345), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n300), .B1(new_n350), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT32), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n352), .B(new_n345), .C1(new_n356), .C2(new_n351), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n334), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n367), .B1(new_n314), .B2(new_n313), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n355), .B1(new_n368), .B2(new_n330), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(new_n345), .ZN(new_n370));
  NOR3_X1   g184(.A1(new_n366), .A2(new_n370), .A3(KEYINPUT29), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT71), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n353), .A2(new_n354), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n351), .B1(new_n339), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n352), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n345), .A2(KEYINPUT29), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n372), .B(new_n189), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n355), .A2(KEYINPUT28), .ZN(new_n379));
  NOR3_X1   g193(.A1(new_n374), .A2(new_n379), .A3(new_n377), .ZN(new_n380));
  OAI21_X1  g194(.A(KEYINPUT71), .B1(new_n380), .B2(G902), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(G472), .B1(new_n371), .B2(new_n382), .ZN(new_n383));
  OAI211_X1 g197(.A(KEYINPUT32), .B(new_n300), .C1(new_n350), .C2(new_n361), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n364), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G234), .ZN(new_n386));
  OAI21_X1  g200(.A(G217), .B1(new_n386), .B2(G902), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(G125), .B(G140), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT16), .ZN(new_n390));
  INV_X1    g204(.A(G125), .ZN(new_n391));
  OR3_X1    g205(.A1(new_n391), .A2(KEYINPUT16), .A3(G140), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n390), .A2(G146), .A3(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(KEYINPUT73), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n389), .A2(new_n193), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT24), .B(G110), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(KEYINPUT72), .ZN(new_n397));
  INV_X1    g211(.A(G119), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G128), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n191), .A2(G119), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT23), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n191), .A2(KEYINPUT23), .A3(G119), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(new_n399), .A3(new_n405), .ZN(new_n406));
  OAI22_X1  g220(.A1(new_n397), .A2(new_n402), .B1(G110), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n394), .A2(new_n395), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n397), .A2(new_n402), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n406), .A2(G110), .ZN(new_n410));
  AOI21_X1  g224(.A(G146), .B1(new_n390), .B2(new_n392), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n409), .B(new_n410), .C1(new_n411), .C2(new_n393), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n261), .A2(G221), .A3(G234), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(KEYINPUT22), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n415), .B(G137), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n408), .A2(new_n412), .A3(new_n416), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n189), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT25), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n420), .A2(new_n421), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n388), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT74), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI211_X1 g241(.A(KEYINPUT74), .B(new_n388), .C1(new_n423), .C2(new_n424), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n418), .A2(new_n419), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n388), .A2(G902), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n427), .A2(new_n428), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n385), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(G214), .B1(G237), .B2(G902), .ZN(new_n435));
  XOR2_X1   g249(.A(new_n435), .B(KEYINPUT82), .Z(new_n436));
  XOR2_X1   g250(.A(G110), .B(G122), .Z(new_n437));
  XOR2_X1   g251(.A(new_n437), .B(KEYINPUT8), .Z(new_n438));
  INV_X1    g252(.A(new_n265), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n325), .A2(KEYINPUT5), .ZN(new_n440));
  INV_X1    g254(.A(G116), .ZN(new_n441));
  OR3_X1    g255(.A1(new_n441), .A2(KEYINPUT5), .A3(G119), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n440), .A2(G113), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n329), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n439), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT84), .ZN(new_n446));
  OR2_X1    g260(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n443), .A2(new_n446), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(new_n329), .A3(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n438), .B(new_n445), .C1(new_n449), .C2(new_n439), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n223), .A2(new_n330), .A3(new_n229), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT83), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n447), .A2(new_n439), .A3(new_n329), .A4(new_n448), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT83), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n223), .A2(new_n330), .A3(new_n454), .A4(new_n229), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n452), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n450), .B1(new_n456), .B2(new_n437), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n226), .A2(G125), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n458), .B1(G125), .B2(new_n200), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n261), .A2(G224), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT7), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n459), .B(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n189), .B1(new_n457), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(KEYINPUT87), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT6), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT85), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n456), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n452), .A2(KEYINPUT85), .A3(new_n453), .A4(new_n455), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n437), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n465), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n470), .B1(new_n467), .B2(new_n468), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n456), .A2(new_n437), .ZN(new_n473));
  OAI21_X1  g287(.A(KEYINPUT6), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n459), .B(new_n460), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(KEYINPUT86), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT86), .ZN(new_n479));
  AOI211_X1 g293(.A(new_n479), .B(new_n476), .C1(new_n471), .C2(new_n474), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n464), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(G210), .B1(G237), .B2(G902), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n482), .B(new_n464), .C1(new_n478), .C2(new_n480), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n436), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OR3_X1    g300(.A1(new_n393), .A2(new_n411), .A3(KEYINPUT92), .ZN(new_n487));
  OAI21_X1  g301(.A(KEYINPUT92), .B1(new_n393), .B2(new_n411), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n341), .A2(new_n261), .A3(G214), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(G143), .ZN(new_n491));
  OR2_X1    g305(.A1(new_n491), .A2(new_n241), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT17), .ZN(new_n493));
  OR2_X1    g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n491), .A2(new_n241), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(KEYINPUT89), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT89), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n491), .A2(new_n497), .A3(new_n241), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n496), .A2(new_n492), .A3(new_n498), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n489), .B(new_n494), .C1(KEYINPUT17), .C2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(KEYINPUT18), .A2(G131), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n491), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n502), .B(KEYINPUT88), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n389), .B(new_n193), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n503), .B(new_n504), .C1(new_n491), .C2(new_n501), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(G113), .B(G122), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT91), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n507), .B(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(KEYINPUT90), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(new_n207), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT93), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n189), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n506), .A2(new_n512), .ZN(new_n515));
  OAI21_X1  g329(.A(G475), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  XOR2_X1   g330(.A(new_n389), .B(KEYINPUT19), .Z(new_n517));
  OAI211_X1 g331(.A(new_n394), .B(new_n499), .C1(G146), .C2(new_n517), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n511), .A2(new_n505), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n511), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n519), .B1(new_n520), .B2(new_n506), .ZN(new_n521));
  INV_X1    g335(.A(G475), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n521), .A2(KEYINPUT20), .A3(new_n522), .A4(new_n189), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n506), .A2(new_n520), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n511), .A2(new_n505), .A3(new_n518), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n524), .A2(new_n522), .A3(new_n189), .A4(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT20), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n516), .A2(new_n523), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n195), .A2(G128), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT13), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n191), .A2(G143), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n530), .A2(new_n531), .ZN(new_n535));
  OAI21_X1  g349(.A(G134), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n530), .A2(new_n533), .A3(new_n235), .ZN(new_n537));
  XNOR2_X1  g351(.A(G116), .B(G122), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(new_n202), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n538), .A2(new_n202), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n536), .B(new_n537), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT14), .B1(new_n441), .B2(G122), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n538), .B1(KEYINPUT14), .B2(new_n202), .ZN(new_n544));
  INV_X1    g358(.A(new_n537), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n235), .B1(new_n530), .B2(new_n533), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n543), .B(new_n544), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n541), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n289), .A2(G217), .A3(new_n261), .ZN(new_n549));
  OR2_X1    g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n549), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n550), .A2(KEYINPUT94), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT94), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n548), .A2(new_n553), .A3(new_n549), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n189), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(G478), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(KEYINPUT15), .ZN(new_n557));
  OR2_X1    g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n555), .A2(new_n557), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT95), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n558), .A2(KEYINPUT95), .A3(new_n559), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n261), .A2(G952), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n565), .B1(G234), .B2(G237), .ZN(new_n566));
  XOR2_X1   g380(.A(KEYINPUT21), .B(G898), .Z(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  OAI211_X1 g382(.A(G902), .B(G953), .C1(new_n386), .C2(new_n341), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n566), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n529), .A2(new_n564), .A3(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n299), .A2(new_n434), .A3(new_n486), .A4(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(G101), .ZN(G3));
  OAI21_X1  g388(.A(new_n189), .B1(new_n350), .B2(new_n361), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(G472), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n362), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n577), .B1(new_n291), .B2(new_n298), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n433), .ZN(new_n579));
  INV_X1    g393(.A(new_n486), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n555), .A2(new_n556), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT33), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n552), .A2(new_n582), .A3(new_n554), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n550), .A2(KEYINPUT33), .A3(new_n551), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n189), .A2(G478), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n581), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n529), .A2(new_n587), .ZN(new_n588));
  NOR4_X1   g402(.A1(new_n579), .A2(new_n580), .A3(new_n571), .A4(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT34), .B(G104), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(G6));
  INV_X1    g405(.A(new_n571), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n523), .A2(new_n516), .A3(new_n528), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n486), .A2(new_n592), .A3(new_n564), .A4(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n579), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g409(.A(KEYINPUT97), .B(G107), .Z(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT96), .B(KEYINPUT35), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(G9));
  AND2_X1   g413(.A1(new_n576), .A2(new_n362), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT99), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n417), .A2(KEYINPUT36), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(KEYINPUT98), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(new_n413), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n430), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n427), .A2(new_n428), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n600), .A2(new_n601), .A3(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n299), .A2(new_n486), .A3(new_n572), .A4(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n601), .B1(new_n600), .B2(new_n606), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(KEYINPUT100), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT37), .B(G110), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G12));
  INV_X1    g427(.A(KEYINPUT101), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n385), .A2(new_n606), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n296), .A2(KEYINPUT81), .A3(new_n297), .ZN(new_n616));
  AOI21_X1  g430(.A(KEYINPUT81), .B1(new_n296), .B2(new_n297), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n436), .ZN(new_n619));
  INV_X1    g433(.A(G900), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n566), .B1(new_n570), .B2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n593), .A2(new_n564), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n476), .B1(new_n471), .B2(new_n474), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT86), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n482), .B1(new_n626), .B2(new_n464), .ZN(new_n627));
  INV_X1    g441(.A(new_n485), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n619), .B(new_n624), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n614), .B1(new_n618), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n385), .A2(new_n606), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n631), .B1(new_n291), .B2(new_n298), .ZN(new_n632));
  AOI211_X1 g446(.A(new_n436), .B(new_n623), .C1(new_n484), .C2(new_n485), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(new_n633), .A3(KEYINPUT101), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G128), .ZN(G30));
  NAND2_X1  g450(.A1(new_n484), .A2(new_n485), .ZN(new_n637));
  XOR2_X1   g451(.A(new_n637), .B(KEYINPUT38), .Z(new_n638));
  AND2_X1   g452(.A1(new_n364), .A2(new_n384), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n347), .A2(new_n349), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n339), .A2(new_n373), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n641), .B1(new_n642), .B2(new_n358), .ZN(new_n643));
  OAI21_X1  g457(.A(G472), .B1(new_n643), .B2(G902), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n639), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n529), .A2(new_n564), .ZN(new_n647));
  NOR4_X1   g461(.A1(new_n638), .A2(new_n646), .A3(new_n436), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n621), .B(KEYINPUT39), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n299), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n606), .B1(new_n651), .B2(KEYINPUT40), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n648), .B(new_n652), .C1(KEYINPUT40), .C2(new_n651), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G143), .ZN(G45));
  NOR2_X1   g468(.A1(new_n588), .A2(new_n621), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n619), .B(new_n655), .C1(new_n627), .C2(new_n628), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT102), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n486), .A2(KEYINPUT102), .A3(new_n655), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n658), .A2(new_n632), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G146), .ZN(G48));
  AOI21_X1  g475(.A(new_n284), .B1(new_n279), .B2(new_n281), .ZN(new_n662));
  OAI21_X1  g476(.A(G469), .B1(new_n662), .B2(G902), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n293), .A2(new_n663), .A3(new_n297), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n664), .A2(new_n385), .A3(new_n433), .ZN(new_n665));
  INV_X1    g479(.A(new_n588), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n665), .A2(new_n486), .A3(new_n592), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT41), .B(G113), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G15));
  AND4_X1   g483(.A1(new_n619), .A2(new_n637), .A3(new_n592), .A4(new_n564), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n670), .A2(KEYINPUT103), .A3(new_n593), .A4(new_n665), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT103), .ZN(new_n672));
  INV_X1    g486(.A(new_n665), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n672), .B1(new_n594), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n675), .B(KEYINPUT104), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(new_n441), .ZN(G18));
  NAND4_X1  g491(.A1(new_n486), .A2(new_n615), .A3(new_n572), .A4(new_n664), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT105), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(new_n398), .ZN(G21));
  AOI211_X1 g494(.A(new_n436), .B(new_n571), .C1(new_n484), .C2(new_n485), .ZN(new_n681));
  INV_X1    g495(.A(new_n664), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n647), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT108), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n348), .B1(new_n369), .B2(new_n345), .ZN(new_n685));
  INV_X1    g499(.A(new_n349), .ZN(new_n686));
  OAI21_X1  g500(.A(KEYINPUT31), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n375), .A2(KEYINPUT106), .A3(new_n352), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n689), .B1(new_n374), .B2(new_n379), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n688), .A2(new_n690), .A3(new_n358), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n687), .A2(KEYINPUT107), .A3(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT107), .ZN(new_n693));
  AND3_X1   g507(.A1(new_n688), .A2(new_n690), .A3(new_n358), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n693), .B1(new_n350), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n692), .A2(new_n360), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n300), .ZN(new_n697));
  AND4_X1   g511(.A1(new_n684), .A2(new_n697), .A3(new_n433), .A4(new_n576), .ZN(new_n698));
  AOI22_X1  g512(.A1(new_n696), .A2(new_n300), .B1(G472), .B2(new_n575), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n684), .B1(new_n699), .B2(new_n433), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n681), .B(new_n683), .C1(new_n698), .C2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT109), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n697), .A2(new_n576), .ZN(new_n703));
  OAI21_X1  g517(.A(KEYINPUT108), .B1(new_n703), .B2(new_n432), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n699), .A2(new_n684), .A3(new_n433), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT109), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n706), .A2(new_n707), .A3(new_n681), .A4(new_n683), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n702), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G122), .ZN(G24));
  AND2_X1   g524(.A1(new_n699), .A2(new_n606), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n711), .A2(new_n486), .A3(new_n655), .A4(new_n664), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G125), .ZN(G27));
  OR2_X1    g527(.A1(new_n276), .A2(KEYINPUT110), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n276), .A2(KEYINPUT110), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n714), .A2(new_n264), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(G469), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n293), .A2(new_n294), .A3(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n718), .A2(new_n719), .A3(new_n297), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n719), .B1(new_n718), .B2(new_n297), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n637), .A2(new_n436), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n722), .A2(new_n723), .A3(new_n434), .A4(new_n655), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT42), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR4_X1   g540(.A1(new_n637), .A2(new_n436), .A3(new_n588), .A4(new_n621), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n727), .A2(KEYINPUT42), .A3(new_n434), .A4(new_n722), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G131), .ZN(G33));
  NAND2_X1  g544(.A1(new_n723), .A2(new_n624), .ZN(new_n731));
  INV_X1    g545(.A(new_n721), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n718), .A2(new_n719), .A3(new_n297), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n732), .A2(new_n434), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(KEYINPUT112), .B1(new_n731), .B2(new_n734), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n637), .A2(new_n436), .A3(new_n623), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT112), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n736), .A2(new_n737), .A3(new_n434), .A4(new_n722), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G134), .ZN(G36));
  AOI21_X1  g554(.A(new_n188), .B1(new_n716), .B2(KEYINPUT45), .ZN(new_n741));
  INV_X1    g555(.A(new_n276), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n742), .B1(new_n259), .B2(new_n263), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n741), .B1(KEYINPUT45), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT46), .B1(new_n744), .B2(new_n294), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n293), .B1(new_n745), .B2(KEYINPUT113), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n746), .B1(KEYINPUT113), .B2(new_n745), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n744), .A2(KEYINPUT46), .A3(new_n294), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n290), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n650), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n593), .A2(new_n587), .ZN(new_n752));
  XOR2_X1   g566(.A(new_n752), .B(KEYINPUT43), .Z(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n577), .A3(new_n606), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n750), .B1(new_n751), .B2(new_n754), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n755), .B(new_n723), .C1(new_n751), .C2(new_n754), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G137), .ZN(G39));
  INV_X1    g571(.A(KEYINPUT47), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n749), .A2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n749), .A2(new_n758), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n385), .A2(new_n433), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n727), .A3(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G140), .ZN(G42));
  NOR3_X1   g579(.A1(new_n637), .A2(new_n682), .A3(new_n436), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n766), .A2(new_n433), .A3(new_n566), .A4(new_n646), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n767), .A2(new_n529), .A3(new_n587), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n706), .A2(new_n566), .A3(new_n753), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n682), .A2(new_n619), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n770), .A2(KEYINPUT118), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(KEYINPUT118), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n769), .A2(new_n638), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT50), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n766), .A2(new_n566), .A3(new_n753), .ZN(new_n775));
  AOI211_X1 g589(.A(new_n768), .B(new_n774), .C1(new_n711), .C2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n293), .A2(new_n663), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n290), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n779), .B1(new_n760), .B2(new_n761), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n769), .A2(new_n723), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n776), .A2(KEYINPUT51), .A3(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n767), .A2(new_n588), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n580), .A2(new_n682), .ZN(new_n785));
  AOI211_X1 g599(.A(new_n565), .B(new_n784), .C1(new_n785), .C2(new_n769), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT117), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n762), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n779), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n762), .A2(new_n788), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n781), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT51), .B1(new_n776), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n787), .A2(new_n793), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n618), .A2(new_n614), .A3(new_n629), .ZN(new_n795));
  AOI21_X1  g609(.A(KEYINPUT101), .B1(new_n632), .B2(new_n633), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n660), .B(new_n712), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n606), .A2(new_n621), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n645), .A2(new_n297), .A3(new_n718), .A4(new_n798), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n799), .A2(new_n580), .A3(new_n647), .ZN(new_n800));
  OAI21_X1  g614(.A(KEYINPUT115), .B1(new_n797), .B2(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n660), .A2(new_n712), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n803));
  INV_X1    g617(.A(new_n800), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n802), .A2(new_n803), .A3(new_n635), .A4(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n801), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n560), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n588), .B1(new_n808), .B2(new_n529), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n578), .A2(new_n681), .A3(new_n433), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n573), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(new_n610), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n667), .A2(new_n678), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n813), .B1(new_n671), .B2(new_n674), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n812), .A2(new_n814), .A3(new_n709), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n529), .A2(new_n621), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n632), .A2(new_n808), .A3(new_n723), .A4(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n727), .A2(new_n711), .A3(new_n722), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n729), .A2(new_n739), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(KEYINPUT52), .B1(new_n797), .B2(new_n800), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n807), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n822), .A2(KEYINPUT53), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n801), .A2(new_n805), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(KEYINPUT52), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(new_n807), .A3(new_n820), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT53), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(KEYINPUT54), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n822), .A2(KEYINPUT53), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n825), .A2(new_n832), .A3(new_n807), .A4(new_n820), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n836), .A2(KEYINPUT116), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(KEYINPUT116), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n794), .A2(new_n830), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n775), .A2(new_n434), .ZN(new_n840));
  XOR2_X1   g654(.A(new_n840), .B(KEYINPUT48), .Z(new_n841));
  OAI22_X1  g655(.A1(new_n839), .A2(new_n841), .B1(G952), .B2(G953), .ZN(new_n842));
  AOI211_X1 g656(.A(new_n290), .B(new_n432), .C1(KEYINPUT49), .C2(new_n777), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n843), .A2(new_n619), .A3(new_n593), .A4(new_n587), .ZN(new_n844));
  XOR2_X1   g658(.A(new_n844), .B(KEYINPUT114), .Z(new_n845));
  INV_X1    g659(.A(KEYINPUT49), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n645), .B1(new_n846), .B2(new_n778), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n845), .A2(new_n638), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n842), .A2(new_n848), .ZN(G75));
  NOR2_X1   g663(.A1(new_n834), .A2(new_n189), .ZN(new_n850));
  AOI21_X1  g664(.A(KEYINPUT56), .B1(new_n850), .B2(G210), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n475), .A2(new_n477), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n852), .A2(new_n625), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(KEYINPUT55), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n851), .B(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n261), .A2(G952), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(G51));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n831), .A2(new_n833), .A3(KEYINPUT54), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT119), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n831), .A2(new_n833), .A3(new_n861), .A4(KEYINPUT54), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n860), .A2(new_n836), .A3(new_n862), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n190), .B(KEYINPUT57), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n858), .B1(new_n865), .B2(new_n292), .ZN(new_n866));
  AOI211_X1 g680(.A(KEYINPUT120), .B(new_n662), .C1(new_n863), .C2(new_n864), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OR3_X1    g682(.A1(new_n834), .A2(new_n189), .A3(new_n744), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n856), .B1(new_n868), .B2(new_n869), .ZN(G54));
  NAND3_X1  g684(.A1(new_n850), .A2(KEYINPUT58), .A3(G475), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(new_n521), .Z(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(new_n856), .ZN(G60));
  INV_X1    g687(.A(new_n585), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n837), .A2(new_n830), .A3(new_n838), .ZN(new_n875));
  NAND2_X1  g689(.A1(G478), .A2(G902), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT59), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n874), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n863), .A2(new_n874), .A3(new_n877), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n878), .A2(new_n856), .A3(new_n879), .ZN(G63));
  NAND2_X1  g694(.A1(G217), .A2(G902), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT60), .Z(new_n882));
  NAND3_X1  g696(.A1(new_n831), .A2(new_n833), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n429), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n856), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n831), .A2(new_n833), .A3(new_n604), .A4(new_n882), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT121), .ZN(new_n887));
  AOI22_X1  g701(.A1(new_n885), .A2(new_n886), .B1(new_n887), .B2(KEYINPUT61), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n887), .A2(KEYINPUT61), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n888), .B(new_n889), .ZN(G66));
  AOI21_X1  g704(.A(new_n261), .B1(new_n567), .B2(G224), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n891), .B1(new_n815), .B2(new_n261), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n471), .B(new_n474), .C1(G898), .C2(new_n261), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n892), .B(new_n893), .Z(G69));
  AOI21_X1  g708(.A(new_n261), .B1(G227), .B2(G900), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n895), .A2(KEYINPUT125), .ZN(new_n896));
  INV_X1    g710(.A(new_n895), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT125), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n368), .B(new_n517), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n261), .A2(G900), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(KEYINPUT123), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n756), .A2(new_n764), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n580), .A2(new_n647), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n749), .A2(new_n434), .A3(new_n650), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n729), .A2(new_n739), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT124), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n797), .B(KEYINPUT122), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n905), .A2(new_n907), .A3(new_n909), .A4(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n904), .B1(new_n911), .B2(new_n261), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n901), .B(new_n903), .C1(new_n912), .C2(new_n902), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n910), .A2(new_n653), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT62), .Z(new_n915));
  INV_X1    g729(.A(new_n651), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n916), .A2(new_n434), .A3(new_n723), .A4(new_n809), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n915), .A2(new_n905), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n918), .A2(new_n261), .A3(new_n900), .ZN(new_n919));
  AOI211_X1 g733(.A(new_n896), .B(new_n899), .C1(new_n913), .C2(new_n919), .ZN(new_n920));
  AND4_X1   g734(.A1(new_n898), .A2(new_n913), .A3(new_n897), .A4(new_n919), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(G72));
  NAND2_X1  g736(.A1(G472), .A2(G902), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT63), .Z(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT126), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(new_n911), .B2(new_n815), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n926), .A2(new_n358), .A3(new_n369), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n829), .B(new_n924), .C1(new_n370), .C2(new_n641), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n927), .B(new_n928), .C1(G952), .C2(new_n261), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n918), .A2(new_n815), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n369), .B1(new_n930), .B2(new_n925), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n929), .B1(new_n931), .B2(new_n345), .ZN(G57));
endmodule


