//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 1 0 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 1 1 1 0 0 0 1 0 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n569, new_n571, new_n572, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  XNOR2_X1  g032(.A(G325), .B(KEYINPUT67), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n460), .A2(G137), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n468), .A3(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n461), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n464), .A2(new_n471), .ZN(G160));
  NAND2_X1  g047(.A1(new_n466), .A2(new_n468), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G136), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n473), .A2(new_n461), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  NAND4_X1  g056(.A1(new_n466), .A2(new_n468), .A3(G138), .A4(new_n461), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n460), .A2(KEYINPUT4), .A3(G138), .A4(new_n461), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n489));
  OAI21_X1  g064(.A(G2105), .B1(new_n489), .B2(G114), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(KEYINPUT68), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n488), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n466), .A2(new_n468), .A3(G126), .A4(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT69), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n493), .A2(new_n497), .A3(new_n494), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n486), .B1(new_n496), .B2(new_n498), .ZN(G164));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT70), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT70), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  OR2_X1    g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g082(.A1(new_n507), .A2(G62), .ZN(new_n508));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  XOR2_X1   g084(.A(new_n509), .B(KEYINPUT72), .Z(new_n510));
  OAI21_X1  g085(.A(new_n504), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n512), .B1(new_n501), .B2(new_n503), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  OAI211_X1 g089(.A(G88), .B(new_n507), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  OAI211_X1 g090(.A(G50), .B(G543), .C1(new_n513), .C2(new_n514), .ZN(new_n516));
  AND3_X1   g091(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT71), .ZN(new_n517));
  AOI21_X1  g092(.A(KEYINPUT71), .B1(new_n515), .B2(new_n516), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n511), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(KEYINPUT73), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n515), .A2(new_n516), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT71), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n525), .A2(new_n526), .A3(new_n511), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n520), .A2(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XOR2_X1   g105(.A(new_n530), .B(KEYINPUT7), .Z(new_n531));
  AOI21_X1  g106(.A(new_n514), .B1(new_n504), .B2(KEYINPUT6), .ZN(new_n532));
  INV_X1    g107(.A(new_n507), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n531), .B1(new_n534), .B2(G89), .ZN(new_n535));
  OAI211_X1 g110(.A(G51), .B(G543), .C1(new_n513), .C2(new_n514), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n537));
  AND3_X1   g112(.A1(new_n536), .A2(KEYINPUT74), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g113(.A(KEYINPUT74), .B1(new_n536), .B2(new_n537), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n535), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g117(.A(new_n535), .B(KEYINPUT75), .C1(new_n538), .C2(new_n539), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(G168));
  INV_X1    g119(.A(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n532), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G52), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n534), .A2(G90), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  XNOR2_X1  g124(.A(KEYINPUT70), .B(G651), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n547), .A2(new_n548), .A3(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  INV_X1    g128(.A(new_n514), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n554), .B1(new_n550), .B2(new_n512), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n555), .A2(G43), .A3(G543), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n555), .A2(G81), .A3(new_n507), .ZN(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n558), .B1(new_n505), .B2(new_n506), .ZN(new_n559));
  AND2_X1   g134(.A1(G68), .A2(G543), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n504), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n556), .A2(new_n557), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT76), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT76), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n556), .A2(new_n557), .A3(new_n564), .A4(new_n561), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  AND3_X1   g143(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G36), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n569), .A2(new_n572), .ZN(G188));
  NAND3_X1  g148(.A1(new_n555), .A2(G53), .A3(G543), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(KEYINPUT9), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n555), .A2(new_n576), .A3(G53), .A4(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(KEYINPUT77), .B1(new_n532), .B2(new_n533), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT77), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n555), .A2(new_n580), .A3(new_n507), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(G91), .A3(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n507), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n583), .A2(new_n500), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n578), .A2(new_n582), .A3(new_n584), .ZN(G299));
  INV_X1    g160(.A(G168), .ZN(G286));
  NAND3_X1  g161(.A1(new_n579), .A2(G87), .A3(new_n581), .ZN(new_n587));
  INV_X1    g162(.A(G74), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n500), .B1(new_n533), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(new_n546), .B2(G49), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n587), .A2(new_n590), .ZN(G288));
  NAND2_X1  g166(.A1(new_n507), .A2(G61), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n550), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AND2_X1   g169(.A1(G48), .A2(G543), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n594), .B1(new_n555), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n579), .A2(G86), .A3(new_n581), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(G305));
  XNOR2_X1  g173(.A(KEYINPUT78), .B(G85), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n534), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n546), .A2(G47), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n602), .A2(new_n550), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(G290));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NOR2_X1   g180(.A1(G301), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n579), .A2(G92), .A3(new_n581), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n579), .A2(KEYINPUT10), .A3(new_n581), .A4(G92), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n533), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n546), .A2(G54), .B1(new_n614), .B2(G651), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT79), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n611), .A2(KEYINPUT79), .A3(new_n615), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n606), .B1(new_n620), .B2(new_n605), .ZN(G321));
  XNOR2_X1  g196(.A(G321), .B(KEYINPUT80), .ZN(G284));
  XNOR2_X1  g197(.A(G299), .B(KEYINPUT81), .ZN(new_n623));
  MUX2_X1   g198(.A(G286), .B(new_n623), .S(new_n605), .Z(G297));
  XNOR2_X1  g199(.A(G297), .B(KEYINPUT82), .ZN(G280));
  XOR2_X1   g200(.A(KEYINPUT83), .B(G559), .Z(new_n626));
  OAI21_X1  g201(.A(new_n620), .B1(G860), .B2(new_n626), .ZN(G148));
  INV_X1    g202(.A(KEYINPUT84), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n605), .B1(new_n620), .B2(new_n626), .ZN(new_n629));
  AOI211_X1 g204(.A(new_n628), .B(new_n629), .C1(new_n605), .C2(new_n566), .ZN(new_n630));
  AND2_X1   g205(.A1(new_n629), .A2(new_n628), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT11), .Z(G282));
  INV_X1    g208(.A(new_n632), .ZN(G323));
  NAND2_X1  g209(.A1(new_n474), .A2(G135), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n476), .A2(G123), .ZN(new_n636));
  OR2_X1    g211(.A1(G99), .A2(G2105), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n637), .B(G2104), .C1(G111), .C2(new_n461), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n635), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT85), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2096), .ZN(new_n641));
  INV_X1    g216(.A(KEYINPUT12), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n474), .A2(new_n642), .A3(G2104), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n460), .A2(new_n461), .ZN(new_n644));
  OAI21_X1  g219(.A(KEYINPUT12), .B1(new_n644), .B2(new_n465), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT13), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2100), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n641), .A2(new_n648), .ZN(G156));
  INV_X1    g224(.A(KEYINPUT14), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n650), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n653), .B2(new_n652), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n655), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  AND3_X1   g238(.A1(new_n662), .A2(G14), .A3(new_n663), .ZN(G401));
  XNOR2_X1  g239(.A(G2072), .B(G2078), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT17), .Z(new_n666));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT86), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n666), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT87), .Z(new_n672));
  NAND3_X1  g247(.A1(new_n668), .A2(new_n665), .A3(new_n669), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT18), .Z(new_n674));
  NOR2_X1   g249(.A1(new_n666), .A2(new_n670), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n665), .A2(new_n669), .ZN(new_n676));
  OR3_X1    g251(.A1(new_n675), .A2(new_n668), .A3(new_n676), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n672), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2096), .B(G2100), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT88), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(new_n680), .ZN(G227));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1956), .B(G2474), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT89), .ZN(new_n686));
  XOR2_X1   g261(.A(G1961), .B(G1966), .Z(new_n687));
  NAND3_X1  g262(.A1(new_n684), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT20), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n684), .B1(new_n686), .B2(new_n687), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n686), .A2(new_n687), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n689), .B(new_n692), .C1(new_n683), .C2(new_n691), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT90), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n693), .B(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(G1991), .B(G1996), .Z(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n696), .A2(new_n698), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1981), .B(G1986), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n699), .A2(new_n702), .A3(new_n700), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(G229));
  NAND2_X1  g281(.A1(new_n474), .A2(G139), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT25), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(G115), .A2(G2104), .ZN(new_n712));
  INV_X1    g287(.A(G127), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n473), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G2105), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n711), .B1(KEYINPUT95), .B2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT95), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n714), .A2(new_n717), .A3(G2105), .ZN(new_n718));
  AOI21_X1  g293(.A(KEYINPUT96), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n715), .A2(KEYINPUT95), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n720), .A2(new_n718), .A3(new_n710), .A4(new_n707), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT96), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(G29), .B1(new_n719), .B2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G33), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(G29), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(new_n442), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n728), .A2(G32), .ZN(new_n729));
  NAND3_X1  g304(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT99), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT98), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT26), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n732), .A2(KEYINPUT98), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n732), .A2(KEYINPUT98), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n736), .A2(KEYINPUT26), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n476), .A2(G129), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n474), .A2(G141), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n735), .A2(new_n738), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n729), .B1(new_n744), .B2(G29), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT27), .B(G1996), .ZN(new_n746));
  AND2_X1   g321(.A1(KEYINPUT24), .A2(G34), .ZN(new_n747));
  NOR2_X1   g322(.A1(KEYINPUT24), .A2(G34), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n728), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT97), .Z(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G29), .B2(G160), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n745), .A2(new_n746), .B1(G2084), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n727), .A2(new_n752), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT100), .Z(new_n754));
  NOR2_X1   g329(.A1(G4), .A2(G16), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n620), .B2(G16), .ZN(new_n756));
  INV_X1    g331(.A(G1348), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n728), .A2(G35), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT103), .Z(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G162), .B2(new_n728), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT29), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G2090), .ZN(new_n763));
  INV_X1    g338(.A(G16), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(G20), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT23), .Z(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G299), .B2(G16), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1956), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n764), .A2(G5), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G171), .B2(new_n764), .ZN(new_n770));
  INV_X1    g345(.A(G1961), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n745), .A2(new_n746), .ZN(new_n773));
  NAND4_X1  g348(.A1(new_n763), .A2(new_n768), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT31), .B(G11), .Z(new_n775));
  INV_X1    g350(.A(G28), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n776), .A2(KEYINPUT30), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT101), .Z(new_n778));
  AOI21_X1  g353(.A(G29), .B1(new_n776), .B2(KEYINPUT30), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n775), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n751), .A2(G2084), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT102), .ZN(new_n782));
  OAI221_X1 g357(.A(new_n780), .B1(new_n728), .B2(new_n639), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n728), .A2(G26), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT94), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT28), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n476), .A2(G128), .ZN(new_n787));
  INV_X1    g362(.A(G140), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(new_n644), .ZN(new_n789));
  OR2_X1    g364(.A1(G104), .A2(G2105), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n790), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT93), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n786), .B1(new_n793), .B2(new_n728), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G2067), .ZN(new_n795));
  AOI211_X1 g370(.A(new_n783), .B(new_n795), .C1(new_n782), .C2(new_n781), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n567), .A2(new_n764), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n764), .B2(G19), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(G1341), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n728), .A2(G27), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G164), .B2(new_n728), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(new_n443), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n796), .A2(new_n800), .A3(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n799), .A2(G1341), .ZN(new_n805));
  NOR3_X1   g380(.A1(new_n774), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n764), .A2(G21), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G168), .B2(new_n764), .ZN(new_n808));
  INV_X1    g383(.A(G1966), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n754), .A2(new_n758), .A3(new_n806), .A4(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(G290), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(G16), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G16), .B2(G24), .ZN(new_n814));
  INV_X1    g389(.A(G1986), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n814), .A2(new_n815), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n728), .A2(G25), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n474), .A2(G131), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n476), .A2(G119), .ZN(new_n821));
  OR2_X1    g396(.A1(G95), .A2(G2105), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n822), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n820), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n819), .B1(new_n825), .B2(new_n728), .ZN(new_n826));
  XOR2_X1   g401(.A(KEYINPUT35), .B(G1991), .Z(new_n827));
  XOR2_X1   g402(.A(new_n826), .B(new_n827), .Z(new_n828));
  NOR3_X1   g403(.A1(new_n817), .A2(new_n818), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(G16), .A2(G23), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT91), .ZN(new_n831));
  AND3_X1   g406(.A1(new_n587), .A2(new_n590), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n831), .B1(new_n587), .B2(new_n590), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n830), .B1(new_n834), .B2(G16), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT33), .B(G1976), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(G303), .A2(G16), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n764), .A2(G22), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT92), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n837), .B1(G1971), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n841), .A2(G1971), .ZN(new_n843));
  MUX2_X1   g418(.A(G6), .B(G305), .S(G16), .Z(new_n844));
  XOR2_X1   g419(.A(KEYINPUT32), .B(G1981), .Z(new_n845));
  XOR2_X1   g420(.A(new_n844), .B(new_n845), .Z(new_n846));
  NOR2_X1   g421(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n842), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n829), .B1(new_n848), .B2(KEYINPUT34), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT34), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(new_n842), .B2(new_n847), .ZN(new_n851));
  NOR3_X1   g426(.A1(new_n849), .A2(KEYINPUT36), .A3(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(KEYINPUT36), .B1(new_n849), .B2(new_n851), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n811), .B1(new_n853), .B2(new_n854), .ZN(G311));
  INV_X1    g430(.A(new_n811), .ZN(new_n856));
  INV_X1    g431(.A(new_n854), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n856), .B1(new_n857), .B2(new_n852), .ZN(G150));
  XOR2_X1   g433(.A(KEYINPUT104), .B(G93), .Z(new_n859));
  NAND3_X1  g434(.A1(new_n555), .A2(new_n507), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n555), .A2(G55), .A3(G543), .ZN(new_n861));
  INV_X1    g436(.A(G67), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n862), .B1(new_n505), .B2(new_n506), .ZN(new_n863));
  AND2_X1   g438(.A1(G80), .A2(G543), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n504), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n860), .A2(new_n861), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(KEYINPUT105), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT105), .ZN(new_n868));
  NAND4_X1  g443(.A1(new_n860), .A2(new_n861), .A3(new_n868), .A4(new_n865), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(G860), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(KEYINPUT37), .Z(new_n872));
  NAND2_X1  g447(.A1(new_n620), .A2(G559), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT38), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n563), .A2(new_n565), .A3(new_n866), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n867), .A2(new_n562), .A3(new_n869), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n874), .B(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT39), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(G860), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n879), .A2(new_n880), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n872), .B1(new_n883), .B2(new_n884), .ZN(G145));
  XNOR2_X1  g460(.A(KEYINPUT107), .B(G37), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n480), .B(G160), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT106), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n474), .A2(G142), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n476), .A2(G130), .ZN(new_n892));
  OR2_X1    g467(.A1(G106), .A2(G2105), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n893), .B(G2104), .C1(G118), .C2(new_n461), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n891), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(new_n646), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n896), .A2(new_n825), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n825), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n890), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n484), .A2(new_n485), .A3(new_n494), .A4(new_n493), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n744), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT98), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n732), .B(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n742), .B1(new_n905), .B2(KEYINPUT26), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n906), .A2(new_n735), .A3(new_n901), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n793), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(new_n719), .B2(new_n723), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n716), .A2(KEYINPUT96), .A3(new_n718), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n721), .A2(new_n722), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n911), .A2(new_n912), .A3(new_n793), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n908), .A2(new_n910), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n908), .B1(new_n910), .B2(new_n913), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n900), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n911), .A2(new_n912), .A3(new_n793), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n793), .B1(new_n911), .B2(new_n912), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n903), .B(new_n907), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n899), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT106), .B1(new_n920), .B2(new_n897), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n908), .A2(new_n910), .A3(new_n913), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n916), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n898), .A2(new_n890), .A3(new_n899), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT108), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n639), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n639), .ZN(new_n929));
  AOI211_X1 g504(.A(new_n929), .B(new_n926), .C1(new_n916), .C2(new_n923), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n889), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n919), .A2(new_n921), .A3(new_n922), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n921), .B1(new_n919), .B2(new_n922), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n927), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n929), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n924), .A2(new_n639), .A3(new_n927), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(new_n936), .A3(new_n888), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n887), .B1(new_n931), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT40), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n938), .B(new_n939), .ZN(G395));
  INV_X1    g515(.A(KEYINPUT110), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n941), .B1(new_n870), .B2(new_n605), .ZN(new_n942));
  XNOR2_X1  g517(.A(KEYINPUT109), .B(KEYINPUT41), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n578), .A2(new_n582), .A3(new_n584), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n945), .A2(new_n611), .A3(new_n615), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n945), .B1(new_n611), .B2(new_n615), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n616), .A2(G299), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT41), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n951), .A3(new_n946), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n619), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT79), .B1(new_n611), .B2(new_n615), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n626), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n878), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n620), .A2(new_n626), .A3(new_n877), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n953), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n950), .A2(new_n946), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n960), .B1(new_n957), .B2(new_n958), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT42), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n953), .A2(new_n957), .A3(new_n958), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT42), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n957), .A2(new_n958), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n963), .B(new_n964), .C1(new_n965), .C2(new_n960), .ZN(new_n966));
  INV_X1    g541(.A(new_n527), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n526), .B1(new_n525), .B2(new_n511), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n834), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n520), .B(new_n527), .C1(new_n833), .C2(new_n832), .ZN(new_n970));
  XNOR2_X1  g545(.A(G305), .B(G290), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n971), .B1(new_n969), .B2(new_n970), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n962), .A2(new_n966), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(G868), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n975), .B1(new_n962), .B2(new_n966), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n942), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n978), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n980), .A2(new_n941), .A3(G868), .A4(new_n976), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n979), .A2(new_n981), .ZN(G295));
  AND2_X1   g557(.A1(new_n979), .A2(new_n981), .ZN(G331));
  INV_X1    g558(.A(new_n539), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n536), .A2(KEYINPUT74), .A3(new_n537), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT75), .B1(new_n986), .B2(new_n535), .ZN(new_n987));
  INV_X1    g562(.A(new_n543), .ZN(new_n988));
  OAI21_X1  g563(.A(G171), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n542), .A2(new_n543), .A3(G301), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n989), .A2(new_n878), .A3(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n990), .ZN(new_n992));
  AOI21_X1  g567(.A(G301), .B1(new_n542), .B2(new_n543), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n877), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n950), .A2(new_n951), .A3(new_n946), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n943), .B1(new_n950), .B2(new_n946), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n991), .B(new_n994), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n960), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n992), .A2(new_n993), .A3(new_n877), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n878), .B1(new_n989), .B2(new_n990), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n974), .A2(new_n997), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G37), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n974), .B1(new_n1001), .B2(new_n997), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT43), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n960), .A2(new_n951), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n950), .A2(new_n946), .A3(new_n944), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1007), .A2(new_n994), .A3(new_n991), .A4(new_n1008), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n1001), .A2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n886), .B(new_n1002), .C1(new_n1010), .C2(new_n974), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1006), .B1(KEYINPUT43), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT44), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1013), .B1(new_n1011), .B2(KEYINPUT43), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n997), .A2(new_n1001), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n975), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT43), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1017), .A2(new_n1018), .A3(new_n1003), .A4(new_n1002), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT111), .B1(new_n1015), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1002), .A2(new_n886), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n974), .B1(new_n1001), .B2(new_n1009), .ZN(new_n1022));
  OAI21_X1  g597(.A(KEYINPUT43), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AND4_X1   g598(.A1(KEYINPUT111), .A2(new_n1023), .A3(KEYINPUT44), .A4(new_n1019), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1014), .B1(new_n1020), .B2(new_n1024), .ZN(G397));
  INV_X1    g600(.A(G1384), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n901), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT45), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n469), .A2(new_n470), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(G2105), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1031), .A2(G40), .A3(new_n463), .A4(new_n462), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G1996), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n744), .B(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(new_n793), .B(G2067), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n825), .A2(new_n827), .ZN(new_n1039));
  OR2_X1    g614(.A1(new_n825), .A2(new_n827), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g616(.A(G290), .B(G1986), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1033), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT49), .ZN(new_n1044));
  INV_X1    g619(.A(G1981), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n555), .A2(G48), .A3(G543), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n555), .A2(G86), .A3(new_n507), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n594), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1046), .A2(new_n1047), .A3(KEYINPUT116), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1045), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n596), .A2(new_n597), .A3(new_n1045), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1044), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1051), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT116), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1056), .A2(new_n1057), .A3(new_n594), .ZN(new_n1058));
  OAI211_X1 g633(.A(KEYINPUT49), .B(new_n1053), .C1(new_n1058), .C2(new_n1045), .ZN(new_n1059));
  INV_X1    g634(.A(G8), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1027), .ZN(new_n1061));
  INV_X1    g636(.A(G40), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n464), .A2(new_n471), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1060), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1055), .A2(new_n1059), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1064), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1066), .B1(new_n834), .B2(G1976), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n1068));
  INV_X1    g643(.A(G288), .ZN(new_n1069));
  XNOR2_X1  g644(.A(KEYINPUT114), .B(G1976), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1067), .B(new_n1068), .C1(KEYINPUT52), .C2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(G288), .A2(KEYINPUT91), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n587), .A2(new_n590), .A3(new_n831), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1073), .A2(G1976), .A3(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1075), .A2(new_n1064), .A3(new_n1071), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1075), .A2(new_n1068), .A3(new_n1064), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1065), .B1(new_n1072), .B2(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT112), .B(G1971), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n484), .A2(new_n485), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n493), .A2(new_n497), .A3(new_n494), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n497), .B1(new_n493), .B2(new_n494), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1083), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT45), .B1(new_n1086), .B2(new_n1026), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n901), .A2(KEYINPUT45), .A3(new_n1026), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n1063), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1082), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT50), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n901), .A2(new_n1091), .A3(new_n1026), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1092), .A2(new_n1063), .ZN(new_n1093));
  NOR2_X1   g668(.A1(G164), .A2(G1384), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1093), .B1(new_n1094), .B2(new_n1091), .ZN(new_n1095));
  XOR2_X1   g670(.A(KEYINPUT113), .B(G2090), .Z(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1090), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n520), .A2(new_n527), .A3(G8), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT55), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1102));
  OAI211_X1 g677(.A(G8), .B(new_n1098), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1099), .B(KEYINPUT55), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1028), .B1(G164), .B2(G1384), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1088), .A2(new_n1063), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1081), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1086), .A2(new_n1091), .A3(new_n1026), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1032), .B1(new_n1027), .B2(KEYINPUT50), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n1109), .A2(new_n1110), .A3(new_n1096), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1105), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1090), .B(KEYINPUT118), .C1(new_n1097), .C2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1112), .A2(new_n1114), .A3(G8), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1104), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1092), .A2(new_n1063), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1086), .A2(new_n1026), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1117), .B1(new_n1118), .B2(KEYINPUT50), .ZN(new_n1119));
  INV_X1    g694(.A(G2084), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1086), .A2(KEYINPUT45), .A3(new_n1026), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1032), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1119), .A2(new_n1120), .B1(new_n1123), .B2(new_n809), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n1124), .A2(G286), .A3(new_n1060), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1080), .A2(new_n1103), .A3(new_n1116), .A4(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g701(.A(KEYINPUT119), .B(KEYINPUT63), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1125), .A2(KEYINPUT63), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1098), .A2(G8), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1104), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1080), .A2(new_n1129), .A3(new_n1103), .A4(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1128), .A2(new_n1132), .ZN(new_n1133));
  OR2_X1    g708(.A1(G288), .A2(G1976), .ZN(new_n1134));
  OR2_X1    g709(.A1(new_n1065), .A2(new_n1134), .ZN(new_n1135));
  XOR2_X1   g710(.A(new_n1053), .B(KEYINPUT117), .Z(new_n1136));
  AOI21_X1  g711(.A(new_n1066), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1103), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1137), .B1(new_n1138), .B2(new_n1080), .ZN(new_n1139));
  NAND2_X1  g714(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT57), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n578), .A2(new_n1141), .A3(new_n582), .A4(new_n584), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g718(.A(KEYINPUT56), .B(G2072), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1106), .A2(new_n1107), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(G1956), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1143), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(G1956), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1113), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1106), .A2(new_n1107), .A3(new_n1144), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1149), .A2(new_n1140), .A3(new_n1142), .A4(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1147), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1154), .A2(KEYINPUT61), .A3(new_n1140), .A4(new_n1142), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1087), .A2(G1996), .A3(new_n1089), .ZN(new_n1157));
  XNOR2_X1  g732(.A(KEYINPUT58), .B(G1341), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1158), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n567), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT59), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT60), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1162), .B1(new_n618), .B2(new_n619), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1027), .A2(new_n1032), .A3(G2067), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT120), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1164), .B(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1095), .A2(new_n757), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n618), .A2(new_n1162), .A3(new_n619), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1163), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  AND4_X1   g745(.A1(KEYINPUT60), .A2(new_n620), .A3(new_n1167), .A4(new_n1166), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1156), .B(new_n1161), .C1(new_n1170), .C2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1168), .B1(new_n618), .B2(new_n619), .ZN(new_n1173));
  OR2_X1    g748(.A1(new_n1143), .A2(KEYINPUT121), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1154), .B1(KEYINPUT121), .B2(new_n1143), .ZN(new_n1175));
  AOI22_X1  g750(.A1(new_n1173), .A2(new_n1151), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1172), .A2(new_n1176), .ZN(new_n1177));
  XOR2_X1   g752(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1178));
  INV_X1    g753(.A(KEYINPUT53), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1106), .A2(new_n1107), .A3(new_n443), .ZN(new_n1180));
  AOI22_X1  g755(.A1(new_n1179), .A2(new_n1180), .B1(new_n1095), .B2(new_n771), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n443), .A2(KEYINPUT53), .ZN(new_n1182));
  OR2_X1    g757(.A1(new_n1123), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(G301), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1180), .A2(new_n1179), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1095), .A2(new_n771), .ZN(new_n1186));
  OR2_X1    g761(.A1(new_n1032), .A2(KEYINPUT123), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1182), .B1(new_n1032), .B2(KEYINPUT123), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1187), .A2(new_n1188), .A3(new_n1029), .A4(new_n1088), .ZN(new_n1189));
  AND4_X1   g764(.A1(G301), .A2(new_n1185), .A3(new_n1186), .A4(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1178), .B1(new_n1184), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1191), .A2(KEYINPUT124), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT124), .ZN(new_n1193));
  OAI211_X1 g768(.A(new_n1193), .B(new_n1178), .C1(new_n1184), .C2(new_n1190), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1177), .A2(new_n1195), .ZN(new_n1196));
  AND3_X1   g771(.A1(new_n1080), .A2(new_n1103), .A3(new_n1116), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1181), .A2(new_n1189), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT125), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1181), .A2(KEYINPUT125), .A3(new_n1189), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1200), .A2(new_n1201), .A3(G171), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1181), .A2(G301), .A3(new_n1183), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1202), .A2(KEYINPUT54), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1123), .A2(new_n809), .ZN(new_n1205));
  OAI211_X1 g780(.A(new_n1093), .B(new_n1120), .C1(new_n1094), .C2(new_n1091), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g782(.A(G8), .B1(new_n1207), .B2(G286), .ZN(new_n1208));
  NOR2_X1   g783(.A1(new_n1124), .A2(G168), .ZN(new_n1209));
  OAI21_X1  g784(.A(KEYINPUT51), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1060), .B1(new_n1124), .B2(G168), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT51), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1210), .A2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g789(.A1(new_n1197), .A2(new_n1204), .A3(new_n1214), .ZN(new_n1215));
  OAI211_X1 g790(.A(new_n1133), .B(new_n1139), .C1(new_n1196), .C2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1207), .A2(G286), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1212), .B1(new_n1211), .B2(new_n1217), .ZN(new_n1218));
  NOR2_X1   g793(.A1(new_n1208), .A2(KEYINPUT51), .ZN(new_n1219));
  OAI21_X1  g794(.A(KEYINPUT62), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g795(.A(KEYINPUT62), .ZN(new_n1221));
  NAND3_X1  g796(.A1(new_n1210), .A2(new_n1221), .A3(new_n1213), .ZN(new_n1222));
  NAND3_X1  g797(.A1(new_n1220), .A2(new_n1184), .A3(new_n1222), .ZN(new_n1223));
  NAND3_X1  g798(.A1(new_n1080), .A2(new_n1103), .A3(new_n1116), .ZN(new_n1224));
  OAI21_X1  g799(.A(KEYINPUT126), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g800(.A(new_n1184), .ZN(new_n1226));
  AOI21_X1  g801(.A(new_n1226), .B1(new_n1214), .B2(KEYINPUT62), .ZN(new_n1227));
  INV_X1    g802(.A(KEYINPUT126), .ZN(new_n1228));
  NAND4_X1  g803(.A1(new_n1227), .A2(new_n1228), .A3(new_n1197), .A4(new_n1222), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1225), .A2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g805(.A(new_n1043), .B1(new_n1216), .B2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g806(.A1(new_n1036), .A2(new_n735), .A3(new_n906), .ZN(new_n1232));
  INV_X1    g807(.A(KEYINPUT46), .ZN(new_n1233));
  NAND2_X1  g808(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1234));
  AOI22_X1  g809(.A1(new_n1232), .A2(new_n1033), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g810(.A(new_n1235), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1236));
  XNOR2_X1  g811(.A(new_n1236), .B(KEYINPUT47), .ZN(new_n1237));
  AND2_X1   g812(.A1(new_n1041), .A2(new_n1033), .ZN(new_n1238));
  NAND3_X1  g813(.A1(new_n1033), .A2(new_n815), .A3(new_n812), .ZN(new_n1239));
  XOR2_X1   g814(.A(new_n1239), .B(KEYINPUT48), .Z(new_n1240));
  OAI21_X1  g815(.A(new_n1237), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g816(.A(new_n1039), .B1(new_n1037), .B2(new_n1033), .ZN(new_n1242));
  INV_X1    g817(.A(G2067), .ZN(new_n1243));
  AOI21_X1  g818(.A(new_n1242), .B1(new_n1243), .B2(new_n793), .ZN(new_n1244));
  OR2_X1    g819(.A1(new_n1244), .A2(KEYINPUT127), .ZN(new_n1245));
  INV_X1    g820(.A(new_n1033), .ZN(new_n1246));
  AOI21_X1  g821(.A(new_n1246), .B1(new_n1244), .B2(KEYINPUT127), .ZN(new_n1247));
  AOI21_X1  g822(.A(new_n1241), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g823(.A1(new_n1231), .A2(new_n1248), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g824(.A(G319), .ZN(new_n1251));
  NOR3_X1   g825(.A1(G401), .A2(G227), .A3(new_n1251), .ZN(new_n1252));
  NAND3_X1  g826(.A1(new_n704), .A2(new_n705), .A3(new_n1252), .ZN(new_n1253));
  NAND2_X1  g827(.A1(new_n931), .A2(new_n937), .ZN(new_n1254));
  AOI21_X1  g828(.A(new_n1253), .B1(new_n1254), .B2(new_n886), .ZN(new_n1255));
  AND2_X1   g829(.A1(new_n1255), .A2(new_n1012), .ZN(G308));
  NAND2_X1  g830(.A1(new_n1255), .A2(new_n1012), .ZN(G225));
endmodule


