//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 1 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1297,
    new_n1298, new_n1299, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n202), .A2(G50), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G107), .ZN(new_n223));
  INV_X1    g0023(.A(G264), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n205), .B1(new_n219), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n208), .B1(new_n212), .B2(new_n213), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XOR2_X1   g0038(.A(G107), .B(G116), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(G169), .ZN(new_n245));
  NOR2_X1   g0045(.A1(new_n245), .A2(KEYINPUT74), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT3), .B(G33), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n247), .A2(G226), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(G33), .A2(G97), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n247), .A2(G1698), .ZN(new_n251));
  OAI211_X1 g0051(.A(new_n249), .B(new_n250), .C1(new_n251), .C2(new_n230), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n209), .B1(G33), .B2(G41), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT13), .ZN(new_n255));
  INV_X1    g0055(.A(G274), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n258));
  NOR3_X1   g0058(.A1(new_n253), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  OAI211_X1 g0061(.A(G1), .B(G13), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n258), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n259), .B1(G238), .B2(new_n264), .ZN(new_n265));
  AND3_X1   g0065(.A1(new_n254), .A2(new_n255), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n255), .B1(new_n254), .B2(new_n265), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n246), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OR2_X1    g0068(.A1(new_n268), .A2(KEYINPUT14), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n266), .A2(new_n267), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G179), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n268), .A2(KEYINPUT14), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n257), .A2(G13), .A3(G20), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n215), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n276), .B(KEYINPUT12), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT65), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(new_n205), .B2(new_n260), .ZN(new_n279));
  NAND4_X1  g0079(.A1(KEYINPUT65), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n279), .A2(new_n209), .A3(new_n280), .A4(new_n274), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n210), .A2(G1), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n282), .A2(G68), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(KEYINPUT73), .B1(new_n277), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n279), .A2(new_n209), .A3(new_n280), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G20), .A2(G33), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G50), .ZN(new_n290));
  OAI22_X1  g0090(.A1(new_n289), .A2(new_n290), .B1(new_n210), .B2(G68), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n260), .A2(new_n221), .A3(G20), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n287), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT11), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n277), .A2(KEYINPUT73), .A3(new_n285), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n273), .B1(new_n286), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n270), .A2(G190), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n296), .A2(new_n286), .ZN(new_n299));
  INV_X1    g0099(.A(G200), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n298), .B(new_n299), .C1(new_n300), .C2(new_n270), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n259), .B1(G244), .B2(new_n264), .ZN(new_n303));
  NOR2_X1   g0103(.A1(G232), .A2(G1698), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n248), .A2(G238), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n247), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n306), .B(new_n253), .C1(G107), .C2(new_n247), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT68), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n303), .A2(KEYINPUT68), .A3(new_n307), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OR2_X1    g0112(.A1(new_n312), .A2(G179), .ZN(new_n313));
  INV_X1    g0113(.A(new_n287), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n288), .A2(KEYINPUT69), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT8), .B(G58), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n288), .A2(KEYINPUT69), .ZN(new_n317));
  OR3_X1    g0117(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT15), .B(G87), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n260), .A2(G20), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n320), .A2(new_n321), .B1(G20), .B2(G77), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n314), .B1(new_n318), .B2(new_n322), .ZN(new_n323));
  NOR3_X1   g0123(.A1(new_n281), .A2(new_n221), .A3(new_n283), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n274), .A2(G77), .ZN(new_n325));
  NOR3_X1   g0125(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n312), .A2(new_n245), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n313), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n310), .A2(G200), .A3(new_n311), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(KEYINPUT70), .A3(new_n326), .ZN(new_n332));
  INV_X1    g0132(.A(G190), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n332), .B1(new_n333), .B2(new_n312), .ZN(new_n334));
  AOI21_X1  g0134(.A(KEYINPUT70), .B1(new_n331), .B2(new_n326), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OR3_X1    g0136(.A1(new_n330), .A2(new_n336), .A3(KEYINPUT71), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n282), .A2(G50), .A3(new_n284), .ZN(new_n338));
  OAI21_X1  g0138(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n339));
  INV_X1    g0139(.A(G150), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n339), .B1(new_n340), .B2(new_n289), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n316), .B(KEYINPUT66), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n341), .B1(new_n342), .B2(new_n321), .ZN(new_n343));
  OAI221_X1 g0143(.A(new_n338), .B1(G50), .B2(new_n274), .C1(new_n343), .C2(new_n314), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n259), .B1(G226), .B2(new_n264), .ZN(new_n345));
  INV_X1    g0145(.A(G223), .ZN(new_n346));
  OAI22_X1  g0146(.A1(new_n251), .A2(new_n346), .B1(new_n221), .B2(new_n247), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n247), .A2(G222), .A3(new_n248), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT64), .ZN(new_n349));
  OR2_X1    g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n349), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n347), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n345), .B1(new_n352), .B2(new_n262), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n344), .B1(new_n354), .B2(G169), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n353), .A2(G179), .ZN(new_n356));
  OR2_X1    g0156(.A1(new_n356), .A2(KEYINPUT67), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(KEYINPUT67), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n355), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g0159(.A(new_n344), .B(KEYINPUT9), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n353), .A2(G200), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT72), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n362), .B1(new_n354), .B2(G190), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n360), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT10), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT10), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n360), .A2(new_n366), .A3(new_n361), .A4(new_n363), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n359), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT71), .B1(new_n330), .B2(new_n336), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n302), .A2(new_n337), .A3(new_n368), .A4(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT79), .ZN(new_n371));
  INV_X1    g0171(.A(G58), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n372), .A2(new_n215), .ZN(new_n373));
  OR2_X1    g0173(.A1(new_n373), .A2(new_n201), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n374), .A2(G20), .B1(G159), .B2(new_n288), .ZN(new_n375));
  AND2_X1   g0175(.A1(KEYINPUT75), .A2(G33), .ZN(new_n376));
  NOR2_X1   g0176(.A1(KEYINPUT75), .A2(G33), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT3), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(KEYINPUT3), .A2(G33), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n210), .A2(KEYINPUT7), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT3), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT75), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n260), .ZN(new_n386));
  NAND2_X1  g0186(.A1(KEYINPUT75), .A2(G33), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n384), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NOR3_X1   g0188(.A1(new_n388), .A2(KEYINPUT76), .A3(new_n379), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT76), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n378), .B2(new_n380), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n210), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT7), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n383), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI211_X1 g0194(.A(KEYINPUT16), .B(new_n375), .C1(new_n394), .C2(new_n215), .ZN(new_n395));
  AND2_X1   g0195(.A1(KEYINPUT3), .A2(G33), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n396), .A2(new_n379), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n210), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n382), .A2(new_n396), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n386), .A2(new_n384), .A3(new_n387), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n398), .A2(new_n393), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n375), .B1(new_n401), .B2(new_n215), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT16), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n395), .A2(new_n404), .A3(new_n287), .ZN(new_n405));
  INV_X1    g0205(.A(new_n342), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n406), .A2(new_n283), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n407), .A2(new_n282), .B1(new_n275), .B2(new_n406), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n259), .B1(G232), .B2(new_n264), .ZN(new_n409));
  NOR2_X1   g0209(.A1(G223), .A2(G1698), .ZN(new_n410));
  INV_X1    g0210(.A(G226), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n410), .B1(new_n411), .B2(G1698), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n381), .A2(new_n412), .B1(G33), .B2(G87), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n409), .B1(new_n262), .B2(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n414), .A2(G179), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n386), .A2(new_n387), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n379), .B1(new_n416), .B2(KEYINPUT3), .ZN(new_n417));
  INV_X1    g0217(.A(new_n412), .ZN(new_n418));
  OAI22_X1  g0218(.A1(new_n417), .A2(new_n418), .B1(new_n260), .B2(new_n217), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n253), .ZN(new_n420));
  AOI21_X1  g0220(.A(G169), .B1(new_n420), .B2(new_n409), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT77), .B1(new_n415), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n414), .A2(new_n245), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT77), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n423), .B(new_n424), .C1(G179), .C2(new_n414), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n405), .A2(new_n408), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  XNOR2_X1  g0226(.A(new_n426), .B(KEYINPUT18), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n414), .A2(new_n300), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n428), .B1(G190), .B2(new_n414), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n405), .A2(new_n408), .A3(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT17), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n405), .A2(new_n429), .A3(KEYINPUT17), .A4(new_n408), .ZN(new_n433));
  AND3_X1   g0233(.A1(new_n432), .A2(KEYINPUT78), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT78), .B1(new_n432), .B2(new_n433), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n427), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OR3_X1    g0236(.A1(new_n370), .A2(new_n371), .A3(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n371), .B1(new_n370), .B2(new_n436), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n262), .A2(G274), .ZN(new_n441));
  INV_X1    g0241(.A(G45), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n442), .A2(G1), .ZN(new_n443));
  AND2_X1   g0243(.A1(KEYINPUT5), .A2(G41), .ZN(new_n444));
  NOR2_X1   g0244(.A1(KEYINPUT5), .A2(G41), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n441), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n262), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n447), .B1(G257), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT4), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(new_n222), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n452), .B(new_n248), .C1(new_n379), .C2(new_n396), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G33), .A2(G283), .ZN(new_n454));
  OAI211_X1 g0254(.A(G250), .B(G1698), .C1(new_n396), .C2(new_n379), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n381), .A2(G244), .A3(new_n248), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n456), .B1(new_n457), .B2(new_n451), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n450), .B1(new_n458), .B2(new_n262), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n245), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n223), .A2(KEYINPUT80), .A3(KEYINPUT6), .A4(G97), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT80), .ZN(new_n462));
  NAND2_X1  g0262(.A1(KEYINPUT6), .A2(G97), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n462), .B1(new_n463), .B2(G107), .ZN(new_n464));
  AND2_X1   g0264(.A1(G97), .A2(G107), .ZN(new_n465));
  NOR2_X1   g0265(.A1(G97), .A2(G107), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n461), .B(new_n464), .C1(new_n467), .C2(KEYINPUT6), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G20), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n288), .A2(G77), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n469), .B(new_n470), .C1(new_n401), .C2(new_n223), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n287), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n274), .A2(G97), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n280), .A2(new_n209), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n260), .A2(G1), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n475), .A2(new_n279), .A3(new_n274), .A4(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(G97), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n474), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n472), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(G179), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n483), .B(new_n450), .C1(new_n458), .C2(new_n262), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n460), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n480), .B1(new_n471), .B2(new_n287), .ZN(new_n486));
  OAI211_X1 g0286(.A(G190), .B(new_n450), .C1(new_n458), .C2(new_n262), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n253), .A2(new_n256), .ZN(new_n488));
  OR2_X1    g0288(.A1(new_n444), .A2(new_n445), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(new_n443), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(G257), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n490), .B1(new_n491), .B2(new_n448), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n493));
  AOI211_X1 g0293(.A(new_n222), .B(G1698), .C1(new_n378), .C2(new_n380), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n493), .B1(new_n494), .B2(KEYINPUT4), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n492), .B1(new_n495), .B2(new_n253), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n486), .B(new_n487), .C1(new_n496), .C2(new_n300), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n485), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT81), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n281), .A2(new_n476), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G116), .ZN(new_n501));
  XNOR2_X1  g0301(.A(KEYINPUT82), .B(G116), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n275), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n260), .A2(G97), .ZN(new_n504));
  AOI21_X1  g0304(.A(G20), .B1(G33), .B2(G283), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n502), .A2(G20), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n506), .A2(KEYINPUT20), .A3(new_n287), .ZN(new_n507));
  AOI21_X1  g0307(.A(KEYINPUT20), .B1(new_n506), .B2(new_n287), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n501), .B(new_n503), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n446), .A2(G270), .A3(new_n262), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT86), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n446), .A2(KEYINPUT86), .A3(G270), .A4(new_n262), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n224), .A2(G1698), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(G257), .B2(G1698), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n516), .B1(new_n380), .B2(new_n378), .ZN(new_n517));
  INV_X1    g0317(.A(G303), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n247), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n253), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n514), .A2(new_n490), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n509), .A2(new_n521), .A3(G169), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT21), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n521), .A2(G200), .ZN(new_n525));
  INV_X1    g0325(.A(new_n509), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n514), .A2(new_n520), .A3(G190), .A4(new_n490), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AND4_X1   g0328(.A1(G179), .A2(new_n514), .A3(new_n490), .A4(new_n520), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n509), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n509), .A2(new_n521), .A3(KEYINPUT21), .A4(G169), .ZN(new_n531));
  AND4_X1   g0331(.A1(new_n524), .A2(new_n528), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT81), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n485), .A2(new_n533), .A3(new_n497), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n499), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n216), .A2(G1698), .ZN(new_n536));
  INV_X1    g0336(.A(new_n502), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n381), .A2(new_n536), .B1(new_n416), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n381), .A2(G244), .A3(G1698), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n262), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n443), .A2(new_n218), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n488), .A2(new_n443), .B1(new_n262), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(G169), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n537), .A2(new_n416), .ZN(new_n545));
  INV_X1    g0345(.A(new_n536), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n417), .B2(new_n546), .ZN(new_n547));
  AOI211_X1 g0347(.A(new_n222), .B(new_n248), .C1(new_n378), .C2(new_n380), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n253), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n549), .A2(G179), .A3(new_n542), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n544), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n210), .A2(new_n552), .B1(new_n466), .B2(new_n217), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n210), .A2(G33), .A3(G97), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT19), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT83), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n554), .A2(KEYINPUT83), .A3(new_n555), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n553), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n381), .A2(new_n210), .A3(G68), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n314), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n320), .A2(new_n274), .ZN(new_n563));
  OAI21_X1  g0363(.A(KEYINPUT84), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI211_X1 g0364(.A(G20), .B(new_n215), .C1(new_n378), .C2(new_n380), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n552), .A2(new_n210), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n466), .A2(new_n217), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n554), .A2(KEYINPUT83), .A3(new_n555), .ZN(new_n569));
  AOI21_X1  g0369(.A(KEYINPUT83), .B1(new_n554), .B2(new_n555), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n287), .B1(new_n565), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT84), .ZN(new_n573));
  INV_X1    g0373(.A(new_n563), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n564), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n478), .A2(new_n319), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT85), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT85), .ZN(new_n580));
  AOI211_X1 g0380(.A(new_n580), .B(new_n577), .C1(new_n564), .C2(new_n575), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n551), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n500), .A2(G87), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n562), .A2(KEYINPUT84), .A3(new_n563), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n573), .B1(new_n572), .B2(new_n574), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n549), .A2(G190), .A3(new_n542), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n540), .A2(new_n543), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n587), .B1(new_n588), .B2(new_n300), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n582), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n535), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT91), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT90), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n491), .A2(new_n248), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n388), .B2(new_n379), .ZN(new_n597));
  INV_X1    g0397(.A(G294), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n598), .B1(new_n386), .B2(new_n387), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n248), .A2(G250), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n601), .B1(new_n378), .B2(new_n380), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT89), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n597), .B(new_n600), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n417), .A2(KEYINPUT89), .A3(new_n601), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n595), .B(new_n253), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n448), .A2(new_n224), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n607), .A2(new_n447), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(KEYINPUT89), .B1(new_n417), .B2(new_n601), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n599), .B1(new_n381), .B2(new_n596), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n602), .A2(new_n603), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n595), .B1(new_n613), .B2(new_n253), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n594), .B1(new_n609), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n613), .A2(new_n253), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(KEYINPUT90), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n617), .A2(KEYINPUT91), .A3(new_n606), .A4(new_n608), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n615), .A2(new_n618), .A3(new_n333), .ZN(new_n619));
  AOI211_X1 g0419(.A(new_n607), .B(new_n447), .C1(new_n613), .C2(new_n253), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n619), .B1(G200), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(KEYINPUT22), .A2(G87), .ZN(new_n622));
  AOI211_X1 g0422(.A(G20), .B(new_n622), .C1(new_n378), .C2(new_n380), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n217), .A2(G20), .ZN(new_n624));
  AOI21_X1  g0424(.A(KEYINPUT22), .B1(new_n247), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(KEYINPUT87), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT87), .ZN(new_n627));
  INV_X1    g0427(.A(new_n625), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n381), .A2(new_n210), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n627), .B(new_n628), .C1(new_n629), .C2(new_n622), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT88), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n632), .A2(KEYINPUT24), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n210), .A2(G107), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT23), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n634), .A2(new_n635), .B1(new_n632), .B2(KEYINPUT24), .ZN(new_n636));
  OAI221_X1 g0436(.A(new_n636), .B1(new_n635), .B2(new_n634), .C1(new_n545), .C2(G20), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n631), .A2(new_n633), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n633), .B1(new_n631), .B2(new_n638), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n287), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n275), .A2(new_n223), .ZN(new_n642));
  XNOR2_X1  g0442(.A(new_n642), .B(KEYINPUT25), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n643), .B1(G107), .B2(new_n500), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n621), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n245), .B1(new_n615), .B2(new_n618), .ZN(new_n648));
  INV_X1    g0448(.A(new_n607), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n616), .A2(new_n649), .A3(new_n490), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n650), .A2(new_n483), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n645), .B1(new_n648), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(KEYINPUT92), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT92), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n645), .B(new_n654), .C1(new_n648), .C2(new_n651), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n593), .A2(new_n647), .A3(new_n653), .A4(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n440), .A2(new_n656), .ZN(G372));
  AND3_X1   g0457(.A1(new_n524), .A2(new_n530), .A3(new_n531), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n652), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n578), .B1(new_n584), .B2(new_n585), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n580), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n576), .A2(KEYINPUT85), .A3(new_n578), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT93), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n544), .A2(new_n550), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n664), .B1(new_n544), .B2(new_n550), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI211_X1 g0468(.A(new_n590), .B(new_n498), .C1(new_n663), .C2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n659), .A2(new_n669), .A3(new_n647), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n663), .A2(new_n668), .ZN(new_n671));
  INV_X1    g0471(.A(new_n485), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n582), .A2(new_n591), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(KEYINPUT26), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n671), .A2(new_n675), .A3(new_n591), .A4(new_n672), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n670), .A2(new_n671), .A3(new_n674), .A4(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n439), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n435), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n432), .A2(KEYINPUT78), .A3(new_n433), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n330), .A2(new_n301), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n297), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n427), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n365), .A2(new_n367), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n359), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n678), .A2(new_n687), .ZN(G369));
  AND2_X1   g0488(.A1(new_n653), .A2(new_n655), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n689), .A2(new_n647), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n257), .A2(new_n210), .A3(G13), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G213), .A3(new_n693), .ZN(new_n694));
  XOR2_X1   g0494(.A(new_n694), .B(KEYINPUT94), .Z(new_n695));
  INV_X1    g0495(.A(G343), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n690), .B1(new_n646), .B2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n652), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n697), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n697), .A2(new_n509), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n532), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n658), .B2(new_n703), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G330), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n700), .A2(new_n698), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n658), .A2(new_n697), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n690), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n708), .A2(new_n709), .A3(new_n711), .ZN(G399));
  INV_X1    g0512(.A(new_n206), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G41), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n567), .A2(G116), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(G1), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(new_n213), .B2(new_n715), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT28), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n677), .A2(new_n698), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(KEYINPUT29), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n653), .A2(new_n655), .A3(new_n658), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT98), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n669), .A2(new_n647), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT98), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n653), .A2(new_n725), .A3(new_n655), .A4(new_n658), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n723), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n671), .B1(new_n673), .B2(KEYINPUT26), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n590), .B1(new_n663), .B2(new_n668), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n675), .B1(new_n729), .B2(new_n672), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n698), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n721), .B1(new_n733), .B2(KEYINPUT29), .ZN(new_n734));
  INV_X1    g0534(.A(G330), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n607), .B1(new_n613), .B2(new_n253), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n529), .A2(new_n736), .A3(new_n588), .A4(new_n496), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT95), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(KEYINPUT30), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT96), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(new_n620), .B2(new_n496), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n650), .A2(KEYINPUT96), .A3(new_n459), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n521), .A2(new_n483), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(new_n588), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n742), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT30), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n737), .A2(new_n738), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n740), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(new_n697), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT31), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n749), .A2(KEYINPUT31), .A3(new_n697), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n752), .A2(KEYINPUT97), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(KEYINPUT31), .B1(new_n749), .B2(new_n697), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT97), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n689), .A2(new_n647), .A3(new_n593), .A4(new_n698), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n735), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n734), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n719), .B1(new_n763), .B2(G1), .ZN(G364));
  AND2_X1   g0564(.A1(new_n210), .A2(G13), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n257), .B1(new_n765), .B2(G45), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n714), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n247), .A2(new_n206), .ZN(new_n769));
  INV_X1    g0569(.A(G355), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n769), .A2(new_n770), .B1(G116), .B2(new_n206), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n389), .A2(new_n391), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n713), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n213), .A2(G45), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n774), .B1(new_n243), .B2(G45), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n771), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G13), .A2(G33), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n209), .B1(G20), .B2(new_n245), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n768), .B1(new_n776), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n210), .A2(new_n333), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n784), .A2(G179), .A3(new_n300), .ZN(new_n785));
  INV_X1    g0585(.A(G322), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n210), .A2(G190), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n787), .A2(G179), .A3(new_n300), .ZN(new_n788));
  INV_X1    g0588(.A(G311), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n785), .A2(new_n786), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n300), .A2(G179), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n784), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n247), .B(new_n790), .C1(G303), .C2(new_n793), .ZN(new_n794));
  OR3_X1    g0594(.A1(new_n210), .A2(KEYINPUT100), .A3(G190), .ZN(new_n795));
  OAI21_X1  g0595(.A(KEYINPUT100), .B1(new_n210), .B2(G190), .ZN(new_n796));
  NOR2_X1   g0596(.A1(G179), .A2(G200), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G329), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n795), .A2(new_n796), .A3(new_n791), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G283), .ZN(new_n803));
  AND3_X1   g0603(.A1(new_n794), .A2(new_n800), .A3(new_n803), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n333), .A2(G179), .A3(G200), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n210), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n333), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n807), .A2(G294), .B1(G326), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n808), .A2(G190), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  XOR2_X1   g0612(.A(KEYINPUT33), .B(G317), .Z(new_n813));
  OAI211_X1 g0613(.A(new_n804), .B(new_n810), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n809), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(new_n290), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n806), .A2(new_n479), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n816), .B(new_n817), .C1(G68), .C2(new_n811), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n788), .A2(KEYINPUT99), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n788), .A2(KEYINPUT99), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(G77), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n247), .B1(new_n792), .B2(new_n217), .C1(new_n372), .C2(new_n785), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(G107), .B2(new_n802), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n818), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(G159), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n798), .A2(new_n827), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT32), .Z(new_n829));
  OAI21_X1  g0629(.A(new_n814), .B1(new_n826), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n783), .B1(new_n830), .B2(new_n780), .ZN(new_n831));
  INV_X1    g0631(.A(new_n779), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n831), .B1(new_n705), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n768), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n706), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n705), .A2(G330), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n833), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g0637(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n837), .B(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(G396));
  NOR2_X1   g0640(.A1(new_n780), .A2(new_n777), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n834), .B1(new_n221), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n780), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n817), .B1(G283), .B2(new_n811), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n518), .B2(new_n815), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n821), .A2(new_n502), .B1(new_n789), .B2(new_n798), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n801), .A2(new_n217), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n397), .B1(new_n792), .B2(new_n223), .C1(new_n598), .C2(new_n785), .ZN(new_n848));
  NOR4_X1   g0648(.A1(new_n845), .A2(new_n846), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n807), .A2(G58), .B1(new_n793), .B2(G50), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n812), .A2(new_n340), .ZN(new_n851));
  INV_X1    g0651(.A(G137), .ZN(new_n852));
  INV_X1    g0652(.A(G143), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n852), .A2(new_n815), .B1(new_n785), .B2(new_n853), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n851), .B(new_n854), .C1(G159), .C2(new_n822), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n850), .B1(new_n215), .B2(new_n801), .C1(new_n855), .C2(KEYINPUT34), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(KEYINPUT34), .B2(new_n855), .ZN(new_n857));
  INV_X1    g0657(.A(G132), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n772), .B1(new_n858), .B2(new_n798), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT103), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n849), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n329), .A2(new_n697), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n697), .A2(new_n327), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT104), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n863), .B(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n335), .B2(new_n334), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n862), .B1(new_n866), .B2(new_n329), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n842), .B1(new_n843), .B2(new_n861), .C1(new_n867), .C2(new_n778), .ZN(new_n868));
  AND3_X1   g0668(.A1(new_n659), .A2(new_n669), .A3(new_n647), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n674), .A2(new_n676), .A3(new_n671), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n698), .B(new_n867), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT105), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n677), .A2(KEYINPUT105), .A3(new_n698), .A4(new_n867), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n867), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n720), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n768), .B1(new_n878), .B2(new_n761), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n878), .A2(new_n761), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n868), .B1(new_n880), .B2(new_n881), .ZN(G384));
  INV_X1    g0682(.A(G116), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n883), .B(new_n212), .C1(new_n468), .C2(KEYINPUT35), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(KEYINPUT35), .B2(new_n468), .ZN(new_n885));
  XOR2_X1   g0685(.A(new_n885), .B(KEYINPUT36), .Z(new_n886));
  OR3_X1    g0686(.A1(new_n213), .A2(new_n221), .A3(new_n373), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n290), .A2(G68), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n257), .B(G13), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n698), .A2(new_n299), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n297), .A2(new_n301), .A3(new_n892), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n273), .A2(new_n891), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n862), .B1(new_n873), .B2(new_n874), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT106), .ZN(new_n897));
  INV_X1    g0697(.A(new_n408), .ZN(new_n898));
  INV_X1    g0698(.A(new_n375), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT76), .B1(new_n388), .B2(new_n379), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n378), .A2(new_n390), .A3(new_n380), .ZN(new_n901));
  AOI21_X1  g0701(.A(G20), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI22_X1  g0702(.A1(new_n902), .A2(KEYINPUT7), .B1(new_n382), .B2(new_n381), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n899), .B1(new_n903), .B2(G68), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n314), .B1(new_n904), .B2(KEYINPUT16), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n375), .B1(new_n394), .B2(new_n215), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n403), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n898), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n897), .B1(new_n908), .B2(new_n695), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n395), .A2(new_n287), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n904), .A2(KEYINPUT16), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n408), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n695), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n912), .A2(KEYINPUT106), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n909), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n436), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n422), .A2(new_n425), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n912), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n909), .A2(new_n914), .A3(new_n430), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(KEYINPUT37), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n405), .A2(new_n408), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n917), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n913), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n922), .A2(new_n923), .A3(new_n430), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n924), .A2(KEYINPUT37), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n920), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n916), .A2(new_n926), .A3(KEYINPUT38), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n916), .A2(new_n926), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT38), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI211_X1 g0730(.A(new_n895), .B(new_n896), .C1(new_n927), .C2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT37), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n924), .B(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n432), .A2(new_n433), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n923), .B1(new_n427), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n929), .B1(new_n933), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n927), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT39), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n930), .A2(KEYINPUT39), .A3(new_n927), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n297), .A2(new_n697), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n942), .A2(new_n944), .B1(new_n427), .B2(new_n913), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n931), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n687), .B1(new_n734), .B2(new_n440), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n946), .B(new_n947), .Z(new_n948));
  AND3_X1   g0748(.A1(new_n749), .A2(KEYINPUT31), .A3(new_n697), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n949), .A2(new_n755), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n656), .B2(new_n697), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(KEYINPUT108), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT108), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n953), .B(new_n950), .C1(new_n656), .C2(new_n697), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n895), .A2(new_n876), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n955), .A2(KEYINPUT40), .A3(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT109), .ZN(new_n959));
  AND3_X1   g0759(.A1(new_n927), .A2(new_n937), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n959), .B1(new_n927), .B2(new_n937), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n930), .A2(new_n927), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n963), .A2(new_n955), .A3(new_n956), .ZN(new_n964));
  XOR2_X1   g0764(.A(KEYINPUT107), .B(KEYINPUT40), .Z(new_n965));
  AOI22_X1  g0765(.A1(new_n958), .A2(new_n962), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AND2_X1   g0766(.A1(new_n439), .A2(new_n955), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n735), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n967), .B2(new_n966), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n948), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n257), .B2(new_n765), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n948), .A2(new_n969), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n890), .B1(new_n971), .B2(new_n972), .ZN(G367));
  INV_X1    g0773(.A(new_n773), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n781), .B1(new_n206), .B2(new_n319), .C1(new_n974), .C2(new_n236), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n975), .A2(new_n768), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n822), .A2(G50), .B1(G77), .B2(new_n802), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n812), .A2(new_n827), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n815), .A2(new_n853), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n978), .B(new_n979), .C1(G68), .C2(new_n807), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n247), .B1(new_n792), .B2(new_n372), .C1(new_n340), .C2(new_n785), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(G137), .B2(new_n799), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n977), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n793), .A2(KEYINPUT46), .A3(G116), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n984), .B1(new_n518), .B2(new_n785), .C1(new_n815), .C2(new_n789), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(G283), .B2(new_n822), .ZN(new_n986));
  INV_X1    g0786(.A(G317), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n986), .B1(new_n479), .B2(new_n801), .C1(new_n987), .C2(new_n798), .ZN(new_n988));
  INV_X1    g0788(.A(new_n772), .ZN(new_n989));
  XNOR2_X1  g0789(.A(KEYINPUT111), .B(KEYINPUT46), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n792), .B2(new_n502), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n807), .A2(G107), .B1(G294), .B2(new_n811), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n989), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n983), .B1(new_n988), .B2(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT47), .Z(new_n995));
  NAND2_X1  g0795(.A1(new_n586), .A2(new_n697), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n671), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n729), .A2(new_n996), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n976), .B1(new_n995), .B2(new_n843), .C1(new_n832), .C2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n711), .A2(new_n709), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n485), .B(new_n497), .C1(new_n486), .C2(new_n698), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n485), .B2(new_n698), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT44), .Z(new_n1006));
  NOR2_X1   g0806(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT45), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n708), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1006), .A2(new_n708), .A3(new_n1008), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n702), .A2(new_n710), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n711), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n707), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1014), .A2(new_n706), .A3(new_n711), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n763), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n763), .B1(new_n1013), .B2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n714), .B(KEYINPUT41), .Z(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n767), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n711), .A2(new_n1004), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT42), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n485), .B1(new_n689), .B2(new_n1002), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n698), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n999), .A2(KEYINPUT43), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(KEYINPUT110), .B(KEYINPUT43), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n997), .A2(new_n998), .A3(new_n1030), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1028), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1010), .A2(new_n1003), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1033), .B(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1000), .B1(new_n1023), .B2(new_n1035), .ZN(G387));
  NAND3_X1  g0836(.A1(new_n699), .A2(new_n701), .A3(new_n779), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n769), .A2(new_n716), .B1(G107), .B2(new_n206), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n233), .A2(new_n442), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n716), .B(new_n442), .C1(new_n215), .C2(new_n221), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT50), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n316), .B2(G50), .ZN(new_n1042));
  OR3_X1    g0842(.A1(new_n316), .A2(new_n1041), .A3(G50), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1040), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n974), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1038), .B1(new_n1039), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n768), .B1(new_n1046), .B2(new_n782), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n806), .A2(new_n319), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n788), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n1049), .A2(G68), .B1(new_n793), .B2(G77), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n290), .B2(new_n785), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n1048), .B(new_n1051), .C1(G159), .C2(new_n809), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n799), .A2(G150), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n342), .A2(new_n811), .B1(new_n802), .B2(G97), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1052), .A2(new_n772), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(G326), .A2(new_n799), .B1(new_n802), .B2(new_n537), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n785), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n1057), .A2(G317), .B1(G311), .B2(new_n811), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n786), .B2(new_n815), .C1(new_n821), .C2(new_n518), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT112), .Z(new_n1060));
  INV_X1    g0860(.A(KEYINPUT48), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n807), .A2(G283), .B1(new_n793), .B2(G294), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT49), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n989), .B(new_n1056), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1055), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1047), .B1(new_n1069), .B2(new_n780), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n1018), .A2(new_n767), .B1(new_n1037), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1019), .A2(new_n714), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1018), .A2(new_n763), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1071), .B1(new_n1072), .B2(new_n1073), .ZN(G393));
  AND2_X1   g0874(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1019), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n715), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT114), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n1013), .A2(new_n1078), .A3(new_n1019), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1078), .B1(new_n1013), .B2(new_n1019), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1077), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n773), .A2(new_n240), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1082), .B(new_n781), .C1(new_n479), .C2(new_n206), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n768), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n1057), .A2(G311), .B1(G317), .B2(new_n809), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT52), .ZN(new_n1086));
  INV_X1    g0886(.A(G283), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n397), .B1(new_n792), .B2(new_n1087), .C1(new_n598), .C2(new_n788), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n806), .A2(new_n502), .B1(new_n812), .B2(new_n518), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n223), .A2(new_n801), .B1(new_n798), .B2(new_n786), .ZN(new_n1090));
  OR4_X1    g0890(.A1(new_n1086), .A2(new_n1088), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n821), .A2(new_n316), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n847), .B(new_n1092), .C1(G143), .C2(new_n799), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n792), .A2(new_n215), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n812), .A2(new_n290), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1094), .B(new_n1095), .C1(G77), .C2(new_n807), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1093), .A2(new_n772), .A3(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1057), .A2(G159), .B1(G150), .B2(new_n809), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT51), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1091), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1084), .B1(new_n1100), .B2(new_n780), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n1003), .B2(new_n832), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT113), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n766), .B1(new_n1013), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n1103), .B2(new_n1013), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1081), .A2(new_n1102), .A3(new_n1105), .ZN(G390));
  NOR3_X1   g0906(.A1(new_n960), .A2(new_n961), .A3(new_n943), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n895), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(KEYINPUT115), .ZN(new_n1109));
  OR3_X1    g0909(.A1(new_n893), .A2(KEYINPUT115), .A3(new_n894), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n866), .A2(new_n329), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n697), .B(new_n1113), .C1(new_n727), .C2(new_n731), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1111), .B1(new_n1114), .B2(new_n862), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1107), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n944), .B1(new_n896), .B2(new_n895), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n942), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n760), .A2(new_n867), .A3(new_n1108), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n953), .B1(new_n759), .B2(new_n950), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n954), .ZN(new_n1122));
  OAI211_X1 g0922(.A(G330), .B(new_n956), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1120), .B1(new_n1123), .B2(KEYINPUT116), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1116), .A2(new_n1118), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1123), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(KEYINPUT116), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n767), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n942), .A2(new_n777), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT54), .B(G143), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n822), .A2(new_n1133), .B1(G125), .B2(new_n799), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n792), .A2(new_n340), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT53), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1134), .B(new_n1136), .C1(new_n290), .C2(new_n801), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n397), .B1(new_n1057), .B2(G132), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(G128), .A2(new_n809), .B1(new_n811), .B2(G137), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1138), .B(new_n1139), .C1(new_n827), .C2(new_n806), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(G68), .A2(new_n802), .B1(new_n799), .B2(G294), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n479), .B2(new_n821), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n397), .B1(new_n792), .B2(new_n217), .C1(new_n1087), .C2(new_n815), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G107), .B2(new_n811), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n806), .A2(new_n221), .B1(new_n785), .B2(new_n883), .ZN(new_n1145));
  OR2_X1    g0945(.A1(new_n1145), .A2(KEYINPUT119), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(KEYINPUT119), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1144), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n1137), .A2(new_n1140), .B1(new_n1142), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n780), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n834), .B1(new_n406), .B2(new_n841), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1131), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1130), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT118), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1116), .A2(new_n1118), .A3(new_n1124), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n1115), .A2(new_n1107), .B1(new_n1117), .B2(new_n942), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1155), .B1(new_n1156), .B2(new_n1127), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n735), .B1(new_n952), .B2(new_n954), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n439), .A2(new_n1158), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n687), .B(new_n1159), .C1(new_n734), .C2(new_n440), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n758), .A2(new_n759), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1162), .A2(G330), .A3(new_n867), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n895), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1164), .A2(KEYINPUT117), .B1(new_n1158), .B2(new_n956), .ZN(new_n1165));
  AOI211_X1 g0965(.A(KEYINPUT117), .B(new_n1108), .C1(new_n760), .C2(new_n867), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n896), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n697), .B1(new_n727), .B2(new_n731), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n862), .B1(new_n1169), .B2(new_n1112), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n735), .B(new_n876), .C1(new_n952), .C2(new_n954), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1170), .B(new_n1119), .C1(new_n1171), .C2(new_n1111), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1161), .B1(new_n1168), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1154), .B1(new_n1157), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n896), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1108), .B1(new_n760), .B2(new_n867), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT117), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1123), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1176), .B1(new_n1179), .B2(new_n1166), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1160), .B1(new_n1180), .B2(new_n1172), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1127), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n1117), .A2(new_n942), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1169), .A2(new_n1112), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n862), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n1184), .A2(new_n1185), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n938), .A2(KEYINPUT109), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n927), .A2(new_n937), .A3(new_n959), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n944), .A3(new_n1188), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1186), .A2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1182), .B1(new_n1183), .B2(new_n1190), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1181), .A2(new_n1191), .A3(KEYINPUT118), .A4(new_n1155), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1175), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n715), .B1(new_n1157), .B2(new_n1174), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1153), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(G378));
  NAND2_X1  g0996(.A1(new_n344), .A2(new_n913), .ZN(new_n1197));
  XOR2_X1   g0997(.A(new_n1197), .B(KEYINPUT55), .Z(new_n1198));
  XNOR2_X1  g0998(.A(new_n368), .B(new_n1198), .ZN(new_n1199));
  XOR2_X1   g0999(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1200));
  XOR2_X1   g1000(.A(new_n1199), .B(new_n1200), .Z(new_n1201));
  OR2_X1    g1001(.A1(new_n1201), .A2(KEYINPUT122), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(KEYINPUT122), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n777), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT58), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n801), .A2(new_n372), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n1057), .A2(G107), .B1(new_n793), .B2(G77), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(new_n215), .B2(new_n806), .C1(new_n883), .C2(new_n815), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1207), .B(new_n1209), .C1(G283), .C2(new_n799), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n772), .A2(G41), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n812), .A2(new_n479), .B1(new_n788), .B2(new_n319), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT120), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1210), .A2(new_n1211), .A3(new_n1213), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n806), .A2(new_n340), .B1(new_n812), .B2(new_n858), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1057), .A2(G128), .B1(new_n793), .B2(new_n1133), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n852), .B2(new_n788), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1215), .B(new_n1217), .C1(G125), .C2(new_n809), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(KEYINPUT59), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n802), .A2(G159), .ZN(new_n1221));
  AOI211_X1 g1021(.A(G33), .B(G41), .C1(new_n799), .C2(G124), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1219), .A2(KEYINPUT59), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1206), .A2(new_n1214), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n290), .B1(G33), .B2(G41), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1225), .B1(new_n1206), .B2(new_n1214), .C1(new_n1211), .C2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n780), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n834), .B1(new_n290), .B2(new_n841), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1205), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n958), .A2(new_n962), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n964), .A2(new_n965), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1232), .A2(G330), .A3(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1201), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n966), .A2(G330), .A3(new_n1203), .A4(new_n1202), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT123), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n931), .B2(new_n945), .ZN(new_n1239));
  AND3_X1   g1039(.A1(new_n1236), .A2(new_n1237), .A3(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1239), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1241));
  OR2_X1    g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1231), .B1(new_n1242), .B2(new_n767), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT118), .B1(new_n1129), .B2(new_n1181), .ZN(new_n1244));
  AND4_X1   g1044(.A1(KEYINPUT118), .A2(new_n1181), .A3(new_n1191), .A4(new_n1155), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1161), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(KEYINPUT57), .B1(new_n1246), .B2(new_n1242), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1160), .B1(new_n1175), .B2(new_n1192), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n946), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1236), .B(new_n1237), .C1(new_n931), .C2(new_n945), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1250), .A2(KEYINPUT57), .A3(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n714), .B1(new_n1248), .B2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1243), .B1(new_n1247), .B2(new_n1253), .ZN(G375));
  INV_X1    g1054(.A(KEYINPUT125), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n834), .B1(new_n215), .B2(new_n841), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1111), .A2(new_n778), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n822), .A2(G107), .B1(G303), .B2(new_n799), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n397), .B1(new_n792), .B2(new_n479), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(G283), .B2(new_n1057), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1259), .B(new_n1261), .C1(new_n221), .C2(new_n801), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1048), .B1(new_n537), .B2(new_n811), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n598), .B2(new_n815), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1207), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n1049), .A2(G150), .B1(new_n793), .B2(G159), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n799), .A2(G128), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1057), .A2(G137), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .A4(new_n1268), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n807), .A2(G50), .B1(G132), .B2(new_n809), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n772), .B(new_n1270), .C1(new_n812), .C2(new_n1132), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n1262), .A2(new_n1264), .B1(new_n1269), .B2(new_n1271), .ZN(new_n1272));
  AOI211_X1 g1072(.A(new_n1257), .B(new_n1258), .C1(new_n780), .C2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n766), .B1(new_n1180), .B2(new_n1172), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1274), .B1(new_n1275), .B2(KEYINPUT124), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT124), .ZN(new_n1277));
  AOI211_X1 g1077(.A(new_n1277), .B(new_n766), .C1(new_n1180), .C2(new_n1172), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1255), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n767), .B1(new_n1168), .B2(new_n1173), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1277), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1275), .A2(KEYINPUT124), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1281), .A2(KEYINPUT125), .A3(new_n1282), .A4(new_n1274), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1279), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1180), .A2(new_n1160), .A3(new_n1172), .ZN(new_n1286));
  AND3_X1   g1086(.A1(new_n1174), .A2(new_n1022), .A3(new_n1286), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(G381));
  OR3_X1    g1089(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1290));
  NOR3_X1   g1090(.A1(G390), .A2(G387), .A3(new_n1290), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1291), .A2(new_n1195), .A3(new_n1288), .ZN(new_n1292));
  INV_X1    g1092(.A(G375), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1292), .A2(KEYINPUT126), .A3(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT126), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1295));
  OR2_X1    g1095(.A1(new_n1294), .A2(new_n1295), .ZN(G407));
  INV_X1    g1096(.A(G213), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(G378), .A2(G343), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1297), .B1(new_n1293), .B2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1299), .B1(new_n1294), .B2(new_n1295), .ZN(G409));
  INV_X1    g1100(.A(KEYINPUT61), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1297), .A2(G343), .ZN(new_n1302));
  OAI211_X1 g1102(.A(G378), .B(new_n1243), .C1(new_n1247), .C2(new_n1253), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1304));
  NOR3_X1   g1104(.A1(new_n1248), .A2(new_n1304), .A3(new_n1021), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1250), .A2(new_n767), .A3(new_n1251), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1230), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1195), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1302), .B1(new_n1303), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1302), .A2(G2897), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT127), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n1286), .A2(new_n1312), .A3(KEYINPUT60), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT60), .B1(new_n1286), .B2(new_n1312), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n714), .B(new_n1174), .C1(new_n1313), .C2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1284), .A2(G384), .A3(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(G384), .B1(new_n1284), .B2(new_n1315), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1311), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1284), .A2(new_n1315), .ZN(new_n1320));
  INV_X1    g1120(.A(G384), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1322), .A2(new_n1316), .A3(new_n1310), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1319), .A2(new_n1323), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1301), .B1(new_n1309), .B2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT63), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1303), .A2(new_n1308), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1302), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1327), .B1(new_n1330), .B2(new_n1332), .ZN(new_n1333));
  OR2_X1    g1133(.A1(new_n1023), .A2(new_n1035), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1334), .A2(G390), .A3(new_n1000), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(G387), .A2(new_n1081), .A3(new_n1102), .A4(new_n1105), .ZN(new_n1336));
  XNOR2_X1  g1136(.A(G393), .B(new_n839), .ZN(new_n1337));
  AND3_X1   g1137(.A1(new_n1335), .A2(new_n1336), .A3(new_n1337), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1337), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1309), .A2(KEYINPUT63), .A3(new_n1331), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1326), .A2(new_n1333), .A3(new_n1340), .A4(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT62), .ZN(new_n1343));
  AND3_X1   g1143(.A1(new_n1309), .A2(new_n1343), .A3(new_n1331), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1343), .B1(new_n1309), .B2(new_n1331), .ZN(new_n1345));
  NOR3_X1   g1145(.A1(new_n1344), .A2(new_n1325), .A3(new_n1345), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1342), .B1(new_n1346), .B2(new_n1340), .ZN(G405));
  OR2_X1    g1147(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(G375), .A2(new_n1195), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(new_n1303), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1350), .A2(new_n1331), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1332), .A2(new_n1349), .A3(new_n1303), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1351), .A2(new_n1352), .ZN(new_n1353));
  XNOR2_X1  g1153(.A(new_n1348), .B(new_n1353), .ZN(G402));
endmodule


