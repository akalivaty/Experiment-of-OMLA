//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 0 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n807, new_n809, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(G190gat), .ZN(new_n204));
  AND2_X1   g003(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT28), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT26), .ZN(new_n210));
  INV_X1    g009(.A(G169gat), .ZN(new_n211));
  INV_X1    g010(.A(G176gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n209), .B(new_n213), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT28), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n219), .B(new_n204), .C1(new_n205), .C2(new_n206), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n208), .A2(new_n217), .A3(new_n218), .A4(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n218), .A2(KEYINPUT24), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n223), .B1(G183gat), .B2(G190gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n222), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n211), .A2(new_n212), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n232));
  AOI22_X1  g031(.A1(new_n230), .A2(new_n214), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT25), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n232), .A2(G176gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT64), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n236), .A2(G169gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n211), .A2(KEYINPUT64), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n235), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n227), .A2(new_n233), .A3(new_n234), .A4(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n223), .A2(G183gat), .A3(G190gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT23), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n218), .A2(KEYINPUT24), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n241), .B(new_n242), .C1(new_n243), .C2(new_n225), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n232), .B1(G169gat), .B2(G176gat), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n245), .B1(new_n215), .B2(new_n216), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT25), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n221), .A2(new_n240), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G113gat), .B(G120gat), .ZN(new_n249));
  OAI21_X1  g048(.A(G127gat), .B1(new_n249), .B2(KEYINPUT1), .ZN(new_n250));
  INV_X1    g049(.A(G120gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G113gat), .ZN(new_n252));
  INV_X1    g051(.A(G113gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(G120gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT1), .ZN(new_n256));
  INV_X1    g055(.A(G127gat), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  AND3_X1   g057(.A1(new_n250), .A2(new_n258), .A3(G134gat), .ZN(new_n259));
  AOI21_X1  g058(.A(G134gat), .B1(new_n250), .B2(new_n258), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n248), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G134gat), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n257), .B1(new_n255), .B2(new_n256), .ZN(new_n264));
  AOI211_X1 g063(.A(KEYINPUT1), .B(G127gat), .C1(new_n252), .C2(new_n254), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n250), .A2(new_n258), .A3(G134gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n221), .A2(new_n240), .A3(new_n247), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n203), .B1(new_n262), .B2(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(G15gat), .B(G43gat), .Z(new_n272));
  XNOR2_X1  g071(.A(G71gat), .B(G99gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT33), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n271), .A2(KEYINPUT32), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n248), .A2(new_n261), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n268), .A2(new_n269), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n202), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n274), .B1(new_n279), .B2(KEYINPUT33), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT32), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  OAI211_X1 g081(.A(KEYINPUT66), .B(new_n276), .C1(new_n280), .C2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n271), .A2(KEYINPUT32), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT33), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n271), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT66), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n284), .A2(new_n286), .A3(new_n287), .A4(new_n274), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n283), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n262), .A2(new_n270), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(new_n202), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT34), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT34), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n290), .A2(new_n293), .A3(new_n202), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT67), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT67), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n292), .A2(new_n297), .A3(new_n294), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n289), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n295), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n300), .A2(new_n283), .A3(new_n297), .A4(new_n288), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G78gat), .B(G106gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n303), .B(KEYINPUT31), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n304), .B(G50gat), .ZN(new_n305));
  INV_X1    g104(.A(G22gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT2), .ZN(new_n307));
  INV_X1    g106(.A(G155gat), .ZN(new_n308));
  INV_X1    g107(.A(G162gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311));
  INV_X1    g110(.A(G148gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G141gat), .ZN(new_n313));
  INV_X1    g112(.A(G141gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G148gat), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n310), .A2(new_n311), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n311), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n313), .A2(new_n315), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n317), .B1(new_n318), .B2(new_n307), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT73), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n320), .A2(new_n308), .A3(new_n309), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT73), .B1(G155gat), .B2(G162gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n316), .B1(new_n319), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT74), .B(KEYINPUT3), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT29), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G218gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT68), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT68), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(G218gat), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT22), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(G197gat), .B(G204gat), .Z(new_n334));
  OAI21_X1  g133(.A(G211gat), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G197gat), .B(G204gat), .ZN(new_n336));
  INV_X1    g135(.A(G211gat), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n336), .A2(KEYINPUT22), .A3(new_n337), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n335), .A2(new_n329), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n329), .B1(new_n335), .B2(new_n338), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT69), .ZN(new_n341));
  NOR3_X1   g140(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n330), .A2(new_n332), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT22), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n337), .B1(new_n345), .B2(new_n336), .ZN(new_n346));
  INV_X1    g145(.A(new_n338), .ZN(new_n347));
  OAI21_X1  g146(.A(G218gat), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n335), .A2(new_n329), .A3(new_n338), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT69), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n328), .B1(new_n342), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n325), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT29), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n348), .A2(new_n352), .A3(new_n353), .A4(new_n349), .ZN(new_n354));
  INV_X1    g153(.A(G228gat), .ZN(new_n355));
  INV_X1    g154(.A(G233gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AND2_X1   g156(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT2), .B1(new_n313), .B2(new_n315), .ZN(new_n359));
  NOR3_X1   g158(.A1(new_n359), .A2(new_n323), .A3(new_n317), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT3), .B1(new_n360), .B2(new_n316), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n351), .A2(new_n358), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n348), .A2(new_n353), .A3(new_n349), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n325), .B1(new_n363), .B2(new_n326), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n339), .A2(new_n340), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n365), .A2(new_n327), .ZN(new_n366));
  OAI22_X1  g165(.A1(new_n364), .A2(new_n366), .B1(new_n355), .B2(new_n356), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n306), .B1(new_n362), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n305), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n363), .A2(new_n326), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(new_n352), .ZN(new_n372));
  INV_X1    g171(.A(new_n366), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n357), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n341), .B1(new_n339), .B2(new_n340), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n348), .A2(KEYINPUT69), .A3(new_n349), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n327), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n354), .A2(new_n357), .ZN(new_n378));
  INV_X1    g177(.A(new_n361), .ZN(new_n379));
  NOR3_X1   g178(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(G22gat), .B1(new_n374), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n362), .A2(new_n367), .A3(new_n306), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n370), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n381), .A2(new_n382), .A3(new_n369), .A4(new_n305), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n302), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT86), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(KEYINPUT76), .B(KEYINPUT5), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n266), .A2(new_n325), .A3(new_n267), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT4), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n325), .A2(new_n326), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n268), .A2(new_n395), .A3(new_n361), .ZN(new_n396));
  NAND2_X1  g195(.A1(G225gat), .A2(G233gat), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n266), .A2(new_n325), .A3(KEYINPUT4), .A4(new_n267), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n394), .A2(new_n396), .A3(new_n397), .A4(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n391), .B1(new_n399), .B2(KEYINPUT75), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n394), .A2(new_n398), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT75), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n401), .A2(new_n402), .A3(new_n397), .A4(new_n396), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n268), .A2(new_n352), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n392), .ZN(new_n405));
  INV_X1    g204(.A(new_n397), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n400), .A2(new_n403), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT79), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n409), .B1(new_n399), .B2(new_n390), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n394), .A2(new_n396), .A3(new_n398), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n411), .A2(KEYINPUT79), .A3(new_n397), .A4(new_n391), .ZN(new_n412));
  XNOR2_X1  g211(.A(G1gat), .B(G29gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(KEYINPUT78), .ZN(new_n414));
  XNOR2_X1  g213(.A(G57gat), .B(G85gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n416), .B(new_n417), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n408), .A2(new_n410), .A3(new_n412), .A4(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT6), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n408), .A2(new_n410), .A3(new_n412), .ZN(new_n422));
  INV_X1    g221(.A(new_n418), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n422), .A2(KEYINPUT6), .A3(new_n423), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n269), .A2(new_n353), .ZN(new_n427));
  INV_X1    g226(.A(G226gat), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n428), .A2(new_n356), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT71), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT72), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n269), .A2(new_n429), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n431), .A2(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n269), .A2(KEYINPUT72), .A3(new_n429), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n427), .A2(KEYINPUT71), .A3(new_n430), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n435), .A2(new_n365), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT70), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n269), .A2(KEYINPUT70), .A3(new_n429), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n431), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n375), .A2(new_n376), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n438), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT30), .ZN(new_n447));
  XNOR2_X1  g246(.A(G8gat), .B(G36gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(G64gat), .B(G92gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n448), .B(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n446), .A2(new_n447), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n446), .A2(new_n451), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n447), .B1(new_n445), .B2(new_n450), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n425), .A2(new_n426), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n302), .A2(new_n386), .A3(KEYINPUT86), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n389), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT35), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n412), .A2(new_n410), .ZN(new_n460));
  AOI211_X1 g259(.A(KEYINPUT82), .B(new_n418), .C1(new_n460), .C2(new_n408), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT82), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n462), .B1(new_n422), .B2(new_n423), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n421), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT83), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g265(.A(KEYINPUT83), .B(new_n421), .C1(new_n461), .C2(new_n463), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(new_n426), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n455), .A2(new_n452), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n470), .A2(KEYINPUT35), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n299), .A2(KEYINPUT85), .A3(new_n301), .ZN(new_n472));
  INV_X1    g271(.A(new_n386), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT85), .B1(new_n299), .B2(new_n301), .ZN(new_n474));
  NOR3_X1   g273(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n468), .A2(new_n471), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n476), .ZN(new_n477));
  OR3_X1    g276(.A1(new_n442), .A2(KEYINPUT84), .A3(new_n443), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT84), .B1(new_n442), .B2(new_n443), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n481));
  INV_X1    g280(.A(new_n365), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT37), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT37), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n438), .A2(new_n485), .A3(new_n444), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT38), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n486), .A2(new_n487), .A3(new_n450), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n484), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n486), .A2(new_n450), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n485), .B1(new_n438), .B2(new_n444), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT38), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n489), .A2(new_n453), .A3(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n466), .A2(new_n493), .A3(new_n426), .A4(new_n467), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT39), .B1(new_n405), .B2(new_n406), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT81), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n394), .A2(new_n396), .A3(new_n398), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n406), .ZN(new_n499));
  OAI211_X1 g298(.A(KEYINPUT81), .B(KEYINPUT39), .C1(new_n405), .C2(new_n406), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n499), .A2(KEYINPUT39), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(new_n418), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT40), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n504), .ZN(new_n506));
  AND4_X1   g305(.A1(new_n452), .A2(new_n455), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n461), .A2(new_n463), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n473), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n425), .A2(new_n426), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n386), .B1(new_n511), .B2(new_n469), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT36), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n302), .B(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT87), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n477), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n517), .B1(new_n477), .B2(new_n516), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT15), .ZN(new_n521));
  XOR2_X1   g320(.A(G43gat), .B(G50gat), .Z(new_n522));
  INV_X1    g321(.A(KEYINPUT89), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(G29gat), .A2(G36gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT14), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n526), .B1(G29gat), .B2(G36gat), .ZN(new_n527));
  INV_X1    g326(.A(G29gat), .ZN(new_n528));
  INV_X1    g327(.A(G36gat), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(new_n529), .A3(KEYINPUT14), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n524), .A2(new_n525), .A3(new_n527), .A4(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(new_n527), .A3(new_n525), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n522), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n521), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n532), .B1(new_n523), .B2(new_n522), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n535), .A2(KEYINPUT15), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(KEYINPUT17), .ZN(new_n538));
  XNOR2_X1  g337(.A(G15gat), .B(G22gat), .ZN(new_n539));
  INV_X1    g338(.A(G1gat), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n539), .A2(KEYINPUT16), .A3(new_n540), .ZN(new_n541));
  OAI221_X1 g340(.A(new_n541), .B1(KEYINPUT90), .B2(G8gat), .C1(new_n540), .C2(new_n539), .ZN(new_n542));
  NAND2_X1  g341(.A1(KEYINPUT90), .A2(G8gat), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n542), .B(new_n543), .Z(new_n544));
  NAND2_X1  g343(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  OR3_X1    g344(.A1(new_n544), .A2(new_n534), .A3(new_n536), .ZN(new_n546));
  NAND2_X1  g345(.A1(G229gat), .A2(G233gat), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT18), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n544), .B(new_n537), .Z(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(new_n547), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n545), .A2(KEYINPUT18), .A3(new_n546), .A4(new_n547), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n550), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G113gat), .B(G141gat), .ZN(new_n557));
  INV_X1    g356(.A(G197gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(KEYINPUT11), .B(G169gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT88), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT12), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n556), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n556), .A2(new_n563), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n565), .A2(KEYINPUT92), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT92), .ZN(new_n567));
  NOR3_X1   g366(.A1(new_n556), .A2(new_n567), .A3(new_n563), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n564), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G99gat), .B(G106gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT95), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT96), .ZN(new_n572));
  OR2_X1    g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n572), .ZN(new_n574));
  NAND2_X1  g373(.A1(G99gat), .A2(G106gat), .ZN(new_n575));
  INV_X1    g374(.A(G85gat), .ZN(new_n576));
  INV_X1    g375(.A(G92gat), .ZN(new_n577));
  AOI22_X1  g376(.A1(KEYINPUT8), .A2(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT94), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G85gat), .A2(G92gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT7), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n573), .A2(new_n574), .A3(new_n580), .A4(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n580), .A2(new_n582), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n584), .A2(new_n572), .A3(new_n571), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT97), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(new_n538), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n537), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT41), .ZN(new_n591));
  NAND2_X1  g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n589), .B(new_n590), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G190gat), .B(G218gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G134gat), .B(G162gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n592), .A2(new_n591), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n595), .A2(new_n599), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT21), .ZN(new_n604));
  XOR2_X1   g403(.A(G71gat), .B(G78gat), .Z(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G57gat), .B(G64gat), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n605), .B1(new_n607), .B2(new_n608), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n544), .B1(new_n604), .B2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(G183gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(G127gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n612), .A2(new_n604), .ZN(new_n616));
  XNOR2_X1  g415(.A(KEYINPUT93), .B(G211gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n618), .B(new_n619), .Z(new_n620));
  XNOR2_X1  g419(.A(new_n615), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(G155gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n621), .B(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT100), .ZN(new_n625));
  INV_X1    g424(.A(new_n612), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n587), .A2(KEYINPUT10), .A3(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT10), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n629), .A2(KEYINPUT99), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n629), .A2(KEYINPUT99), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT98), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n612), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n612), .A2(new_n632), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n586), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n583), .A2(KEYINPUT98), .A3(new_n626), .A4(new_n585), .ZN(new_n637));
  AOI211_X1 g436(.A(new_n630), .B(new_n631), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n625), .B1(new_n628), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G230gat), .A2(G233gat), .ZN(new_n640));
  INV_X1    g439(.A(new_n638), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n641), .A2(KEYINPUT100), .A3(new_n627), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n639), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n636), .A2(new_n637), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n644), .A2(new_n640), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G120gat), .B(G148gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(G176gat), .B(G204gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n643), .A2(new_n646), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n640), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n652), .B1(new_n641), .B2(new_n627), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n649), .B1(new_n653), .B2(new_n645), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n603), .A2(new_n624), .A3(new_n655), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n520), .A2(KEYINPUT101), .A3(new_n569), .A4(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n477), .A2(new_n516), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT87), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n477), .A2(new_n516), .A3(new_n517), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n659), .A2(new_n660), .A3(new_n569), .A4(new_n656), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT101), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n657), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(new_n511), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(new_n540), .ZN(G1324gat));
  OAI21_X1  g466(.A(G8gat), .B1(new_n665), .B2(new_n469), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n469), .B1(new_n657), .B2(new_n663), .ZN(new_n669));
  OR2_X1    g468(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n670));
  NAND2_X1  g469(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n669), .A2(KEYINPUT42), .A3(new_n670), .A4(new_n671), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(KEYINPUT102), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT102), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n674), .A2(new_n678), .A3(new_n675), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n673), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(KEYINPUT103), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n673), .A2(new_n677), .A3(new_n682), .A4(new_n679), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(G1325gat));
  INV_X1    g483(.A(G15gat), .ZN(new_n685));
  INV_X1    g484(.A(new_n514), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n665), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n472), .A2(new_n474), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n685), .B1(new_n665), .B2(new_n689), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n690), .A2(KEYINPUT104), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(KEYINPUT104), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n687), .B1(new_n691), .B2(new_n692), .ZN(G1326gat));
  NAND2_X1  g492(.A1(new_n664), .A2(new_n473), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT43), .B(G22gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1327gat));
  INV_X1    g495(.A(new_n624), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n697), .A2(new_n655), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n520), .A2(new_n569), .A3(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n603), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n511), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(new_n528), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT45), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n518), .A2(new_n519), .A3(new_n700), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706));
  OAI21_X1  g505(.A(KEYINPUT106), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n659), .A2(new_n660), .A3(new_n603), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT106), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n708), .A2(new_n709), .A3(KEYINPUT44), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT107), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n512), .A2(new_n711), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n456), .A2(KEYINPUT107), .A3(new_n386), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n510), .B(new_n686), .C1(new_n712), .C2(new_n713), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n459), .A2(new_n476), .A3(KEYINPUT108), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT108), .B1(new_n459), .B2(new_n476), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n718), .B1(new_n601), .B2(new_n602), .ZN(new_n719));
  INV_X1    g518(.A(new_n602), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n720), .A2(KEYINPUT109), .A3(new_n600), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n717), .A2(new_n706), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(KEYINPUT110), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT110), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n717), .A2(new_n725), .A3(new_n706), .A4(new_n722), .ZN(new_n726));
  AOI22_X1  g525(.A1(new_n707), .A2(new_n710), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n698), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n565), .B(KEYINPUT92), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n729), .A2(KEYINPUT105), .A3(new_n564), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n569), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n728), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n727), .A2(new_n511), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n704), .B1(new_n528), .B2(new_n737), .ZN(G1328gat));
  AND3_X1   g537(.A1(new_n708), .A2(new_n709), .A3(KEYINPUT44), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n709), .B1(new_n708), .B2(KEYINPUT44), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n468), .A2(new_n471), .A3(new_n475), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT35), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n302), .A2(new_n386), .A3(KEYINPUT86), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT86), .B1(new_n302), .B2(new_n386), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n743), .B1(new_n746), .B2(new_n456), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n741), .B1(new_n742), .B2(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n459), .A2(new_n476), .A3(KEYINPUT108), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(KEYINPUT44), .B1(new_n750), .B2(new_n714), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n725), .B1(new_n751), .B2(new_n722), .ZN(new_n752));
  INV_X1    g551(.A(new_n726), .ZN(new_n753));
  OAI22_X1  g552(.A1(new_n739), .A2(new_n740), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n754), .A2(new_n470), .A3(new_n735), .ZN(new_n755));
  OR2_X1    g554(.A1(new_n755), .A2(KEYINPUT112), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(KEYINPUT112), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n756), .A2(new_n757), .A3(G36gat), .ZN(new_n758));
  NAND2_X1  g557(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n701), .A2(new_n529), .A3(new_n470), .A4(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n758), .A2(new_n762), .ZN(G1329gat));
  NAND2_X1  g562(.A1(new_n514), .A2(G43gat), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n727), .A2(new_n736), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(G43gat), .B1(new_n701), .B2(new_n688), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT113), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT47), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(KEYINPUT113), .A2(KEYINPUT47), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n767), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n770), .B1(new_n767), .B2(new_n771), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(G1330gat));
  NAND3_X1  g573(.A1(new_n754), .A2(new_n473), .A3(new_n735), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT115), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n754), .A2(KEYINPUT115), .A3(new_n473), .A4(new_n735), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n777), .A2(G50gat), .A3(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(G50gat), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n701), .A2(new_n780), .A3(new_n473), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n779), .A2(KEYINPUT48), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT114), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n727), .A2(new_n386), .A3(new_n736), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n781), .B1(new_n784), .B2(new_n780), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT48), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n783), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n781), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n788), .B1(new_n775), .B2(G50gat), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n789), .A2(KEYINPUT114), .A3(KEYINPUT48), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n782), .B1(new_n787), .B2(new_n790), .ZN(G1331gat));
  AND3_X1   g590(.A1(new_n717), .A2(new_n697), .A3(new_n700), .ZN(new_n792));
  INV_X1    g591(.A(new_n655), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n733), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  XOR2_X1   g595(.A(new_n511), .B(KEYINPUT116), .Z(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g598(.A1(new_n795), .A2(new_n469), .ZN(new_n800));
  NOR2_X1   g599(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n801));
  AND2_X1   g600(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n803), .B1(new_n800), .B2(new_n801), .ZN(G1333gat));
  OAI21_X1  g603(.A(G71gat), .B1(new_n795), .B2(new_n686), .ZN(new_n805));
  OR2_X1    g604(.A1(new_n689), .A2(G71gat), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n805), .B1(new_n795), .B2(new_n806), .ZN(new_n807));
  XOR2_X1   g606(.A(new_n807), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g607(.A1(new_n796), .A2(new_n473), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g609(.A1(new_n697), .A2(new_n733), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n754), .A2(new_n655), .A3(new_n811), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n812), .A2(new_n576), .A3(new_n511), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n717), .A2(new_n603), .A3(new_n811), .ZN(new_n814));
  OR2_X1    g613(.A1(new_n814), .A2(KEYINPUT51), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(KEYINPUT51), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n815), .A2(new_n655), .A3(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(G85gat), .B1(new_n818), .B2(new_n702), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n813), .A2(new_n819), .ZN(G1336gat));
  NOR2_X1   g619(.A1(new_n817), .A2(G92gat), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT117), .B1(new_n821), .B2(new_n470), .ZN(new_n822));
  INV_X1    g621(.A(new_n811), .ZN(new_n823));
  NOR4_X1   g622(.A1(new_n727), .A2(new_n469), .A3(new_n793), .A4(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n822), .B1(new_n577), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(KEYINPUT52), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n822), .B(new_n827), .C1(new_n577), .C2(new_n824), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(G1337gat));
  OAI21_X1  g628(.A(G99gat), .B1(new_n812), .B2(new_n686), .ZN(new_n830));
  OR3_X1    g629(.A1(new_n817), .A2(G99gat), .A3(new_n689), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(G1338gat));
  INV_X1    g631(.A(G106gat), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n833), .B1(new_n817), .B2(new_n386), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n754), .A2(new_n473), .A3(new_n655), .A4(new_n811), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n835), .B1(new_n837), .B2(KEYINPUT118), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n833), .B1(new_n836), .B2(KEYINPUT118), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n838), .A2(new_n840), .A3(KEYINPUT53), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n834), .B1(new_n836), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n842), .B1(new_n844), .B2(new_n839), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n841), .A2(new_n845), .ZN(G1339gat));
  INV_X1    g645(.A(new_n797), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n641), .A2(new_n652), .A3(new_n627), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n643), .A2(new_n848), .A3(KEYINPUT54), .ZN(new_n849));
  XNOR2_X1  g648(.A(KEYINPUT119), .B(KEYINPUT54), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n653), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n849), .A2(KEYINPUT55), .A3(new_n649), .A4(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n849), .A2(new_n649), .A3(new_n851), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT55), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n733), .A2(new_n651), .A3(new_n852), .A4(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n551), .A2(new_n553), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n547), .B1(new_n545), .B2(new_n546), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n561), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  XOR2_X1   g658(.A(new_n859), .B(KEYINPUT120), .Z(new_n860));
  AND2_X1   g659(.A1(new_n729), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n655), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n722), .B1(new_n856), .B2(new_n862), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n719), .A2(new_n721), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n861), .A2(new_n651), .A3(new_n852), .A4(new_n855), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n624), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n656), .A2(new_n734), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n847), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n869), .A2(new_n746), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n870), .A2(new_n469), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(new_n253), .A3(new_n733), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n473), .B1(new_n867), .B2(new_n868), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n511), .A2(new_n470), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n873), .A2(new_n688), .A3(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n569), .ZN(new_n876));
  OAI21_X1  g675(.A(G113gat), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n872), .A2(new_n877), .ZN(G1340gat));
  NAND3_X1  g677(.A1(new_n871), .A2(new_n251), .A3(new_n655), .ZN(new_n879));
  OAI21_X1  g678(.A(G120gat), .B1(new_n875), .B2(new_n793), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(G1341gat));
  NAND3_X1  g680(.A1(new_n871), .A2(new_n257), .A3(new_n697), .ZN(new_n882));
  OAI21_X1  g681(.A(G127gat), .B1(new_n875), .B2(new_n624), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(G1342gat));
  NOR2_X1   g683(.A1(new_n700), .A2(new_n470), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n870), .A2(new_n263), .A3(new_n885), .ZN(new_n886));
  XOR2_X1   g685(.A(new_n886), .B(KEYINPUT56), .Z(new_n887));
  OAI21_X1  g686(.A(G134gat), .B1(new_n875), .B2(new_n700), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(G1343gat));
  NAND2_X1  g688(.A1(new_n686), .A2(new_n874), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n867), .A2(new_n868), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT57), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(new_n893), .A3(new_n473), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT121), .B1(new_n855), .B2(new_n852), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n896), .B1(new_n853), .B2(new_n854), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n569), .A3(new_n651), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n603), .B1(new_n899), .B2(new_n862), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n624), .B1(new_n900), .B2(new_n866), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n386), .B1(new_n901), .B2(new_n868), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n891), .B(new_n894), .C1(new_n902), .C2(new_n893), .ZN(new_n903));
  OAI21_X1  g702(.A(G141gat), .B1(new_n903), .B2(new_n876), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT58), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT122), .B1(new_n514), .B2(new_n386), .ZN(new_n906));
  OR3_X1    g705(.A1(new_n514), .A2(KEYINPUT122), .A3(new_n386), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n869), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(KEYINPUT123), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n876), .A2(G141gat), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n869), .A2(new_n911), .A3(new_n906), .A4(new_n907), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n909), .A2(new_n469), .A3(new_n910), .A4(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n904), .A2(new_n905), .A3(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n651), .ZN(new_n915));
  NOR4_X1   g714(.A1(new_n895), .A2(new_n876), .A3(new_n915), .A4(new_n897), .ZN(new_n916));
  INV_X1    g715(.A(new_n862), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n700), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(new_n866), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n697), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n868), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n473), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n890), .B1(new_n922), .B2(KEYINPUT57), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n733), .A3(new_n894), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n908), .A2(new_n470), .ZN(new_n925));
  AOI22_X1  g724(.A1(new_n924), .A2(G141gat), .B1(new_n910), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n914), .B1(new_n926), .B2(new_n905), .ZN(G1344gat));
  NAND2_X1  g726(.A1(new_n473), .A2(new_n893), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n865), .A2(new_n700), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n624), .B1(new_n900), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n656), .A2(new_n876), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n893), .B1(new_n892), .B2(new_n473), .ZN(new_n933));
  NOR4_X1   g732(.A1(new_n932), .A2(new_n933), .A3(new_n793), .A4(new_n890), .ZN(new_n934));
  OAI21_X1  g733(.A(KEYINPUT59), .B1(new_n934), .B2(new_n312), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT59), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n936), .B(G148gat), .C1(new_n903), .C2(new_n793), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n909), .A2(new_n912), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n939), .A2(new_n470), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n940), .A2(new_n312), .A3(new_n655), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n938), .A2(new_n941), .ZN(G1345gat));
  INV_X1    g741(.A(new_n903), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n697), .A2(G155gat), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT124), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n909), .A2(new_n469), .A3(new_n697), .A4(new_n912), .ZN(new_n946));
  AOI22_X1  g745(.A1(new_n943), .A2(new_n945), .B1(new_n946), .B2(new_n308), .ZN(G1346gat));
  OAI21_X1  g746(.A(G162gat), .B1(new_n903), .B2(new_n864), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n885), .A2(new_n309), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(new_n939), .B2(new_n949), .ZN(G1347gat));
  AOI21_X1  g749(.A(new_n702), .B1(new_n867), .B2(new_n868), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n951), .A2(new_n470), .A3(new_n746), .ZN(new_n952));
  OAI211_X1 g751(.A(new_n952), .B(new_n733), .C1(new_n237), .C2(new_n238), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n797), .A2(new_n469), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g754(.A(KEYINPUT125), .B1(new_n955), .B2(new_n689), .ZN(new_n956));
  OR3_X1    g755(.A1(new_n955), .A2(KEYINPUT125), .A3(new_n689), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n873), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(G169gat), .B1(new_n958), .B2(new_n876), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n953), .A2(new_n959), .ZN(G1348gat));
  AOI21_X1  g759(.A(G176gat), .B1(new_n952), .B2(new_n655), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n958), .A2(new_n212), .A3(new_n793), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n961), .A2(new_n962), .ZN(G1349gat));
  OAI21_X1  g762(.A(G183gat), .B1(new_n958), .B2(new_n624), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n952), .B1(new_n206), .B2(new_n205), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n965), .B2(new_n624), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g766(.A1(new_n952), .A2(new_n204), .A3(new_n722), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT61), .ZN(new_n969));
  INV_X1    g768(.A(new_n958), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(new_n603), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n969), .B1(new_n971), .B2(G190gat), .ZN(new_n972));
  AOI211_X1 g771(.A(KEYINPUT61), .B(new_n204), .C1(new_n970), .C2(new_n603), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n968), .B1(new_n972), .B2(new_n973), .ZN(G1351gat));
  NOR2_X1   g773(.A1(new_n514), .A2(new_n386), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n951), .A2(new_n470), .A3(new_n975), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n976), .A2(new_n558), .A3(new_n733), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n955), .A2(new_n514), .ZN(new_n978));
  INV_X1    g777(.A(new_n978), .ZN(new_n979));
  NOR4_X1   g778(.A1(new_n932), .A2(new_n933), .A3(new_n876), .A4(new_n979), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n977), .B1(new_n980), .B2(new_n558), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(KEYINPUT126), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT126), .ZN(new_n983));
  OAI211_X1 g782(.A(new_n977), .B(new_n983), .C1(new_n980), .C2(new_n558), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n982), .A2(new_n984), .ZN(G1352gat));
  INV_X1    g784(.A(G204gat), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n976), .A2(new_n986), .A3(new_n655), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT62), .ZN(new_n988));
  OR2_X1    g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n987), .A2(new_n988), .ZN(new_n990));
  NOR4_X1   g789(.A1(new_n932), .A2(new_n933), .A3(new_n793), .A4(new_n979), .ZN(new_n991));
  OAI211_X1 g790(.A(new_n989), .B(new_n990), .C1(new_n986), .C2(new_n991), .ZN(G1353gat));
  NOR4_X1   g791(.A1(new_n932), .A2(new_n933), .A3(new_n624), .A4(new_n979), .ZN(new_n993));
  INV_X1    g792(.A(new_n993), .ZN(new_n994));
  OR2_X1    g793(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n995));
  NAND2_X1  g794(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n996));
  NAND4_X1  g795(.A1(new_n994), .A2(G211gat), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  OAI211_X1 g796(.A(KEYINPUT127), .B(KEYINPUT63), .C1(new_n993), .C2(new_n337), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n976), .A2(new_n337), .A3(new_n697), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(G1354gat));
  AOI21_X1  g799(.A(G218gat), .B1(new_n976), .B2(new_n722), .ZN(new_n1001));
  NOR3_X1   g800(.A1(new_n932), .A2(new_n933), .A3(new_n979), .ZN(new_n1002));
  NOR2_X1   g801(.A1(new_n700), .A2(new_n343), .ZN(new_n1003));
  AOI21_X1  g802(.A(new_n1001), .B1(new_n1002), .B2(new_n1003), .ZN(G1355gat));
endmodule


