//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 0 1 1 1 0 0 0 1 1 0 0 1 0 0 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1294, new_n1295, new_n1296, new_n1297,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n207), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT1), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n207), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT0), .Z(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(new_n201), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(G50), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  AOI211_X1 g0024(.A(new_n215), .B(new_n218), .C1(new_n221), .C2(new_n224), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(KEYINPUT2), .B(G226), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G264), .B(G270), .Z(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XNOR2_X1  g0034(.A(G87), .B(G97), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT65), .ZN(new_n236));
  XOR2_X1   g0036(.A(G107), .B(G116), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G351));
  INV_X1    g0042(.A(G274), .ZN(new_n243));
  AND2_X1   g0043(.A1(G1), .A2(G13), .ZN(new_n244));
  NAND2_X1  g0044(.A1(G33), .A2(G41), .ZN(new_n245));
  AOI21_X1  g0045(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G41), .ZN(new_n247));
  INV_X1    g0047(.A(G45), .ZN(new_n248));
  AOI21_X1  g0048(.A(G1), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(new_n249), .ZN(new_n253));
  AND2_X1   g0053(.A1(new_n253), .A2(G226), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n259), .A2(new_n262), .A3(G222), .ZN(new_n263));
  INV_X1    g0063(.A(G77), .ZN(new_n264));
  INV_X1    g0064(.A(G1698), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n265), .B1(new_n257), .B2(new_n258), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  XOR2_X1   g0067(.A(KEYINPUT67), .B(G223), .Z(new_n268));
  OAI221_X1 g0068(.A(new_n263), .B1(new_n264), .B2(new_n259), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  AOI211_X1 g0069(.A(new_n251), .B(new_n254), .C1(new_n269), .C2(new_n252), .ZN(new_n270));
  NOR2_X1   g0070(.A1(G20), .A2(G33), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT8), .ZN(new_n273));
  INV_X1    g0073(.A(G58), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT68), .B(G58), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n275), .B1(new_n276), .B2(new_n273), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n220), .A2(G33), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n272), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n219), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G1), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n281), .B1(new_n283), .B2(G20), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G50), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n283), .A2(G13), .A3(G20), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n285), .B1(G50), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n282), .A2(new_n287), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n270), .A2(G190), .B1(new_n288), .B2(KEYINPUT9), .ZN(new_n289));
  INV_X1    g0089(.A(G200), .ZN(new_n290));
  OAI221_X1 g0090(.A(new_n289), .B1(KEYINPUT9), .B2(new_n288), .C1(new_n290), .C2(new_n270), .ZN(new_n291));
  XNOR2_X1  g0091(.A(new_n291), .B(KEYINPUT10), .ZN(new_n292));
  OR2_X1    g0092(.A1(new_n270), .A2(G169), .ZN(new_n293));
  INV_X1    g0093(.A(new_n288), .ZN(new_n294));
  INV_X1    g0094(.A(G179), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n270), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n293), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  AND2_X1   g0098(.A1(KEYINPUT3), .A2(G33), .ZN(new_n299));
  NOR2_X1   g0099(.A1(KEYINPUT3), .A2(G33), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n262), .A2(G226), .ZN(new_n302));
  NAND2_X1  g0102(.A1(G232), .A2(G1698), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(G33), .A2(G97), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n252), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT69), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n250), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n246), .A2(KEYINPUT69), .A3(new_n249), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n309), .A2(new_n310), .B1(G238), .B2(new_n253), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT13), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT13), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n307), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n313), .A2(G179), .A3(new_n315), .ZN(new_n316));
  AND3_X1   g0116(.A1(new_n307), .A2(new_n311), .A3(new_n314), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n314), .B1(new_n307), .B2(new_n311), .ZN(new_n318));
  OAI21_X1  g0118(.A(G169), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(KEYINPUT72), .A2(KEYINPUT14), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n316), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n313), .A2(new_n315), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n320), .B1(new_n323), .B2(G169), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT73), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n319), .A2(new_n321), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n323), .A2(G169), .A3(new_n320), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT73), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n326), .A2(new_n327), .A3(new_n328), .A4(new_n316), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT70), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n286), .A2(G68), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n331), .B1(new_n333), .B2(KEYINPUT71), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n334), .A2(KEYINPUT12), .B1(G68), .B2(new_n284), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT12), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n336), .B1(new_n332), .B2(KEYINPUT70), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n335), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n271), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(new_n202), .ZN(new_n340));
  OAI22_X1  g0140(.A1(new_n278), .A2(new_n264), .B1(new_n220), .B2(G68), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n281), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  XOR2_X1   g0142(.A(new_n342), .B(KEYINPUT11), .Z(new_n343));
  NOR2_X1   g0143(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n330), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n323), .A2(G200), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n313), .A2(G190), .A3(new_n315), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n347), .A2(new_n344), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G159), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n339), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G68), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n222), .B1(new_n276), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n352), .B1(new_n354), .B2(G20), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n257), .A2(KEYINPUT7), .A3(new_n220), .A4(new_n258), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT74), .B1(new_n299), .B2(new_n300), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT74), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n257), .A2(new_n359), .A3(new_n258), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n358), .A2(new_n360), .A3(new_n220), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT7), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n357), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI211_X1 g0163(.A(KEYINPUT16), .B(new_n355), .C1(new_n363), .C2(new_n353), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT16), .ZN(new_n365));
  INV_X1    g0165(.A(new_n352), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n274), .A2(KEYINPUT68), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT68), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G58), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n201), .B1(new_n370), .B2(G68), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n366), .B1(new_n371), .B2(new_n220), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n257), .A2(new_n220), .A3(new_n258), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n362), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n353), .B1(new_n374), .B2(new_n356), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n365), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n364), .A2(new_n281), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n277), .A2(new_n286), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(new_n284), .B2(new_n277), .ZN(new_n379));
  OAI211_X1 g0179(.A(G226), .B(G1698), .C1(new_n299), .C2(new_n300), .ZN(new_n380));
  NAND2_X1  g0180(.A1(G33), .A2(G87), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT66), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n265), .ZN(new_n383));
  NAND2_X1  g0183(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n383), .B(new_n384), .C1(new_n299), .C2(new_n300), .ZN(new_n385));
  INV_X1    g0185(.A(G223), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n380), .B(new_n381), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n252), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT77), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n244), .A2(new_n245), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n283), .B1(G41), .B2(G45), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(G232), .A3(new_n391), .ZN(new_n392));
  AND2_X1   g0192(.A1(KEYINPUT76), .A2(G190), .ZN(new_n393));
  NOR2_X1   g0193(.A1(KEYINPUT76), .A2(G190), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AND3_X1   g0195(.A1(new_n250), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n388), .A2(new_n389), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n250), .A2(new_n392), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n398), .B1(new_n387), .B2(new_n252), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n397), .B1(G200), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n389), .B1(new_n388), .B2(new_n396), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n377), .B(new_n379), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT17), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n379), .ZN(new_n405));
  INV_X1    g0205(.A(new_n281), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n374), .A2(new_n356), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G68), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n355), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n406), .B1(new_n409), .B2(new_n365), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n405), .B1(new_n410), .B2(new_n364), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n388), .A2(new_n250), .A3(new_n392), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n290), .ZN(new_n413));
  INV_X1    g0213(.A(new_n401), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(new_n414), .A3(new_n397), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n411), .A2(new_n415), .A3(KEYINPUT17), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n404), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n376), .A2(new_n281), .ZN(new_n418));
  OAI211_X1 g0218(.A(KEYINPUT16), .B(new_n366), .C1(new_n371), .C2(new_n220), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n361), .A2(new_n362), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n356), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n419), .B1(new_n421), .B2(G68), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n379), .B1(new_n418), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n399), .A2(G179), .ZN(new_n424));
  INV_X1    g0224(.A(G169), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n424), .B1(new_n425), .B2(new_n399), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n423), .A2(KEYINPUT18), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT75), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n423), .A2(new_n426), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT18), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n430), .A2(new_n428), .A3(new_n431), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n417), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n284), .A2(G77), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(G77), .B2(new_n286), .ZN(new_n438));
  XOR2_X1   g0238(.A(KEYINPUT8), .B(G58), .Z(new_n439));
  AOI22_X1  g0239(.A1(new_n439), .A2(new_n271), .B1(G20), .B2(G77), .ZN(new_n440));
  XNOR2_X1  g0240(.A(KEYINPUT15), .B(G87), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n440), .B1(new_n278), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n438), .B1(new_n281), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n301), .A2(G107), .ZN(new_n445));
  INV_X1    g0245(.A(G238), .ZN(new_n446));
  OAI221_X1 g0246(.A(new_n445), .B1(new_n385), .B2(new_n227), .C1(new_n267), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n252), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n251), .B1(G244), .B2(new_n253), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n444), .B1(new_n451), .B2(G169), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n450), .A2(G179), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G190), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n443), .B1(new_n450), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n456), .B1(G200), .B2(new_n450), .ZN(new_n457));
  OR2_X1    g0257(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  NOR4_X1   g0258(.A1(new_n298), .A2(new_n350), .A3(new_n436), .A4(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT89), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n266), .A2(G264), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n259), .A2(new_n262), .A3(G257), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n301), .A2(G303), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n252), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n283), .B(G45), .C1(new_n247), .C2(KEYINPUT5), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT81), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n248), .A2(G1), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT81), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT5), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G41), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n469), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n247), .A2(KEYINPUT5), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n468), .A2(new_n473), .A3(new_n474), .A4(new_n246), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n469), .A2(new_n474), .A3(new_n472), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n476), .A2(G270), .A3(new_n390), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n475), .A2(KEYINPUT87), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(KEYINPUT87), .B1(new_n475), .B2(new_n477), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n466), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT88), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT20), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G283), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n220), .ZN(new_n484));
  INV_X1    g0284(.A(G97), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT78), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT78), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G97), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n484), .B1(new_n489), .B2(new_n256), .ZN(new_n490));
  INV_X1    g0290(.A(G116), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n280), .A2(new_n219), .B1(G20), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n482), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(G33), .B1(new_n486), .B2(new_n488), .ZN(new_n495));
  OAI211_X1 g0295(.A(KEYINPUT20), .B(new_n492), .C1(new_n495), .C2(new_n484), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(G13), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n498), .A2(G1), .ZN(new_n499));
  AOI21_X1  g0299(.A(G116), .B1(new_n499), .B2(G20), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n283), .A2(G33), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n286), .A2(new_n501), .A3(new_n219), .A4(new_n280), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n500), .B1(G116), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n481), .B1(new_n497), .B2(new_n504), .ZN(new_n505));
  AOI211_X1 g0305(.A(KEYINPUT88), .B(new_n503), .C1(new_n494), .C2(new_n496), .ZN(new_n506));
  OAI211_X1 g0306(.A(G169), .B(new_n480), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT21), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n461), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n480), .A2(G169), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n497), .A2(new_n504), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT88), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n497), .A2(new_n481), .A3(new_n504), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n510), .A2(new_n514), .A3(KEYINPUT89), .A4(KEYINPUT21), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n509), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT90), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n505), .A2(new_n506), .ZN(new_n518));
  OAI211_X1 g0318(.A(G179), .B(new_n466), .C1(new_n478), .C2(new_n479), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n519), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n514), .A2(KEYINPUT90), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n516), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT91), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT91), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n516), .A2(new_n526), .A3(new_n523), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n507), .A2(new_n508), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n480), .A2(G200), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n518), .B(new_n529), .C1(new_n480), .C2(new_n395), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n525), .A2(new_n527), .A3(new_n528), .A4(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n339), .A2(new_n264), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT6), .ZN(new_n533));
  AND2_X1   g0333(.A1(G97), .A2(G107), .ZN(new_n534));
  NOR2_X1   g0334(.A1(G97), .A2(G107), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  XNOR2_X1  g0336(.A(KEYINPUT78), .B(G97), .ZN(new_n537));
  INV_X1    g0337(.A(G107), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT6), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n536), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n532), .B1(new_n540), .B2(G20), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n538), .B1(new_n374), .B2(new_n356), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT79), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AOI211_X1 g0344(.A(KEYINPUT79), .B(new_n538), .C1(new_n374), .C2(new_n356), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n281), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n286), .A2(G97), .ZN(new_n547));
  INV_X1    g0347(.A(new_n502), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n547), .B1(new_n548), .B2(G97), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT84), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n546), .A2(KEYINPUT84), .A3(new_n549), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n471), .A2(G41), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n390), .B(G257), .C1(new_n467), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(KEYINPUT82), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT82), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n476), .A2(new_n558), .A3(G257), .A4(new_n390), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n475), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT83), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n259), .A2(new_n262), .A3(G244), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT80), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT4), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n266), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n565), .B1(new_n563), .B2(new_n564), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n252), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT83), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n560), .A2(new_n571), .A3(new_n475), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n562), .A2(new_n570), .A3(G179), .A4(new_n572), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n562), .A2(new_n572), .A3(new_n570), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n573), .B1(new_n574), .B2(new_n425), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n554), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n259), .A2(new_n220), .A3(G87), .ZN(new_n577));
  XNOR2_X1  g0377(.A(new_n577), .B(KEYINPUT22), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT24), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n256), .A2(new_n491), .A3(G20), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT23), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n220), .B2(G107), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n538), .A2(KEYINPUT23), .A3(G20), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n580), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n578), .A2(new_n579), .A3(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n579), .B1(new_n578), .B2(new_n584), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n281), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n259), .A2(G257), .A3(G1698), .ZN(new_n589));
  NAND2_X1  g0389(.A1(G33), .A2(G294), .ZN(new_n590));
  INV_X1    g0390(.A(G250), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n589), .B(new_n590), .C1(new_n591), .C2(new_n385), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n476), .A2(new_n390), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n592), .A2(new_n252), .B1(G264), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n594), .A2(G190), .A3(new_n475), .ZN(new_n595));
  INV_X1    g0395(.A(new_n286), .ZN(new_n596));
  AOI21_X1  g0396(.A(KEYINPUT25), .B1(new_n596), .B2(new_n538), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n596), .A2(KEYINPUT25), .A3(new_n538), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n598), .A2(new_n599), .B1(G107), .B2(new_n548), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n594), .A2(new_n475), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(G200), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n588), .A2(new_n595), .A3(new_n600), .A4(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n562), .A2(new_n572), .A3(new_n570), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n550), .B1(G200), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n574), .A2(G190), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n576), .A2(new_n603), .A3(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n601), .A2(G179), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n609), .B1(new_n425), .B2(new_n601), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n588), .A2(new_n600), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n385), .A2(new_n446), .ZN(new_n613));
  NAND2_X1  g0413(.A1(G244), .A2(G1698), .ZN(new_n614));
  OAI22_X1  g0414(.A1(new_n301), .A2(new_n614), .B1(new_n256), .B2(new_n491), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n252), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n469), .A2(new_n243), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n591), .B1(new_n248), .B2(G1), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n617), .A2(new_n390), .A3(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n616), .A2(KEYINPUT85), .A3(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT85), .ZN(new_n621));
  INV_X1    g0421(.A(new_n614), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n259), .A2(new_n622), .B1(G33), .B2(G116), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n259), .A2(new_n262), .A3(G238), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n390), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n619), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n621), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n620), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(G200), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n620), .A2(new_n627), .A3(G190), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT19), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n220), .B1(new_n305), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(G87), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n538), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n632), .B1(new_n489), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n631), .B1(new_n537), .B2(new_n278), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n259), .A2(new_n220), .A3(G68), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n441), .ZN(new_n639));
  OAI22_X1  g0439(.A1(new_n638), .A2(new_n406), .B1(new_n286), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n502), .A2(new_n633), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n629), .A2(new_n630), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n620), .A2(new_n627), .A3(new_n295), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(KEYINPUT86), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n628), .A2(new_n425), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n502), .A2(new_n441), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n640), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT86), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n620), .A2(new_n627), .A3(new_n649), .A4(new_n295), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n645), .A2(new_n646), .A3(new_n648), .A4(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n612), .A2(new_n643), .A3(new_n651), .ZN(new_n652));
  NOR4_X1   g0452(.A1(new_n460), .A2(new_n531), .A3(new_n608), .A4(new_n652), .ZN(new_n653));
  XOR2_X1   g0453(.A(new_n653), .B(KEYINPUT92), .Z(G372));
  INV_X1    g0454(.A(new_n297), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n432), .A2(new_n427), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n344), .B1(new_n325), .B2(new_n329), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n657), .B1(new_n349), .B2(new_n454), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n656), .B1(new_n658), .B2(new_n417), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n655), .B1(new_n659), .B2(new_n292), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n563), .A2(new_n564), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(KEYINPUT4), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n662), .A2(new_n566), .A3(new_n567), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n252), .A2(new_n663), .B1(new_n561), .B2(KEYINPUT83), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n425), .B1(new_n664), .B2(new_n572), .ZN(new_n665));
  INV_X1    g0465(.A(new_n573), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n550), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT93), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT26), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n425), .B1(new_n625), .B2(new_n626), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n648), .A2(new_n644), .A3(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n625), .A2(new_n626), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n642), .B(new_n630), .C1(new_n290), .C2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n575), .A2(KEYINPUT93), .A3(new_n550), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n669), .A2(new_n670), .A3(new_n676), .A4(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n672), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n554), .A2(new_n575), .A3(new_n643), .A4(new_n651), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n679), .B1(new_n680), .B2(KEYINPUT26), .ZN(new_n681));
  AND4_X1   g0481(.A1(new_n516), .A2(new_n523), .A3(new_n612), .A4(new_n528), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n576), .A2(new_n676), .A3(new_n607), .A4(new_n603), .ZN(new_n683));
  OAI211_X1 g0483(.A(new_n678), .B(new_n681), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n660), .B1(new_n460), .B2(new_n685), .ZN(G369));
  NAND2_X1  g0486(.A1(new_n499), .A2(new_n220), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n687), .A2(KEYINPUT27), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(KEYINPUT27), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(G213), .A3(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G343), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n518), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n528), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n693), .B1(new_n524), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n531), .B2(new_n693), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n587), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n406), .B1(new_n699), .B2(new_n585), .ZN(new_n700));
  INV_X1    g0500(.A(new_n600), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n601), .A2(new_n425), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(G179), .B2(new_n601), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n692), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT94), .ZN(new_n707));
  INV_X1    g0507(.A(new_n692), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n611), .A2(new_n708), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n709), .A2(new_n603), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n706), .B(new_n707), .C1(new_n710), .C2(new_n705), .ZN(new_n711));
  AOI22_X1  g0511(.A1(new_n709), .A2(new_n603), .B1(new_n610), .B2(new_n611), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n612), .A2(new_n708), .ZN(new_n713));
  OAI21_X1  g0513(.A(KEYINPUT94), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n698), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n694), .B1(new_n524), .B2(KEYINPUT91), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n708), .B1(new_n717), .B2(new_n527), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n715), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n716), .A2(new_n706), .A3(new_n719), .ZN(G399));
  INV_X1    g0520(.A(new_n216), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(G41), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n224), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n489), .A2(G116), .A3(new_n634), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G1), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n723), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT28), .ZN(new_n727));
  INV_X1    g0527(.A(G330), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT95), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(KEYINPUT30), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n620), .A2(new_n627), .A3(new_n594), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(new_n521), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n730), .B1(new_n732), .B2(new_n604), .ZN(new_n733));
  INV_X1    g0533(.A(new_n730), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n574), .A2(new_n521), .A3(new_n731), .A4(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n673), .A2(G179), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n604), .A2(new_n480), .A3(new_n601), .A4(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n733), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(KEYINPUT31), .B1(new_n738), .B2(new_n708), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n738), .A2(KEYINPUT31), .A3(new_n708), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n739), .B1(KEYINPUT96), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n738), .A2(new_n708), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT31), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n742), .A2(KEYINPUT96), .A3(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n608), .A2(new_n652), .A3(new_n708), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n747), .A2(new_n527), .A3(new_n717), .A4(new_n530), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n728), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n525), .A2(new_n527), .A3(new_n528), .A4(new_n612), .ZN(new_n750));
  INV_X1    g0550(.A(new_n683), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n675), .B1(new_n667), .B2(new_n668), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n670), .B1(new_n753), .B2(new_n677), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n672), .B1(new_n680), .B2(KEYINPUT26), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n708), .B1(new_n752), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(KEYINPUT29), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n684), .A2(new_n692), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT29), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n749), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n727), .B1(new_n762), .B2(G1), .ZN(G364));
  NOR2_X1   g0563(.A1(new_n498), .A2(G20), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n283), .B1(new_n764), .B2(G45), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n722), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n698), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(G330), .B2(new_n696), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n721), .A2(new_n301), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G355), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(G116), .B2(new_n216), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n358), .A2(new_n360), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n721), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(new_n248), .B2(new_n224), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n241), .A2(G45), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n772), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n220), .B1(KEYINPUT97), .B2(new_n425), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n425), .A2(KEYINPUT97), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n219), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G13), .A2(G33), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G20), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n767), .B1(new_n778), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n220), .A2(new_n295), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n290), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n789), .A2(new_n395), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n790), .A2(KEYINPUT98), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(KEYINPUT98), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n370), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n788), .A2(G200), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(G190), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n301), .B1(new_n797), .B2(G68), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n796), .A2(new_n395), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n220), .A2(G179), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n801), .A2(G190), .A3(G200), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n800), .A2(new_n202), .B1(new_n633), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n789), .A2(G190), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(G179), .A2(G200), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n220), .B1(new_n806), .B2(G190), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n805), .A2(new_n264), .B1(new_n807), .B2(new_n485), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n803), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n806), .A2(G20), .A3(new_n455), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n810), .A2(KEYINPUT32), .A3(new_n351), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT32), .ZN(new_n812));
  INV_X1    g0612(.A(new_n810), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n812), .B1(new_n813), .B2(G159), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n801), .A2(new_n455), .A3(G200), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n811), .B(new_n814), .C1(G107), .C2(new_n816), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n795), .A2(new_n798), .A3(new_n809), .A4(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(G322), .ZN(new_n819));
  INV_X1    g0619(.A(new_n797), .ZN(new_n820));
  XOR2_X1   g0620(.A(KEYINPUT33), .B(G317), .Z(new_n821));
  OAI22_X1  g0621(.A1(new_n793), .A2(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT99), .ZN(new_n823));
  INV_X1    g0623(.A(G311), .ZN(new_n824));
  INV_X1    g0624(.A(G294), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n805), .A2(new_n824), .B1(new_n807), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(G283), .ZN(new_n827));
  INV_X1    g0627(.A(G303), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n815), .A2(new_n827), .B1(new_n802), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n799), .A2(G326), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n259), .B1(new_n813), .B2(G329), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n818), .B1(new_n823), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n787), .B1(new_n834), .B2(new_n781), .ZN(new_n835));
  INV_X1    g0635(.A(new_n784), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n835), .B1(new_n696), .B2(new_n836), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n769), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(G396));
  AOI21_X1  g0639(.A(new_n457), .B1(new_n444), .B2(new_n708), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(new_n454), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n454), .A2(new_n692), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n684), .A2(new_n692), .A3(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n840), .A2(new_n454), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n842), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT103), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n849), .A2(new_n759), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT104), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n846), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n851), .B2(new_n850), .ZN(new_n853));
  INV_X1    g0653(.A(new_n749), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n767), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n854), .B2(new_n853), .ZN(new_n856));
  INV_X1    g0656(.A(new_n802), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n857), .A2(G107), .B1(new_n816), .B2(G87), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n828), .B2(new_n800), .ZN(new_n859));
  OAI22_X1  g0659(.A1(new_n805), .A2(new_n491), .B1(new_n820), .B2(new_n827), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n301), .B1(new_n810), .B2(new_n824), .C1(new_n485), .C2(new_n807), .ZN(new_n861));
  NOR3_X1   g0661(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n825), .B2(new_n793), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT101), .ZN(new_n864));
  AOI22_X1  g0664(.A1(G137), .A2(new_n799), .B1(new_n804), .B2(G159), .ZN(new_n865));
  INV_X1    g0665(.A(G150), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n865), .B1(new_n866), .B2(new_n820), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n794), .B2(G143), .ZN(new_n868));
  XOR2_X1   g0668(.A(new_n868), .B(KEYINPUT34), .Z(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n870), .A2(KEYINPUT102), .ZN(new_n871));
  INV_X1    g0671(.A(new_n773), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n857), .A2(G50), .B1(new_n816), .B2(G68), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n276), .B2(new_n807), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n872), .B(new_n874), .C1(G132), .C2(new_n813), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n870), .B2(KEYINPUT102), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n864), .B1(new_n871), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n781), .ZN(new_n878));
  INV_X1    g0678(.A(new_n767), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n781), .A2(new_n782), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n880), .B(KEYINPUT100), .Z(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n879), .B1(new_n882), .B2(new_n264), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n878), .B(new_n883), .C1(new_n844), .C2(new_n783), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n856), .A2(new_n884), .ZN(G384));
  OR2_X1    g0685(.A1(new_n540), .A2(KEYINPUT35), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n540), .A2(KEYINPUT35), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n886), .A2(G116), .A3(new_n221), .A4(new_n887), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n888), .B(KEYINPUT36), .Z(new_n889));
  OAI211_X1 g0689(.A(new_n224), .B(G77), .C1(new_n353), .C2(new_n276), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n202), .A2(G68), .ZN(new_n891));
  AOI211_X1 g0691(.A(new_n283), .B(G13), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n742), .A2(new_n743), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n894), .A2(new_n740), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n576), .A2(new_n607), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n612), .A2(new_n643), .A3(new_n651), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n896), .A2(new_n897), .A3(new_n603), .A4(new_n692), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n895), .B1(new_n531), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n344), .A2(new_n692), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n346), .A2(new_n349), .A3(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n349), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n900), .B1(new_n657), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n848), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n899), .A2(new_n905), .A3(KEYINPUT40), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT105), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n423), .A2(new_n907), .A3(new_n691), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT105), .B1(new_n411), .B2(new_n690), .ZN(new_n909));
  INV_X1    g0709(.A(new_n656), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n908), .B(new_n909), .C1(new_n910), .C2(new_n417), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT106), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n400), .A2(new_n401), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n913), .B1(new_n914), .B2(new_n423), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n411), .A2(new_n415), .A3(KEYINPUT106), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT107), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n915), .A2(new_n916), .A3(new_n917), .A4(new_n430), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n909), .A2(new_n908), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n402), .A2(new_n913), .B1(new_n423), .B2(new_n426), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n917), .B1(new_n921), .B2(new_n916), .ZN(new_n922));
  OAI21_X1  g0722(.A(KEYINPUT37), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT37), .B1(new_n411), .B2(new_n415), .ZN(new_n924));
  INV_X1    g0724(.A(new_n908), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n907), .B1(new_n423), .B2(new_n691), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n430), .B(new_n924), .C1(new_n925), .C2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT108), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n912), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n927), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n915), .A2(new_n430), .A3(new_n916), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT107), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n933), .A2(new_n919), .A3(new_n918), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n931), .B1(new_n934), .B2(KEYINPUT37), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT108), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT38), .B1(new_n930), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n421), .A2(G68), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT16), .B1(new_n938), .B2(new_n355), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n364), .A2(new_n281), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n379), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n691), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n426), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n942), .A2(new_n943), .A3(new_n402), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(KEYINPUT37), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n927), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n946), .B(KEYINPUT38), .C1(new_n435), .C2(new_n942), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n906), .B1(new_n937), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n946), .B1(new_n435), .B2(new_n942), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT38), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n947), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n953), .A2(new_n899), .A3(new_n905), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT40), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n949), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n459), .A2(new_n899), .ZN(new_n958));
  OAI21_X1  g0758(.A(G330), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(new_n957), .B2(new_n958), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n902), .A2(new_n904), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(new_n842), .B2(new_n845), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n963), .A2(new_n953), .B1(new_n910), .B2(new_n690), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n911), .B1(new_n935), .B2(KEYINPUT108), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n928), .A2(new_n929), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n951), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n948), .A2(KEYINPUT39), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n967), .A2(new_n968), .B1(KEYINPUT39), .B2(new_n953), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n657), .A2(new_n692), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n964), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n758), .A2(new_n459), .A3(new_n761), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n972), .A2(new_n660), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n971), .B(new_n973), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n960), .A2(new_n974), .B1(new_n283), .B2(new_n764), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n960), .A2(new_n974), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n893), .B1(new_n975), .B2(new_n976), .ZN(G367));
  NOR2_X1   g0777(.A1(new_n642), .A2(new_n692), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n679), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n675), .B2(new_n978), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n550), .A2(new_n708), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n896), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n575), .A2(new_n550), .A3(new_n708), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n718), .A2(new_n715), .A3(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT42), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n985), .A2(new_n705), .B1(new_n575), .B2(new_n554), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n987), .A2(new_n988), .B1(new_n708), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(KEYINPUT109), .B1(new_n987), .B2(new_n988), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n987), .A2(KEYINPUT109), .A3(new_n988), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n990), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT110), .Z(new_n996));
  OAI21_X1  g0796(.A(new_n981), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n985), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n716), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n981), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n996), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n993), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1002), .A2(new_n991), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1000), .B(new_n1001), .C1(new_n1003), .C2(new_n990), .ZN(new_n1004));
  AND3_X1   g0804(.A1(new_n997), .A2(new_n999), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n999), .B1(new_n997), .B2(new_n1004), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n722), .B(KEYINPUT41), .Z(new_n1008));
  INV_X1    g0808(.A(new_n716), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n719), .A2(new_n706), .A3(new_n985), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(KEYINPUT111), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT111), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n719), .A2(new_n1012), .A3(new_n706), .A4(new_n985), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1011), .A2(KEYINPUT45), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n719), .A2(new_n706), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n998), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT44), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(KEYINPUT44), .B1(new_n1015), .B2(new_n998), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1014), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(KEYINPUT45), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1009), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n718), .B(new_n715), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n698), .B(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n762), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1016), .B(new_n1017), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1021), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1027), .A2(new_n1028), .A3(new_n716), .A4(new_n1014), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1022), .A2(new_n1026), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1008), .B1(new_n1030), .B2(new_n762), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1007), .B1(new_n1031), .B2(new_n766), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT112), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1007), .B(KEYINPUT112), .C1(new_n1031), .C2(new_n766), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n775), .A2(new_n233), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n785), .B1(new_n216), .B2(new_n441), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n767), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n807), .A2(new_n353), .ZN(new_n1040));
  INV_X1    g0840(.A(G137), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n259), .B1(new_n810), .B2(new_n1041), .C1(new_n805), .C2(new_n202), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1040), .B(new_n1042), .C1(G143), .C2(new_n799), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n802), .A2(new_n276), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n815), .A2(new_n264), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1044), .B(new_n1045), .C1(G159), .C2(new_n797), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1043), .B(new_n1046), .C1(new_n866), .C2(new_n793), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n827), .A2(new_n805), .B1(new_n800), .B2(new_n824), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n773), .B(new_n1048), .C1(G317), .C2(new_n813), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n857), .A2(G116), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT46), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n794), .A2(G303), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n820), .A2(new_n825), .B1(new_n537), .B2(new_n815), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n807), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1053), .B1(G107), .B2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1049), .A2(new_n1051), .A3(new_n1052), .A4(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1047), .A2(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT47), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1039), .B1(new_n1058), .B2(new_n781), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n980), .A2(new_n836), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1036), .A2(new_n1061), .ZN(G387));
  INV_X1    g0862(.A(KEYINPUT115), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1024), .A2(new_n762), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1025), .A2(new_n1064), .A3(new_n247), .A4(new_n216), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n715), .A2(new_n836), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n230), .A2(new_n248), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n724), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1067), .A2(new_n774), .B1(new_n1068), .B2(new_n770), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n439), .A2(new_n202), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT50), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n248), .B1(new_n353), .B2(new_n264), .ZN(new_n1072));
  NOR3_X1   g0872(.A1(new_n1071), .A2(new_n1068), .A3(new_n1072), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1069), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n538), .B2(new_n721), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n767), .B1(new_n1075), .B2(new_n786), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n353), .A2(new_n805), .B1(new_n820), .B2(new_n277), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT113), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n800), .A2(new_n351), .B1(new_n485), .B2(new_n815), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n773), .B1(new_n866), .B2(new_n810), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n802), .A2(new_n264), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n807), .A2(new_n441), .ZN(new_n1082));
  NOR4_X1   g0882(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1078), .B(new_n1083), .C1(new_n202), .C2(new_n793), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n794), .A2(G317), .B1(G303), .B2(new_n804), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n1085), .A2(KEYINPUT114), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(KEYINPUT114), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(G322), .A2(new_n799), .B1(new_n797), .B2(G311), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT48), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n802), .A2(new_n825), .B1(new_n807), .B2(new_n827), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1091), .A2(KEYINPUT49), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n773), .B1(G326), .B2(new_n813), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1094), .B(new_n1095), .C1(new_n491), .C2(new_n815), .ZN(new_n1096));
  AOI21_X1  g0896(.A(KEYINPUT49), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1084), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n1066), .B(new_n1076), .C1(new_n1098), .C2(new_n781), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(new_n1024), .B2(new_n766), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1063), .B1(new_n1065), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1065), .A2(new_n1063), .A3(new_n1100), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(G393));
  NAND3_X1  g0904(.A1(new_n1022), .A2(new_n1029), .A3(new_n766), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n238), .A2(new_n775), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n785), .B1(new_n216), .B2(new_n537), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n767), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n794), .A2(G311), .B1(G317), .B2(new_n799), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT52), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n301), .B1(new_n810), .B2(new_n819), .C1(new_n815), .C2(new_n538), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n805), .A2(new_n825), .B1(new_n820), .B2(new_n828), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n802), .A2(new_n827), .B1(new_n807), .B2(new_n491), .ZN(new_n1113));
  OR4_X1    g0913(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n872), .B1(G143), .B2(new_n813), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1115), .B1(new_n353), .B2(new_n802), .C1(new_n633), .C2(new_n815), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n807), .A2(new_n264), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n804), .B2(new_n439), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n202), .B2(new_n820), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n794), .A2(G159), .B1(G150), .B2(new_n799), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1120), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT117), .ZN(new_n1126));
  OR2_X1    g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1114), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1108), .B1(new_n1129), .B2(new_n781), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n985), .B2(new_n836), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1030), .A2(new_n722), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1026), .B1(new_n1022), .B2(new_n1029), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1105), .B(new_n1131), .C1(new_n1132), .C2(new_n1133), .ZN(G390));
  XOR2_X1   g0934(.A(new_n970), .B(KEYINPUT118), .Z(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(new_n967), .B2(new_n947), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n708), .B(new_n841), .C1(new_n752), .C2(new_n756), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n961), .B1(new_n1137), .B2(new_n843), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n845), .A2(new_n842), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n961), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n970), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n967), .A2(new_n968), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n953), .A2(KEYINPUT39), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n749), .A2(new_n844), .A3(new_n961), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n1139), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n728), .B1(new_n748), .B2(new_n895), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1148), .A2(new_n905), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n1139), .B2(new_n1145), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1147), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n969), .A2(new_n782), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n882), .A2(new_n277), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n827), .A2(new_n800), .B1(new_n805), .B2(new_n537), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(G107), .B2(new_n797), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n301), .B1(new_n810), .B2(new_n825), .C1(new_n802), .C2(new_n633), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1117), .B(new_n1157), .C1(G68), .C2(new_n816), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1156), .B(new_n1158), .C1(new_n491), .C2(new_n793), .ZN(new_n1159));
  INV_X1    g0959(.A(G128), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n1160), .A2(new_n800), .B1(new_n820), .B2(new_n1041), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(G159), .B2(new_n1054), .ZN(new_n1162));
  OAI21_X1  g0962(.A(KEYINPUT53), .B1(new_n802), .B2(new_n866), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n813), .A2(G125), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT54), .B(G143), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1163), .B(new_n1164), .C1(new_n805), .C2(new_n1165), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n802), .A2(KEYINPUT53), .A3(new_n866), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(G132), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1162), .B(new_n1168), .C1(new_n1169), .C2(new_n793), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n259), .B1(new_n815), .B2(new_n202), .ZN(new_n1171));
  XOR2_X1   g0971(.A(new_n1171), .B(KEYINPUT120), .Z(new_n1172));
  OAI21_X1  g0972(.A(new_n1159), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n879), .B(new_n1154), .C1(new_n1173), .C2(new_n781), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n1152), .A2(new_n766), .B1(new_n1153), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n459), .A2(new_n1148), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n972), .A2(new_n660), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n740), .A2(KEYINPUT96), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n894), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1179), .B(new_n744), .C1(new_n531), .C2(new_n898), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1180), .A2(G330), .A3(new_n844), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1181), .A2(new_n962), .B1(new_n905), .B2(new_n1148), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1140), .ZN(new_n1183));
  OAI21_X1  g0983(.A(KEYINPUT119), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT119), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n961), .B1(new_n749), .B2(new_n844), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1185), .B(new_n1140), .C1(new_n1186), .C2(new_n1149), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1184), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n899), .A2(G330), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n962), .B1(new_n1189), .B2(new_n849), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n843), .B1(new_n757), .B2(new_n847), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n1190), .A2(new_n1146), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1177), .B1(new_n1188), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n722), .B1(new_n1152), .B2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1139), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n969), .A2(new_n1142), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1196), .B1(new_n1197), .B2(new_n1150), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1192), .B1(new_n1184), .B2(new_n1187), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n1198), .A2(new_n1177), .A3(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1175), .B1(new_n1195), .B2(new_n1200), .ZN(G378));
  AOI21_X1  g1001(.A(new_n728), .B1(new_n954), .B2(new_n955), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n288), .A2(new_n690), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n298), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n298), .A2(new_n1205), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1204), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1208), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1210), .A2(new_n1206), .A3(new_n1203), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n949), .A2(new_n1202), .A3(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1212), .B1(new_n949), .B2(new_n1202), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n971), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1212), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n956), .A2(G330), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n899), .A2(new_n905), .A3(KEYINPUT40), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n967), .B2(new_n947), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1216), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n970), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n949), .A2(new_n1202), .A3(new_n1212), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1220), .A2(new_n1223), .A3(new_n964), .A4(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1215), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n766), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n767), .B1(new_n881), .B2(G50), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(G97), .A2(new_n797), .B1(new_n804), .B2(new_n639), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1229), .B1(new_n276), .B2(new_n815), .C1(new_n793), .C2(new_n538), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n872), .A2(new_n247), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n807), .A2(new_n353), .B1(new_n810), .B2(new_n827), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n800), .A2(new_n491), .B1(new_n264), .B2(new_n802), .ZN(new_n1233));
  NOR4_X1   g1033(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .A4(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(KEYINPUT58), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1231), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1236));
  XOR2_X1   g1036(.A(new_n1236), .B(KEYINPUT121), .Z(new_n1237));
  AND2_X1   g1037(.A1(new_n1235), .A2(new_n1237), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n799), .A2(G125), .B1(G150), .B2(new_n1054), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(G132), .B2(new_n797), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1165), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n804), .A2(G137), .B1(new_n857), .B2(new_n1242), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1241), .B(new_n1243), .C1(new_n1160), .C2(new_n793), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1244), .A2(KEYINPUT59), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(KEYINPUT59), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n816), .A2(G159), .ZN(new_n1247));
  AOI211_X1 g1047(.A(G33), .B(G41), .C1(new_n813), .C2(G124), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n1238), .B1(KEYINPUT58), .B2(new_n1234), .C1(new_n1245), .C2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1228), .B1(new_n1250), .B2(new_n781), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n1212), .B2(new_n783), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1227), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1177), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1226), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT57), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n722), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1257), .B1(new_n1215), .B2(new_n1225), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1259), .B1(new_n1255), .B2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1253), .B1(new_n1258), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(G375));
  NAND2_X1  g1063(.A1(new_n1188), .A2(new_n1193), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1264), .A2(new_n1254), .ZN(new_n1265));
  NOR3_X1   g1065(.A1(new_n1265), .A2(new_n1008), .A3(new_n1194), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n962), .A2(new_n782), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n767), .B1(new_n881), .B2(G68), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n805), .A2(new_n866), .B1(new_n815), .B2(new_n276), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n872), .B(new_n1269), .C1(G128), .C2(new_n813), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n794), .A2(G137), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n799), .A2(G132), .B1(G50), .B2(new_n1054), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n797), .A2(new_n1242), .B1(new_n857), .B2(G159), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .A4(new_n1273), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n259), .B(new_n1045), .C1(G303), .C2(new_n813), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n802), .A2(new_n485), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n1082), .B(new_n1276), .C1(G294), .C2(new_n799), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1275), .B(new_n1277), .C1(new_n793), .C2(new_n827), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(G107), .A2(new_n804), .B1(new_n797), .B2(G116), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1279), .B(KEYINPUT122), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1274), .B1(new_n1278), .B2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1268), .B1(new_n1281), .B2(new_n781), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n1264), .A2(new_n766), .B1(new_n1267), .B2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1266), .A2(new_n1284), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1285), .B(KEYINPUT123), .ZN(G381));
  XOR2_X1   g1086(.A(new_n1262), .B(KEYINPUT124), .Z(new_n1287));
  NAND3_X1  g1087(.A1(new_n1102), .A2(new_n838), .A3(new_n1103), .ZN(new_n1288));
  OR3_X1    g1088(.A1(new_n1288), .A2(G384), .A3(G378), .ZN(new_n1289));
  NOR3_X1   g1089(.A1(new_n1287), .A2(G381), .A3(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1061), .ZN(new_n1291));
  AOI211_X1 g1091(.A(new_n1291), .B(G390), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(G407));
  INV_X1    g1093(.A(G378), .ZN(new_n1294));
  INV_X1    g1094(.A(G213), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1295), .A2(G343), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1294), .A2(new_n1296), .ZN(new_n1297));
  OAI211_X1 g1097(.A(G407), .B(G213), .C1(new_n1287), .C2(new_n1297), .ZN(G409));
  INV_X1    g1098(.A(KEYINPUT127), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1103), .ZN(new_n1300));
  OAI21_X1  g1100(.A(G396), .B1(new_n1300), .B2(new_n1101), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1301), .A2(new_n1288), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1291), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1303));
  INV_X1    g1103(.A(G390), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  OAI211_X1 g1105(.A(new_n1299), .B(new_n1302), .C1(new_n1305), .C2(new_n1292), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1299), .B1(new_n1301), .B2(new_n1288), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1307), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(G387), .A2(G390), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1302), .A2(new_n1299), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1308), .A2(new_n1309), .A3(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1306), .A2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT61), .ZN(new_n1313));
  INV_X1    g1113(.A(G384), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1199), .A2(KEYINPUT60), .A3(new_n1177), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(new_n722), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1194), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(KEYINPUT60), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1265), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1316), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1314), .B1(new_n1320), .B2(new_n1284), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1265), .B1(KEYINPUT60), .B2(new_n1317), .ZN(new_n1322));
  OAI211_X1 g1122(.A(G384), .B(new_n1283), .C1(new_n1322), .C2(new_n1316), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1296), .A2(G2897), .ZN(new_n1324));
  AND3_X1   g1124(.A1(new_n1321), .A2(new_n1323), .A3(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1324), .B1(new_n1321), .B2(new_n1323), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT126), .ZN(new_n1328));
  NOR3_X1   g1128(.A1(new_n1213), .A2(new_n971), .A3(new_n1214), .ZN(new_n1329));
  AOI22_X1  g1129(.A1(new_n1220), .A2(new_n1224), .B1(new_n1223), .B2(new_n964), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1328), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1215), .A2(new_n1225), .A3(KEYINPUT126), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1331), .A2(new_n766), .A3(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1008), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1255), .A2(new_n1334), .A3(new_n1226), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1333), .A2(new_n1335), .A3(new_n1252), .ZN(new_n1336));
  AND2_X1   g1136(.A1(new_n1294), .A2(new_n1336), .ZN(new_n1337));
  AND2_X1   g1137(.A1(new_n1227), .A2(new_n1252), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1177), .B1(new_n1152), .B2(new_n1194), .ZN(new_n1339));
  OAI21_X1  g1139(.A(KEYINPUT57), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n722), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1341));
  AOI21_X1  g1141(.A(KEYINPUT57), .B1(new_n1255), .B2(new_n1226), .ZN(new_n1342));
  OAI211_X1 g1142(.A(G378), .B(new_n1338), .C1(new_n1341), .C2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT125), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1258), .A2(new_n1261), .ZN(new_n1346));
  NAND4_X1  g1146(.A1(new_n1346), .A2(KEYINPUT125), .A3(G378), .A4(new_n1338), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1337), .B1(new_n1345), .B2(new_n1347), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1327), .B1(new_n1348), .B2(new_n1296), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1321), .A2(new_n1323), .ZN(new_n1350));
  NOR3_X1   g1150(.A1(new_n1348), .A2(new_n1296), .A3(new_n1350), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT62), .ZN(new_n1352));
  OAI211_X1 g1152(.A(new_n1313), .B(new_n1349), .C1(new_n1351), .C2(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(new_n1296), .ZN(new_n1354));
  INV_X1    g1154(.A(new_n1350), .ZN(new_n1355));
  AOI21_X1  g1155(.A(KEYINPUT125), .B1(new_n1262), .B2(G378), .ZN(new_n1356));
  NOR2_X1   g1156(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1357));
  NOR2_X1   g1157(.A1(new_n1356), .A2(new_n1357), .ZN(new_n1358));
  OAI211_X1 g1158(.A(new_n1354), .B(new_n1355), .C1(new_n1358), .C2(new_n1337), .ZN(new_n1359));
  NOR2_X1   g1159(.A1(new_n1359), .A2(KEYINPUT62), .ZN(new_n1360));
  OAI21_X1  g1160(.A(new_n1312), .B1(new_n1353), .B2(new_n1360), .ZN(new_n1361));
  AND2_X1   g1161(.A1(new_n1349), .A2(new_n1313), .ZN(new_n1362));
  AND2_X1   g1162(.A1(new_n1306), .A2(new_n1311), .ZN(new_n1363));
  INV_X1    g1163(.A(KEYINPUT63), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1359), .A2(new_n1364), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1351), .A2(KEYINPUT63), .ZN(new_n1366));
  NAND4_X1  g1166(.A1(new_n1362), .A2(new_n1363), .A3(new_n1365), .A4(new_n1366), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1361), .A2(new_n1367), .ZN(G405));
  OAI22_X1  g1168(.A1(new_n1356), .A2(new_n1357), .B1(G378), .B2(new_n1262), .ZN(new_n1369));
  AND2_X1   g1169(.A1(new_n1369), .A2(new_n1355), .ZN(new_n1370));
  NOR2_X1   g1170(.A1(new_n1369), .A2(new_n1355), .ZN(new_n1371));
  OR3_X1    g1171(.A1(new_n1312), .A2(new_n1370), .A3(new_n1371), .ZN(new_n1372));
  OAI21_X1  g1172(.A(new_n1312), .B1(new_n1370), .B2(new_n1371), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1372), .A2(new_n1373), .ZN(G402));
endmodule


