//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 0 1 1 0 1 0 0 0 0 0 0 0 1 1 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n541,
    new_n542, new_n543, new_n544, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n554, new_n555, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n571, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT65), .Z(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n451), .A2(new_n456), .B1(new_n457), .B2(new_n452), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT66), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND3_X1   g036(.A1(new_n460), .A2(new_n461), .A3(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n460), .B1(G2104), .B2(new_n461), .ZN(new_n463));
  OAI21_X1  g038(.A(G101), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OR2_X1    g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(G137), .A3(new_n461), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(G125), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n461), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n469), .A2(new_n474), .ZN(G160));
  OAI21_X1  g050(.A(new_n461), .B1(new_n470), .B2(new_n471), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  INV_X1    g053(.A(G124), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n467), .A2(G2105), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n461), .A2(G112), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  OAI221_X1 g057(.A(new_n478), .B1(new_n479), .B2(new_n480), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  XOR2_X1   g058(.A(new_n483), .B(KEYINPUT68), .Z(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  INV_X1    g060(.A(KEYINPUT71), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(KEYINPUT70), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g064(.A(G138), .B1(new_n486), .B2(new_n487), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n489), .B1(new_n476), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n492), .B1(KEYINPUT71), .B2(KEYINPUT4), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n467), .A2(new_n493), .A3(new_n461), .A4(new_n488), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n496));
  OAI211_X1 g071(.A(G126), .B(G2105), .C1(new_n470), .C2(new_n471), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n498), .A2(new_n500), .A3(G2104), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n496), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n497), .A2(new_n496), .A3(new_n501), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n495), .B1(new_n503), .B2(new_n504), .ZN(G164));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT72), .A2(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT72), .A2(G543), .ZN(new_n509));
  OAI211_X1 g084(.A(new_n507), .B(KEYINPUT5), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT72), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT72), .A2(G543), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT73), .B1(new_n515), .B2(KEYINPUT5), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n510), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G62), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n506), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n517), .A2(G88), .A3(new_n523), .ZN(new_n524));
  OAI21_X1  g099(.A(G543), .B1(new_n521), .B2(new_n522), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G50), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n520), .A2(new_n528), .ZN(G166));
  NAND3_X1  g104(.A1(new_n517), .A2(G89), .A3(new_n523), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n525), .A2(KEYINPUT74), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT74), .ZN(new_n533));
  OAI211_X1 g108(.A(new_n533), .B(G543), .C1(new_n521), .C2(new_n522), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G51), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n530), .A2(new_n531), .A3(new_n536), .A4(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  AND2_X1   g115(.A1(new_n517), .A2(new_n523), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G90), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n535), .A2(G52), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  OAI211_X1 g119(.A(new_n542), .B(new_n543), .C1(new_n506), .C2(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  AOI22_X1  g121(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n506), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n541), .A2(G81), .B1(G43), .B2(new_n535), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  INV_X1    g131(.A(G53), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT9), .B1(new_n525), .B2(new_n557), .ZN(new_n558));
  OR3_X1    g133(.A1(new_n525), .A2(KEYINPUT9), .A3(new_n557), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n541), .A2(G91), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT76), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n517), .A2(KEYINPUT75), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT75), .ZN(new_n563));
  OAI211_X1 g138(.A(new_n510), .B(new_n563), .C1(new_n514), .C2(new_n516), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(G65), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n561), .B1(new_n567), .B2(G651), .ZN(new_n568));
  AOI211_X1 g143(.A(KEYINPUT76), .B(new_n506), .C1(new_n565), .C2(new_n566), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n560), .B1(new_n568), .B2(new_n569), .ZN(G299));
  AOI22_X1  g145(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n571));
  OAI211_X1 g146(.A(new_n524), .B(new_n527), .C1(new_n571), .C2(new_n506), .ZN(G303));
  NAND2_X1  g147(.A1(new_n541), .A2(G87), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n526), .A2(G49), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G288));
  INV_X1    g151(.A(KEYINPUT77), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n517), .A2(G61), .ZN(new_n578));
  AND2_X1   g153(.A1(G73), .A2(G543), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n577), .B(G651), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n579), .B1(new_n517), .B2(G61), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT77), .B1(new_n581), .B2(new_n506), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n526), .A2(G48), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n517), .A2(new_n523), .ZN(new_n585));
  INV_X1    g160(.A(G86), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n583), .A2(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n590), .A2(new_n506), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n541), .A2(G85), .B1(G47), .B2(new_n535), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(G290));
  INV_X1    g168(.A(KEYINPUT78), .ZN(new_n594));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(G171), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(G301), .A2(KEYINPUT78), .A3(G868), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n585), .B2(new_n599), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n517), .A2(KEYINPUT10), .A3(G92), .A4(new_n523), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n535), .A2(G54), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AND2_X1   g179(.A1(new_n562), .A2(new_n564), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G66), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n604), .B1(G651), .B2(new_n608), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n596), .B(new_n597), .C1(new_n609), .C2(G868), .ZN(G284));
  XNOR2_X1  g185(.A(G284), .B(KEYINPUT79), .ZN(G321));
  NAND2_X1  g186(.A1(G299), .A2(new_n595), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(new_n595), .B2(G168), .ZN(G297));
  XOR2_X1   g188(.A(G297), .B(KEYINPUT80), .Z(G280));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n609), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND2_X1  g191(.A1(new_n550), .A2(new_n595), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n600), .A2(new_n601), .B1(G54), .B2(new_n535), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n605), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n506), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n620), .A2(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n617), .B1(new_n621), .B2(new_n595), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g198(.A1(new_n462), .A2(new_n463), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(new_n467), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT81), .B(G2100), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT82), .Z(new_n630));
  NAND2_X1  g205(.A1(new_n477), .A2(G135), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT83), .ZN(new_n632));
  OAI21_X1  g207(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n633));
  INV_X1    g208(.A(G111), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n633), .B1(new_n634), .B2(G2105), .ZN(new_n635));
  INV_X1    g210(.A(new_n480), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(G123), .ZN(new_n637));
  AND2_X1   g212(.A1(new_n632), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2096), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n630), .B(new_n639), .C1(new_n628), .C2(new_n627), .ZN(G156));
  XOR2_X1   g215(.A(G2451), .B(G2454), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(KEYINPUT14), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2427), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2430), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n649), .B1(new_n648), .B2(new_n647), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n644), .B(new_n650), .Z(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  AND3_X1   g229(.A1(new_n653), .A2(G14), .A3(new_n654), .ZN(G401));
  XNOR2_X1  g230(.A(G2072), .B(G2078), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT84), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT17), .ZN(new_n659));
  XOR2_X1   g234(.A(G2067), .B(G2678), .Z(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2084), .B(G2090), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n659), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n662), .B1(new_n658), .B2(new_n661), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n659), .B2(new_n661), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n660), .A2(new_n662), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n658), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT18), .ZN(new_n668));
  OR3_X1    g243(.A1(new_n663), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n669), .A2(KEYINPUT85), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(KEYINPUT85), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2096), .B(G2100), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n670), .A2(new_n671), .A3(new_n673), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(G227));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT86), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1956), .B(G2474), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n680), .A2(new_n682), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT20), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n680), .B1(new_n682), .B2(new_n684), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n682), .A2(new_n684), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OAI211_X1 g264(.A(new_n686), .B(new_n689), .C1(new_n679), .C2(new_n688), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1991), .B(G1996), .Z(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n692), .A2(new_n694), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n695), .A2(new_n698), .A3(new_n696), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(G229));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G23), .ZN(new_n705));
  INV_X1    g280(.A(G288), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(new_n704), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT33), .B(G1976), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT87), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n707), .B(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n704), .A2(G6), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n587), .B1(new_n580), .B2(new_n582), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(new_n704), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT32), .B(G1981), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n704), .A2(G22), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G166), .B2(new_n704), .ZN(new_n718));
  INV_X1    g293(.A(G1971), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n710), .A2(new_n715), .A3(new_n716), .A4(new_n720), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n721), .A2(KEYINPUT34), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(KEYINPUT34), .ZN(new_n723));
  MUX2_X1   g298(.A(G24), .B(G290), .S(G16), .Z(new_n724));
  AND2_X1   g299(.A1(new_n724), .A2(G1986), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(G1986), .ZN(new_n726));
  INV_X1    g301(.A(G29), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G25), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n636), .A2(G119), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n477), .A2(G131), .ZN(new_n730));
  OR2_X1    g305(.A1(G95), .A2(G2105), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n731), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n728), .B1(new_n734), .B2(new_n727), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT35), .B(G1991), .Z(new_n736));
  XOR2_X1   g311(.A(new_n735), .B(new_n736), .Z(new_n737));
  NOR3_X1   g312(.A1(new_n725), .A2(new_n726), .A3(new_n737), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n722), .A2(new_n723), .A3(new_n738), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT36), .Z(new_n740));
  NAND2_X1  g315(.A1(new_n704), .A2(G20), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT23), .Z(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G299), .B2(G16), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(G1956), .Z(new_n744));
  NOR2_X1   g319(.A1(G171), .A2(new_n704), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G5), .B2(new_n704), .ZN(new_n746));
  INV_X1    g321(.A(G1961), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT96), .Z(new_n749));
  NAND2_X1  g324(.A1(new_n727), .A2(G27), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT98), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G164), .B2(new_n727), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT99), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G2078), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n727), .A2(G35), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G162), .B2(new_n727), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT100), .B(KEYINPUT29), .ZN(new_n757));
  INV_X1    g332(.A(G2090), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n756), .B(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n747), .B2(new_n746), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n704), .A2(G21), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G168), .B2(new_n704), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT94), .B(G1966), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n749), .A2(new_n754), .A3(new_n761), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n727), .A2(G26), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT28), .Z(new_n768));
  AOI22_X1  g343(.A1(new_n636), .A2(G128), .B1(G140), .B2(new_n477), .ZN(new_n769));
  OAI21_X1  g344(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n770));
  INV_X1    g345(.A(G116), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(G2105), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT90), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n768), .B1(new_n774), .B2(G29), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G2067), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT27), .B(G1996), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n636), .A2(G129), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n624), .A2(G105), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n477), .A2(G141), .ZN(new_n780));
  NAND3_X1  g355(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT26), .Z(new_n782));
  NAND4_X1  g357(.A1(new_n778), .A2(new_n779), .A3(new_n780), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(G29), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n727), .A2(G32), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n777), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT31), .B(G11), .Z(new_n787));
  XOR2_X1   g362(.A(KEYINPUT95), .B(G28), .Z(new_n788));
  OR2_X1    g363(.A1(new_n788), .A2(KEYINPUT30), .ZN(new_n789));
  AOI21_X1  g364(.A(G29), .B1(new_n788), .B2(KEYINPUT30), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n787), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(new_n638), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT25), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n467), .A2(G127), .ZN(new_n795));
  NAND2_X1  g370(.A1(G115), .A2(G2104), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n461), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AOI211_X1 g372(.A(new_n794), .B(new_n797), .C1(G139), .C2(new_n477), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(G29), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G29), .B2(G33), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT91), .B(G2072), .Z(new_n801));
  OAI221_X1 g376(.A(new_n791), .B1(new_n727), .B2(new_n792), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  AOI211_X1 g377(.A(new_n786), .B(new_n802), .C1(new_n800), .C2(new_n801), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT24), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n804), .A2(G34), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(G34), .ZN(new_n806));
  AOI21_X1  g381(.A(G29), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(G160), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(G29), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT92), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(G2084), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n784), .A2(new_n785), .A3(new_n777), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT93), .ZN(new_n813));
  AND4_X1   g388(.A1(new_n776), .A2(new_n803), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(G4), .A2(G16), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT88), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n620), .B2(new_n704), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G1348), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n810), .A2(G2084), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT97), .ZN(new_n820));
  NOR2_X1   g395(.A1(G16), .A2(G19), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n551), .B2(G16), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT89), .B(G1341), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n814), .A2(new_n818), .A3(new_n820), .A4(new_n824), .ZN(new_n825));
  NOR4_X1   g400(.A1(new_n740), .A2(new_n744), .A3(new_n766), .A4(new_n825), .ZN(G311));
  OR4_X1    g401(.A1(new_n740), .A2(new_n744), .A3(new_n766), .A4(new_n825), .ZN(G150));
  NAND3_X1  g402(.A1(new_n517), .A2(G93), .A3(new_n523), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n535), .A2(G55), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(KEYINPUT101), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT101), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n828), .A2(new_n829), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n517), .A2(G67), .ZN(new_n835));
  INV_X1    g410(.A(G80), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n835), .B1(new_n836), .B2(new_n515), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(G651), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(G860), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT37), .Z(new_n841));
  INV_X1    g416(.A(KEYINPUT102), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n551), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  AOI22_X1  g418(.A1(new_n831), .A2(new_n833), .B1(G651), .B2(new_n837), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n844), .A2(KEYINPUT102), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n550), .B1(new_n844), .B2(KEYINPUT102), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n839), .A2(new_n842), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT38), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n620), .A2(new_n615), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n851), .A2(new_n853), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT39), .ZN(new_n857));
  AOI21_X1  g432(.A(G860), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n854), .A2(new_n855), .A3(KEYINPUT39), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n858), .A2(KEYINPUT103), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(KEYINPUT103), .B1(new_n858), .B2(new_n859), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n841), .B1(new_n860), .B2(new_n861), .ZN(G145));
  NAND2_X1  g437(.A1(new_n477), .A2(G142), .ZN(new_n863));
  INV_X1    g438(.A(G130), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n461), .A2(G118), .ZN(new_n865));
  OAI21_X1  g440(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n866));
  OAI221_X1 g441(.A(new_n863), .B1(new_n864), .B2(new_n480), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n626), .B(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n733), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n869), .A2(KEYINPUT104), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(KEYINPUT104), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n798), .B(new_n774), .Z(new_n873));
  NAND4_X1  g448(.A1(new_n491), .A2(new_n494), .A3(new_n497), .A4(new_n501), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n783), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n873), .A2(new_n875), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n877), .B1(new_n876), .B2(new_n878), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n871), .B(new_n872), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n484), .B(new_n808), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n792), .ZN(new_n884));
  INV_X1    g459(.A(new_n881), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n885), .A2(new_n879), .A3(new_n870), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n882), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(G37), .ZN(new_n888));
  INV_X1    g463(.A(new_n869), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n889), .A2(KEYINPUT105), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n890), .B1(new_n885), .B2(new_n879), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n885), .A2(new_n879), .A3(new_n890), .ZN(new_n892));
  INV_X1    g467(.A(new_n884), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n887), .B(new_n888), .C1(new_n891), .C2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT40), .ZN(G395));
  OR2_X1    g471(.A1(new_n568), .A2(new_n569), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n897), .A2(new_n560), .A3(new_n620), .ZN(new_n898));
  NAND2_X1  g473(.A1(G299), .A2(new_n609), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n897), .A2(KEYINPUT106), .A3(new_n560), .A4(new_n620), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n902), .B1(G299), .B2(new_n609), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n901), .A2(new_n903), .A3(new_n899), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT41), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n905), .B1(G299), .B2(new_n609), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n898), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n850), .B(new_n621), .ZN(new_n910));
  MUX2_X1   g485(.A(new_n900), .B(new_n909), .S(new_n910), .Z(new_n911));
  INV_X1    g486(.A(KEYINPUT108), .ZN(new_n912));
  XNOR2_X1  g487(.A(G290), .B(G303), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT107), .ZN(new_n914));
  NAND2_X1  g489(.A1(G288), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n573), .A2(KEYINPUT107), .A3(new_n574), .A4(new_n575), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n712), .ZN(new_n918));
  NAND3_X1  g493(.A1(G305), .A2(new_n915), .A3(new_n916), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n913), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n913), .B1(new_n919), .B2(new_n918), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n912), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n918), .A2(new_n919), .ZN(new_n924));
  INV_X1    g499(.A(new_n913), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n926), .A2(KEYINPUT108), .A3(new_n920), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT109), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(new_n929), .A3(KEYINPUT42), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n928), .A2(KEYINPUT42), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n921), .A2(new_n922), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT109), .B1(new_n932), .B2(KEYINPUT42), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n930), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n911), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n911), .A2(new_n934), .ZN(new_n936));
  OAI21_X1  g511(.A(G868), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n839), .A2(new_n595), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(G295));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n938), .ZN(G331));
  INV_X1    g515(.A(new_n928), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n542), .A2(new_n543), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n544), .A2(new_n506), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n943), .A2(KEYINPUT111), .A3(G286), .A4(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT111), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(G301), .B2(G168), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT110), .B1(G301), .B2(G168), .ZN(new_n950));
  NAND3_X1  g525(.A1(G301), .A2(KEYINPUT110), .A3(G168), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n949), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n843), .A2(new_n845), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n847), .A2(new_n848), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n950), .ZN(new_n957));
  AOI22_X1  g532(.A1(new_n957), .A2(new_n951), .B1(new_n948), .B2(new_n946), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n958), .A2(new_n846), .A3(new_n849), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT112), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n900), .A2(new_n905), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n901), .A2(new_n903), .A3(new_n907), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n961), .A2(new_n962), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n960), .A2(new_n900), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT112), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n960), .B1(new_n963), .B2(new_n964), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n941), .B(new_n966), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  AOI22_X1  g545(.A1(new_n904), .A2(new_n905), .B1(new_n898), .B2(new_n907), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n967), .B(new_n928), .C1(new_n971), .C2(new_n960), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n970), .A2(KEYINPUT43), .A3(new_n888), .A4(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT43), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n888), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n909), .A2(new_n961), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n928), .B1(new_n976), .B2(new_n967), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n974), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n973), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT44), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n970), .A2(new_n974), .A3(new_n888), .A4(new_n972), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT43), .B1(new_n975), .B2(new_n977), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT44), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n980), .A2(new_n985), .ZN(G397));
  INV_X1    g561(.A(G1384), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n874), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G40), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n469), .A2(new_n989), .A3(new_n474), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT45), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n988), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G2067), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n774), .B(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n992), .B1(new_n994), .B2(new_n877), .ZN(new_n995));
  INV_X1    g570(.A(new_n992), .ZN(new_n996));
  INV_X1    g571(.A(G1996), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n996), .A2(KEYINPUT46), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT46), .B1(new_n996), .B2(new_n997), .ZN(new_n999));
  OR3_X1    g574(.A1(new_n995), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT47), .ZN(new_n1001));
  OR2_X1    g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(G290), .A2(G1986), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1004), .A2(new_n992), .ZN(new_n1005));
  OR2_X1    g580(.A1(new_n1005), .A2(KEYINPUT48), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n783), .B(new_n997), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n994), .A2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g583(.A(new_n733), .B(new_n736), .Z(new_n1009));
  OAI21_X1  g584(.A(new_n996), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1005), .A2(KEYINPUT48), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1006), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n734), .A2(new_n736), .ZN(new_n1014));
  OAI22_X1  g589(.A1(new_n1008), .A2(new_n1014), .B1(G2067), .B2(new_n774), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n996), .ZN(new_n1016));
  AND4_X1   g591(.A1(new_n1002), .A2(new_n1012), .A3(new_n1013), .A4(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G1981), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n583), .A2(new_n1018), .A3(new_n588), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n581), .A2(new_n506), .ZN(new_n1020));
  OAI21_X1  g595(.A(G1981), .B1(new_n1020), .B2(new_n587), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT49), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1019), .A2(KEYINPUT49), .A3(new_n1021), .ZN(new_n1025));
  INV_X1    g600(.A(new_n474), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1026), .A2(G40), .A3(new_n464), .A4(new_n468), .ZN(new_n1027));
  OAI21_X1  g602(.A(G8), .B1(new_n988), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1024), .A2(new_n1025), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G8), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT50), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n497), .A2(new_n496), .A3(new_n501), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n491), .B(new_n494), .C1(new_n1033), .C2(new_n502), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1032), .B1(new_n1034), .B2(new_n987), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n874), .A2(new_n1032), .A3(new_n987), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n990), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n758), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT45), .B1(new_n1034), .B2(new_n987), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n991), .A2(G1384), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n874), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n990), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n719), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1031), .B1(new_n1039), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT114), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(G166), .B2(new_n1031), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT114), .ZN(new_n1050));
  NAND4_X1  g625(.A1(G303), .A2(new_n1050), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1047), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1045), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n706), .A2(G1976), .ZN(new_n1054));
  INV_X1    g629(.A(G1976), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT52), .B1(G288), .B2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1054), .A2(new_n1056), .A3(new_n1029), .ZN(new_n1057));
  NOR2_X1   g632(.A1(G288), .A2(new_n1055), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT52), .B1(new_n1058), .B2(new_n1028), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1030), .A2(new_n1053), .A3(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n991), .B1(G164), .B2(G1384), .ZN(new_n1063));
  INV_X1    g638(.A(G2078), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1027), .B1(new_n874), .B2(new_n1041), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n747), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1041), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT116), .B1(G164), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1027), .B1(new_n988), .B2(new_n991), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1034), .A2(new_n1073), .A3(new_n1041), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1067), .A2(G2078), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1071), .A2(new_n1072), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1068), .A2(new_n1069), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(G171), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT123), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1077), .A2(KEYINPUT123), .A3(G171), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1047), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1027), .B1(new_n988), .B2(KEYINPUT50), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1034), .A2(new_n1032), .A3(new_n987), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1084), .A2(new_n758), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1044), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(G8), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1083), .A2(new_n1088), .A3(KEYINPUT115), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT115), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1031), .B1(new_n1044), .B2(new_n1086), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1090), .B1(new_n1052), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1089), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1062), .A2(new_n1082), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1071), .A2(new_n1074), .A3(new_n1072), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(new_n764), .ZN(new_n1097));
  INV_X1    g672(.A(G2084), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1038), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1100), .A2(G8), .A3(G286), .ZN(new_n1101));
  OAI21_X1  g676(.A(G8), .B1(KEYINPUT121), .B2(KEYINPUT51), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1096), .A2(new_n764), .B1(new_n1038), .B2(new_n1098), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1102), .B1(new_n1103), .B2(G168), .ZN(new_n1104));
  NAND2_X1  g679(.A1(KEYINPUT121), .A2(KEYINPUT51), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1101), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1105), .ZN(new_n1107));
  AOI211_X1 g682(.A(new_n1102), .B(new_n1107), .C1(new_n1103), .C2(G168), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1095), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1102), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1110), .B1(new_n1100), .B2(G286), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n1107), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1112), .A2(KEYINPUT122), .A3(new_n1113), .A4(new_n1101), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1109), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1094), .B1(new_n1115), .B2(KEYINPUT62), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1109), .A2(new_n1114), .A3(new_n1117), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1116), .A2(KEYINPUT125), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT125), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT119), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n1103), .A2(new_n1031), .A3(G286), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT118), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1083), .B1(new_n1045), .B2(new_n1123), .ZN(new_n1124));
  AOI211_X1 g699(.A(KEYINPUT118), .B(new_n1031), .C1(new_n1039), .C2(new_n1044), .ZN(new_n1125));
  OAI211_X1 g700(.A(KEYINPUT63), .B(new_n1122), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1028), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1060), .B1(new_n1127), .B2(new_n1025), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n1053), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1121), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1093), .A2(new_n1128), .A3(new_n1053), .A4(new_n1122), .ZN(new_n1131));
  XOR2_X1   g706(.A(KEYINPUT117), .B(KEYINPUT63), .Z(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  OR2_X1    g708(.A1(new_n1045), .A2(new_n1123), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1125), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1134), .A2(new_n1135), .A3(new_n1083), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1122), .A2(KEYINPUT63), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1062), .A2(new_n1136), .A3(KEYINPUT119), .A4(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1130), .A2(new_n1133), .A3(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1030), .A2(new_n1055), .A3(new_n706), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1028), .B1(new_n1140), .B2(new_n1019), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1053), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1141), .B1(new_n1142), .B2(new_n1128), .ZN(new_n1143));
  OR2_X1    g718(.A1(KEYINPUT124), .A2(G2078), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1067), .B1(KEYINPUT124), .B2(G2078), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1072), .A2(new_n1042), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n1040), .A2(new_n1043), .A3(G2078), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1069), .B(new_n1146), .C1(new_n1147), .C2(KEYINPUT53), .ZN(new_n1148));
  OR2_X1    g723(.A1(new_n1148), .A2(G171), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1080), .A2(new_n1081), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT54), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1148), .A2(G171), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1068), .A2(G301), .A3(new_n1069), .A4(new_n1076), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1153), .A2(new_n1154), .A3(KEYINPUT54), .ZN(new_n1155));
  AND4_X1   g730(.A1(new_n1053), .A2(new_n1093), .A3(new_n1128), .A4(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1031), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n1111), .A2(new_n1107), .B1(G286), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(KEYINPUT122), .B1(new_n1158), .B2(new_n1113), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1106), .A2(new_n1095), .A3(new_n1108), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1152), .B(new_n1156), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(G1956), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1163));
  XNOR2_X1  g738(.A(KEYINPUT56), .B(G2072), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1162), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT57), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n1167), .B(new_n560), .C1(new_n568), .C2(new_n569), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1165), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n988), .A2(new_n1027), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n993), .ZN(new_n1171));
  INV_X1    g746(.A(G1348), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1172), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n620), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1174), .A2(new_n1166), .A3(new_n1168), .A4(new_n1165), .ZN(new_n1175));
  AND2_X1   g750(.A1(new_n1173), .A2(new_n1171), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(new_n620), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1166), .A2(new_n1168), .A3(new_n1165), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(new_n1174), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT60), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1176), .A2(new_n1181), .A3(new_n609), .ZN(new_n1182));
  NOR3_X1   g757(.A1(new_n1040), .A2(new_n1043), .A3(G1996), .ZN(new_n1183));
  XNOR2_X1  g758(.A(KEYINPUT58), .B(G1341), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1170), .A2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n551), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT59), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  OAI211_X1 g763(.A(KEYINPUT59), .B(new_n551), .C1(new_n1183), .C2(new_n1185), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1182), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  AOI22_X1  g765(.A1(new_n1178), .A2(KEYINPUT60), .B1(new_n1180), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1179), .A2(KEYINPUT120), .A3(new_n1192), .ZN(new_n1193));
  OAI211_X1 g768(.A(new_n1193), .B(new_n1180), .C1(new_n1192), .C2(new_n1179), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1169), .B1(new_n1191), .B2(new_n1194), .ZN(new_n1195));
  OAI211_X1 g770(.A(new_n1139), .B(new_n1143), .C1(new_n1161), .C2(new_n1195), .ZN(new_n1196));
  NOR3_X1   g771(.A1(new_n1119), .A2(new_n1120), .A3(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT113), .ZN(new_n1198));
  NAND2_X1  g773(.A1(G290), .A2(G1986), .ZN(new_n1199));
  AND3_X1   g774(.A1(new_n1004), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n996), .B1(new_n1199), .B2(new_n1198), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1010), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1017), .B1(new_n1197), .B2(new_n1202), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g778(.A1(new_n675), .A2(G319), .A3(new_n676), .ZN(new_n1205));
  INV_X1    g779(.A(KEYINPUT126), .ZN(new_n1206));
  XNOR2_X1  g780(.A(new_n1205), .B(new_n1206), .ZN(new_n1207));
  INV_X1    g781(.A(G401), .ZN(new_n1208));
  NAND2_X1  g782(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g783(.A1(new_n1209), .A2(KEYINPUT127), .ZN(new_n1210));
  AND2_X1   g784(.A1(new_n895), .A2(new_n702), .ZN(new_n1211));
  INV_X1    g785(.A(KEYINPUT127), .ZN(new_n1212));
  NAND3_X1  g786(.A1(new_n1207), .A2(new_n1212), .A3(new_n1208), .ZN(new_n1213));
  AND4_X1   g787(.A1(new_n983), .A2(new_n1210), .A3(new_n1211), .A4(new_n1213), .ZN(G308));
  NAND4_X1  g788(.A1(new_n983), .A2(new_n1210), .A3(new_n1211), .A4(new_n1213), .ZN(G225));
endmodule


