//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 0 1 0 0 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 0 1 1 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1250, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1298, new_n1299,
    new_n1300;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  INV_X1    g0002(.A(G58), .ZN(new_n203));
  INV_X1    g0003(.A(G68), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NOR3_X1   g0005(.A1(new_n202), .A2(G77), .A3(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT0), .Z(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n205), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n211), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT65), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n208), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  OR2_X1    g0025(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n217), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT66), .Z(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G226), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XOR2_X1   g0038(.A(G50), .B(G58), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G97), .B(G107), .Z(new_n241));
  XNOR2_X1  g0041(.A(G87), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  INV_X1    g0044(.A(KEYINPUT72), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT10), .ZN(new_n246));
  NOR2_X1   g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NOR2_X1   g0047(.A1(KEYINPUT72), .A2(KEYINPUT10), .ZN(new_n248));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(new_n212), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g0051(.A(G20), .B1(new_n202), .B2(new_n205), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT8), .B(G58), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  AND3_X1   g0054(.A1(new_n213), .A2(KEYINPUT69), .A3(G33), .ZN(new_n255));
  AOI21_X1  g0055(.A(KEYINPUT69), .B1(new_n213), .B2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n213), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n254), .A2(new_n258), .B1(G150), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n251), .B1(new_n252), .B2(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(KEYINPUT68), .A2(G1), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT68), .A2(G1), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n250), .B1(new_n266), .B2(G20), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G50), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n266), .A2(G13), .A3(G20), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n268), .B1(G50), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n263), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT9), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n271), .B(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT3), .B(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G222), .A2(G1698), .ZN(new_n275));
  INV_X1    g0075(.A(G1698), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(G223), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n274), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G1), .A3(G13), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n278), .B(new_n281), .C1(G77), .C2(new_n274), .ZN(new_n282));
  INV_X1    g0082(.A(G274), .ZN(new_n283));
  AND2_X1   g0083(.A1(G1), .A2(G13), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n283), .B1(new_n284), .B2(new_n279), .ZN(new_n285));
  INV_X1    g0085(.A(G1), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n285), .B(new_n286), .C1(G41), .C2(G45), .ZN(new_n287));
  INV_X1    g0087(.A(G226), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT68), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n286), .ZN(new_n290));
  NAND2_X1  g0090(.A1(KEYINPUT68), .A2(G1), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G41), .A2(G45), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n280), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n282), .B(new_n287), .C1(new_n288), .C2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G190), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n297), .B1(G200), .B2(new_n295), .ZN(new_n298));
  AOI211_X1 g0098(.A(new_n247), .B(new_n248), .C1(new_n273), .C2(new_n298), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n273), .A2(KEYINPUT72), .A3(KEYINPUT10), .A4(new_n298), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G232), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n287), .B1(new_n294), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n274), .A2(G1698), .ZN(new_n306));
  INV_X1    g0106(.A(G87), .ZN(new_n307));
  OAI22_X1  g0107(.A1(new_n306), .A2(new_n288), .B1(new_n259), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT77), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n274), .A2(new_n309), .A3(G223), .A4(new_n276), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT3), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G33), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n311), .A2(new_n313), .A3(G223), .A4(new_n276), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT77), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n308), .B1(new_n310), .B2(new_n315), .ZN(new_n316));
  OAI211_X1 g0116(.A(G179), .B(new_n305), .C1(new_n316), .C2(new_n280), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n311), .A2(new_n313), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n318), .A2(new_n276), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n319), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n315), .A2(new_n310), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n280), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(G169), .B1(new_n322), .B2(new_n304), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n317), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT78), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT78), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n317), .A2(new_n323), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT16), .ZN(new_n328));
  NAND2_X1  g0128(.A1(G58), .A2(G68), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(G58), .A2(G68), .ZN(new_n331));
  OAI21_X1  g0131(.A(G20), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G159), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n332), .B(KEYINPUT75), .C1(new_n333), .C2(new_n260), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT75), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n213), .B1(new_n205), .B2(new_n329), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n260), .A2(new_n333), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT76), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(new_n312), .B2(G33), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n259), .A2(KEYINPUT76), .A3(KEYINPUT3), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n341), .A2(new_n313), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT7), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n344), .A2(G20), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n344), .B1(new_n274), .B2(G20), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n204), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n328), .B1(new_n339), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n318), .A2(KEYINPUT7), .A3(new_n213), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n204), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n339), .A2(new_n351), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n349), .B(new_n250), .C1(new_n352), .C2(new_n328), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n267), .A2(new_n253), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n354), .B1(new_n253), .B2(new_n269), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n325), .A2(new_n327), .A3(new_n357), .ZN(new_n358));
  AND2_X1   g0158(.A1(KEYINPUT79), .A2(KEYINPUT18), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(KEYINPUT79), .A2(KEYINPUT18), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n325), .A2(new_n327), .A3(new_n357), .A4(new_n362), .ZN(new_n363));
  OAI211_X1 g0163(.A(G190), .B(new_n305), .C1(new_n316), .C2(new_n280), .ZN(new_n364));
  OAI21_X1  g0164(.A(G200), .B1(new_n322), .B2(new_n304), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n353), .A2(new_n356), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT17), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AND4_X1   g0168(.A1(new_n353), .A2(new_n356), .A3(new_n364), .A4(new_n365), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT17), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n360), .A2(new_n363), .A3(new_n368), .A4(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n269), .A2(G68), .ZN(new_n373));
  XOR2_X1   g0173(.A(new_n373), .B(KEYINPUT12), .Z(new_n374));
  AOI22_X1  g0174(.A1(new_n261), .A2(G50), .B1(G20), .B2(new_n204), .ZN(new_n375));
  INV_X1    g0175(.A(G77), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n375), .B1(new_n257), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n250), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT11), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n267), .A2(G68), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n377), .A2(KEYINPUT11), .A3(new_n250), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n374), .A2(new_n380), .A3(new_n381), .A4(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G238), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n287), .B1(new_n294), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n303), .A2(G1698), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n274), .B(new_n387), .C1(G226), .C2(G1698), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G33), .A2(G97), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n280), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT13), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT13), .B1(new_n386), .B2(new_n390), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n384), .B1(new_n296), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G200), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n397), .B1(new_n393), .B2(new_n394), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n393), .A2(G179), .A3(new_n394), .ZN(new_n400));
  XNOR2_X1  g0200(.A(new_n400), .B(KEYINPUT74), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n395), .A2(G169), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n402), .A2(KEYINPUT73), .A3(KEYINPUT14), .ZN(new_n403));
  NAND2_X1  g0203(.A1(KEYINPUT73), .A2(KEYINPUT14), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n395), .A2(G169), .A3(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n401), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n399), .B1(new_n406), .B2(new_n383), .ZN(new_n407));
  INV_X1    g0207(.A(new_n271), .ZN(new_n408));
  OR2_X1    g0208(.A1(new_n295), .A2(G179), .ZN(new_n409));
  INV_X1    g0209(.A(G169), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n295), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n408), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n274), .A2(G232), .A3(new_n276), .ZN(new_n413));
  INV_X1    g0213(.A(G107), .ZN(new_n414));
  OAI221_X1 g0214(.A(new_n413), .B1(new_n414), .B2(new_n274), .C1(new_n306), .C2(new_n385), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n280), .B1(new_n415), .B2(KEYINPUT70), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n416), .B1(KEYINPUT70), .B2(new_n415), .ZN(new_n417));
  INV_X1    g0217(.A(new_n294), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(G244), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n419), .A2(new_n287), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n422), .A2(new_n397), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT71), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n253), .B1(new_n424), .B2(new_n260), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n424), .B2(new_n260), .ZN(new_n426));
  XNOR2_X1  g0226(.A(KEYINPUT15), .B(G87), .ZN(new_n427));
  OAI221_X1 g0227(.A(new_n426), .B1(new_n213), .B2(new_n376), .C1(new_n257), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n250), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n269), .A2(G77), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n430), .B1(G77), .B2(new_n267), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n429), .B(new_n431), .C1(new_n421), .C2(new_n296), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n412), .B1(new_n423), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n429), .A2(new_n431), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n422), .B2(G169), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n421), .A2(G179), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n302), .A2(new_n372), .A3(new_n407), .A4(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n269), .A2(G107), .ZN(new_n441));
  XNOR2_X1  g0241(.A(new_n441), .B(KEYINPUT25), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n250), .B1(new_n266), .B2(G33), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n269), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n442), .B1(new_n414), .B2(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n311), .A2(new_n313), .A3(new_n213), .A4(G87), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT22), .ZN(new_n447));
  OR2_X1    g0247(.A1(new_n447), .A2(KEYINPUT88), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n274), .A2(new_n213), .A3(new_n448), .A4(G87), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n213), .A2(G33), .A3(G116), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT23), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n454), .A2(new_n414), .A3(G20), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT23), .B1(new_n213), .B2(G107), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT89), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n453), .B(new_n455), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n456), .A2(new_n457), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT24), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n452), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n461), .B1(new_n452), .B2(new_n460), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n250), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT90), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g0266(.A(KEYINPUT90), .B(new_n250), .C1(new_n462), .C2(new_n463), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n445), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n274), .A2(G257), .A3(G1698), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G294), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n311), .A2(new_n313), .A3(G250), .A4(new_n276), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n281), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT91), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n472), .A2(KEYINPUT91), .A3(new_n281), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n290), .A2(G45), .A3(new_n291), .ZN(new_n477));
  AND2_X1   g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  NOR2_X1   g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(G264), .B(new_n280), .C1(new_n477), .C2(new_n480), .ZN(new_n481));
  XNOR2_X1  g0281(.A(KEYINPUT5), .B(G41), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n285), .A2(new_n266), .A3(new_n482), .A4(G45), .ZN(new_n483));
  AND2_X1   g0283(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n475), .A2(new_n476), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n473), .A2(new_n483), .A3(new_n481), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n485), .A2(G169), .B1(new_n487), .B2(G179), .ZN(new_n488));
  OR2_X1    g0288(.A1(new_n468), .A2(new_n488), .ZN(new_n489));
  OAI22_X1  g0289(.A1(new_n485), .A2(G190), .B1(new_n487), .B2(G200), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n468), .A2(new_n490), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n274), .A2(G244), .A3(G1698), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G116), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n311), .A2(new_n313), .A3(G238), .A4(new_n276), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n281), .ZN(new_n497));
  AND2_X1   g0297(.A1(G33), .A2(G41), .ZN(new_n498));
  OAI21_X1  g0298(.A(G274), .B1(new_n498), .B2(new_n212), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n499), .A2(G45), .A3(new_n266), .ZN(new_n500));
  OAI21_X1  g0300(.A(G250), .B1(new_n498), .B2(new_n212), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n477), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT82), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n500), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n503), .B1(new_n500), .B2(new_n502), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n497), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n410), .ZN(new_n507));
  INV_X1    g0307(.A(G179), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n477), .A2(new_n285), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n266), .A2(G45), .B1(new_n280), .B2(G250), .ZN(new_n510));
  OAI21_X1  g0310(.A(KEYINPUT82), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n500), .A2(new_n502), .A3(new_n503), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n511), .A2(new_n512), .B1(new_n281), .B2(new_n496), .ZN(new_n513));
  INV_X1    g0313(.A(new_n427), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n269), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(G97), .B1(new_n255), .B2(new_n256), .ZN(new_n516));
  OR2_X1    g0316(.A1(KEYINPUT83), .A2(KEYINPUT19), .ZN(new_n517));
  NAND2_X1  g0317(.A1(KEYINPUT83), .A2(KEYINPUT19), .ZN(new_n518));
  AND2_X1   g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(KEYINPUT84), .A2(G87), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(G97), .A2(G107), .ZN(new_n523));
  NAND2_X1  g0323(.A1(KEYINPUT84), .A2(G87), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n389), .B1(new_n517), .B2(new_n518), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n525), .B1(new_n526), .B2(G20), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n274), .A2(new_n213), .A3(G68), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n520), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n515), .B1(new_n529), .B2(new_n250), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n443), .A2(new_n269), .A3(new_n514), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n508), .A2(new_n513), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n497), .B(G190), .C1(new_n504), .C2(new_n505), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT85), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n444), .B2(new_n307), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n443), .A2(new_n269), .A3(KEYINPUT85), .A4(G87), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n533), .A2(new_n537), .A3(new_n530), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n506), .A2(G200), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n507), .A2(new_n532), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n443), .A2(G116), .A3(new_n269), .ZN(new_n541));
  INV_X1    g0341(.A(G116), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n266), .A2(G13), .A3(G20), .A4(new_n542), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n249), .A2(new_n212), .B1(G20), .B2(new_n542), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G33), .A2(G283), .ZN(new_n545));
  INV_X1    g0345(.A(G97), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n545), .B(new_n213), .C1(G33), .C2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT20), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n544), .A2(KEYINPUT20), .A3(new_n547), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n541), .B(new_n543), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(G270), .B(new_n280), .C1(new_n477), .C2(new_n480), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n551), .A2(new_n483), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n312), .A2(G33), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n554));
  OAI21_X1  g0354(.A(G303), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n311), .A2(new_n313), .A3(G264), .A4(G1698), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n311), .A2(new_n313), .A3(G257), .A4(new_n276), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n281), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n552), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n550), .B1(new_n560), .B2(G200), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT87), .ZN(new_n562));
  OR2_X1    g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n560), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G190), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n561), .A2(new_n562), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n563), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n560), .A2(new_n550), .A3(G169), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT21), .ZN(new_n569));
  OAI21_X1  g0369(.A(KEYINPUT86), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n410), .B1(new_n552), .B2(new_n559), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT86), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT21), .A4(new_n550), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n559), .A2(G179), .A3(new_n483), .A4(new_n551), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n568), .A2(new_n569), .B1(new_n576), .B2(new_n550), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n567), .A2(new_n574), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT81), .ZN(new_n579));
  OAI211_X1 g0379(.A(G257), .B(new_n280), .C1(new_n477), .C2(new_n480), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n580), .A2(new_n483), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n311), .A2(new_n313), .A3(G244), .A4(new_n276), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT4), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n545), .ZN(new_n585));
  NAND2_X1  g0385(.A1(G250), .A2(G1698), .ZN(new_n586));
  NAND2_X1  g0386(.A1(KEYINPUT4), .A2(G244), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n586), .B1(new_n587), .B2(G1698), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n585), .B1(new_n274), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n281), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n581), .A2(new_n591), .A3(new_n508), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n346), .A2(new_n347), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(G107), .ZN(new_n594));
  XNOR2_X1  g0394(.A(G97), .B(G107), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT6), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n596), .A2(new_n546), .A3(G107), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n600), .A2(G20), .B1(G77), .B2(new_n261), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n251), .B1(new_n594), .B2(new_n601), .ZN(new_n602));
  OR2_X1    g0402(.A1(new_n269), .A2(G97), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n443), .A2(G97), .A3(new_n269), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n592), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT80), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n581), .A2(new_n591), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n280), .B1(new_n584), .B2(new_n589), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n580), .A2(new_n483), .ZN(new_n610));
  OAI21_X1  g0410(.A(KEYINPUT80), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(G169), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n579), .B1(new_n606), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n602), .A2(new_n605), .ZN(new_n614));
  OAI21_X1  g0414(.A(G200), .B1(new_n609), .B2(new_n610), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n608), .A2(new_n611), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n614), .B(new_n615), .C1(new_n296), .C2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n607), .B1(new_n581), .B2(new_n591), .ZN(new_n618));
  NOR3_X1   g0418(.A1(new_n609), .A2(new_n610), .A3(KEYINPUT80), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n410), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n598), .B1(new_n596), .B2(new_n595), .ZN(new_n621));
  OAI22_X1  g0421(.A1(new_n621), .A2(new_n213), .B1(new_n376), .B2(new_n260), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n414), .B1(new_n346), .B2(new_n347), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n250), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n605), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n609), .A2(new_n610), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n624), .A2(new_n625), .B1(new_n626), .B2(new_n508), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n620), .A2(KEYINPUT81), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n613), .A2(new_n617), .A3(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n578), .A2(new_n629), .ZN(new_n630));
  AND4_X1   g0430(.A1(new_n440), .A2(new_n492), .A3(new_n540), .A4(new_n630), .ZN(G372));
  INV_X1    g0431(.A(new_n412), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n302), .A2(KEYINPUT95), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT95), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n299), .B2(new_n301), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n353), .A2(new_n356), .B1(new_n317), .B2(new_n323), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT18), .ZN(new_n638));
  XNOR2_X1  g0438(.A(new_n637), .B(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n399), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n641), .A2(new_n437), .B1(new_n406), .B2(new_n383), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n370), .A2(new_n368), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT94), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n636), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n632), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(KEYINPUT92), .B1(new_n504), .B2(new_n505), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT92), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n511), .A2(new_n650), .A3(new_n512), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n649), .A2(new_n497), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n410), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n532), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n574), .B(new_n577), .C1(new_n468), .C2(new_n488), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n652), .A2(G200), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n538), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT93), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n654), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n658), .B1(new_n654), .B2(new_n657), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n629), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n491), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n654), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n606), .A2(new_n612), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n665), .B(new_n666), .C1(new_n659), .C2(new_n660), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n613), .A2(new_n628), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n540), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT26), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n664), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n440), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n648), .A2(new_n673), .ZN(G369));
  AND2_X1   g0474(.A1(new_n574), .A2(new_n577), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n213), .A2(G13), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n266), .A2(new_n676), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G213), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n550), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n675), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n675), .A2(new_n567), .A3(new_n683), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G330), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n492), .ZN(new_n689));
  INV_X1    g0489(.A(new_n682), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n468), .A2(new_n690), .ZN(new_n691));
  OAI22_X1  g0491(.A1(new_n689), .A2(new_n691), .B1(new_n489), .B2(new_n690), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n489), .A2(new_n682), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n675), .A2(new_n682), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n694), .B1(new_n492), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n693), .A2(new_n696), .ZN(G399));
  INV_X1    g0497(.A(new_n209), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(G41), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n525), .A2(G116), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(G1), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n215), .B2(new_n700), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT28), .ZN(new_n704));
  OAI211_X1 g0504(.A(KEYINPUT26), .B(new_n666), .C1(new_n659), .C2(new_n660), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT100), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n706), .B1(new_n669), .B2(new_n665), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n529), .A2(new_n250), .ZN(new_n709));
  INV_X1    g0509(.A(new_n515), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(new_n710), .A3(new_n531), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n497), .B(new_n508), .C1(new_n504), .C2(new_n505), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n713), .B1(new_n410), .B2(new_n652), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n533), .A2(new_n537), .A3(new_n530), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n715), .B1(G200), .B2(new_n652), .ZN(new_n716));
  OAI21_X1  g0516(.A(KEYINPUT93), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n654), .A2(new_n657), .A3(new_n658), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n719), .A2(new_n491), .A3(new_n662), .A4(new_n655), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n719), .A2(new_n706), .A3(KEYINPUT26), .A4(new_n666), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n708), .A2(new_n654), .A3(new_n720), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n690), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT29), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n672), .A2(new_n690), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n724), .B1(new_n725), .B2(KEYINPUT29), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n473), .A2(new_n481), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n506), .A2(new_n575), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n618), .A2(new_n619), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n728), .A2(new_n729), .A3(KEYINPUT30), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT97), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n728), .A2(new_n729), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT30), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n728), .A2(new_n729), .A3(KEYINPUT97), .A4(KEYINPUT30), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n564), .A2(G179), .A3(new_n626), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(new_n486), .A3(new_n652), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n732), .A2(new_n735), .A3(new_n736), .A4(new_n738), .ZN(new_n739));
  XOR2_X1   g0539(.A(KEYINPUT96), .B(KEYINPUT31), .Z(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AND3_X1   g0541(.A1(new_n739), .A2(new_n682), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(KEYINPUT31), .B1(new_n739), .B2(new_n682), .ZN(new_n743));
  OAI21_X1  g0543(.A(KEYINPUT98), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n739), .A2(new_n682), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT31), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT98), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n739), .A2(new_n682), .A3(new_n741), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n492), .A2(new_n630), .A3(new_n540), .A4(new_n690), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n744), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT99), .ZN(new_n753));
  AND3_X1   g0553(.A1(new_n752), .A2(new_n753), .A3(G330), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n753), .B1(new_n752), .B2(G330), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n726), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n704), .B1(new_n756), .B2(G1), .ZN(G364));
  XNOR2_X1  g0557(.A(new_n687), .B(KEYINPUT101), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n286), .B1(new_n676), .B2(G45), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n699), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n758), .B(new_n762), .C1(G330), .C2(new_n686), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G13), .A2(G33), .ZN(new_n764));
  XOR2_X1   g0564(.A(new_n764), .B(KEYINPUT102), .Z(new_n765));
  OR2_X1    g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  XOR2_X1   g0566(.A(new_n766), .B(KEYINPUT103), .Z(new_n767));
  AOI21_X1  g0567(.A(new_n212), .B1(G20), .B2(new_n410), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n274), .A2(new_n209), .ZN(new_n771));
  INV_X1    g0571(.A(G355), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n771), .A2(new_n772), .B1(G116), .B2(new_n209), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n240), .A2(G45), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n318), .A2(new_n209), .ZN(new_n775));
  INV_X1    g0575(.A(G45), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n775), .B1(new_n776), .B2(new_n216), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n773), .B1(new_n774), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n761), .B1(new_n770), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n213), .A2(G179), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n780), .A2(G190), .A3(G200), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT105), .Z(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G303), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n213), .A2(new_n508), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G190), .A2(G200), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n780), .A2(new_n785), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI22_X1  g0589(.A1(G311), .A2(new_n787), .B1(new_n789), .B2(G329), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n784), .A2(G190), .A3(new_n397), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n274), .B1(new_n792), .B2(G322), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n784), .A2(G200), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n296), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n780), .A2(new_n296), .A3(G200), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n796), .A2(G326), .B1(new_n798), .B2(G283), .ZN(new_n799));
  NOR3_X1   g0599(.A1(new_n296), .A2(G179), .A3(G200), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n213), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n795), .A2(G190), .ZN(new_n803));
  XNOR2_X1  g0603(.A(KEYINPUT33), .B(G317), .ZN(new_n804));
  AOI22_X1  g0604(.A1(G294), .A2(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n783), .A2(new_n794), .A3(new_n799), .A4(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT106), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n797), .A2(new_n414), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n522), .A2(new_n524), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n810), .A2(new_n781), .B1(new_n801), .B2(new_n546), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n809), .B(new_n811), .C1(G50), .C2(new_n796), .ZN(new_n812));
  XNOR2_X1  g0612(.A(KEYINPUT104), .B(G159), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n789), .A2(new_n813), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n814), .A2(KEYINPUT32), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n814), .A2(KEYINPUT32), .B1(new_n803), .B2(G68), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n274), .B1(new_n791), .B2(new_n203), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(G77), .B2(new_n787), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n812), .A2(new_n815), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n806), .A2(new_n807), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n808), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n779), .B1(new_n821), .B2(new_n768), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n686), .B2(new_n767), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n763), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(G396));
  NOR2_X1   g0625(.A1(new_n754), .A2(new_n755), .ZN(new_n826));
  INV_X1    g0626(.A(new_n437), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n434), .A2(new_n682), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n423), .B2(new_n432), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NOR3_X1   g0630(.A1(new_n435), .A2(new_n436), .A3(new_n682), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n725), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n831), .B1(new_n827), .B2(new_n829), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n690), .B(new_n835), .C1(new_n664), .C2(new_n671), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n761), .B1(new_n826), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n826), .B2(new_n837), .ZN(new_n839));
  INV_X1    g0639(.A(new_n803), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n840), .A2(KEYINPUT107), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n840), .A2(KEYINPUT107), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n844), .A2(G283), .B1(G116), .B2(new_n787), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n845), .A2(KEYINPUT108), .B1(G303), .B2(new_n796), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(KEYINPUT108), .B2(new_n845), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT109), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n782), .A2(G107), .ZN(new_n849));
  INV_X1    g0649(.A(G294), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n318), .B1(new_n791), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(G311), .B2(new_n789), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n797), .A2(new_n307), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(G97), .B2(new_n802), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n849), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n792), .A2(G143), .B1(new_n787), .B2(new_n813), .ZN(new_n856));
  INV_X1    g0656(.A(new_n796), .ZN(new_n857));
  INV_X1    g0657(.A(G137), .ZN(new_n858));
  INV_X1    g0658(.A(G150), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n856), .B1(new_n857), .B2(new_n858), .C1(new_n859), .C2(new_n840), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT34), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n860), .A2(new_n861), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n782), .A2(G50), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n797), .A2(new_n204), .ZN(new_n865));
  INV_X1    g0665(.A(G132), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n274), .B1(new_n788), .B2(new_n866), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n865), .B(new_n867), .C1(G58), .C2(new_n802), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n863), .A2(new_n864), .A3(new_n868), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n848), .A2(new_n855), .B1(new_n862), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n768), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n768), .A2(new_n764), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n762), .B1(new_n376), .B2(new_n872), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n871), .B(new_n873), .C1(new_n765), .C2(new_n835), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n839), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(G384));
  OR2_X1    g0676(.A1(new_n600), .A2(KEYINPUT35), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n600), .A2(KEYINPUT35), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n877), .A2(G116), .A3(new_n214), .A4(new_n878), .ZN(new_n879));
  XOR2_X1   g0679(.A(new_n879), .B(KEYINPUT36), .Z(new_n880));
  NAND3_X1  g0680(.A1(new_n216), .A2(G77), .A3(new_n329), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n201), .A2(G68), .ZN(new_n882));
  AOI211_X1 g0682(.A(G13), .B(new_n266), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT39), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n680), .B1(new_n353), .B2(new_n356), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n369), .A2(new_n637), .A3(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT110), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n886), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n358), .A2(new_n888), .A3(new_n366), .A4(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n637), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n892), .A2(new_n890), .A3(new_n366), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT110), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n893), .A2(new_n894), .A3(KEYINPUT37), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n889), .A2(new_n891), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n886), .B1(new_n639), .B2(new_n643), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT38), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT38), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n352), .A2(new_n328), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n339), .A2(new_n351), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n251), .B1(new_n901), .B2(KEYINPUT16), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n355), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n317), .A2(new_n323), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n366), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n903), .A2(new_n680), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT37), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AOI221_X4 g0707(.A(new_n899), .B1(new_n907), .B2(new_n891), .C1(new_n371), .C2(new_n906), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n885), .B1(new_n898), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n371), .A2(new_n906), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n907), .A2(new_n891), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n899), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n910), .A2(KEYINPUT38), .A3(new_n911), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n913), .A2(KEYINPUT39), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n909), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n406), .A2(new_n383), .A3(new_n690), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n384), .A2(new_n690), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n407), .B(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n922), .B1(new_n836), .B2(new_n832), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n913), .A2(new_n914), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n923), .A2(new_n924), .B1(new_n639), .B2(new_n680), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n920), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n726), .A2(new_n440), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n648), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n926), .B(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(G330), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n745), .A2(new_n746), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(new_n740), .B2(new_n745), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n751), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n407), .B1(new_n384), .B2(new_n690), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n383), .B(new_n682), .C1(new_n406), .C2(new_n399), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n833), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n898), .A2(new_n908), .ZN(new_n938));
  OAI21_X1  g0738(.A(KEYINPUT40), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT40), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n924), .A2(new_n940), .A3(new_n933), .A4(new_n936), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n439), .B1(new_n932), .B2(new_n751), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n930), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n943), .B2(new_n942), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n929), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n266), .B2(new_n676), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n929), .A2(new_n945), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n884), .B1(new_n947), .B2(new_n948), .ZN(G367));
  NAND2_X1  g0749(.A1(new_n537), .A2(new_n530), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n682), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n654), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(new_n719), .B2(new_n951), .ZN(new_n953));
  INV_X1    g0753(.A(new_n767), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n236), .A2(new_n775), .B1(new_n209), .B2(new_n427), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n761), .B1(new_n770), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n844), .A2(new_n813), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n201), .A2(new_n786), .B1(new_n788), .B2(new_n858), .ZN(new_n959));
  AOI211_X1 g0759(.A(new_n318), .B(new_n959), .C1(G150), .C2(new_n792), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n801), .A2(new_n204), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(G143), .B2(new_n796), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n797), .A2(new_n376), .ZN(new_n963));
  INV_X1    g0763(.A(new_n781), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n963), .B1(G58), .B2(new_n964), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n958), .A2(new_n960), .A3(new_n962), .A4(new_n965), .ZN(new_n966));
  AOI22_X1  g0766(.A1(G283), .A2(new_n787), .B1(new_n789), .B2(G317), .ZN(new_n967));
  INV_X1    g0767(.A(G303), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n967), .B(new_n318), .C1(new_n968), .C2(new_n791), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n796), .A2(G311), .B1(new_n798), .B2(G97), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n414), .B2(new_n801), .ZN(new_n971));
  AOI21_X1  g0771(.A(KEYINPUT46), .B1(new_n964), .B2(G116), .ZN(new_n972));
  NOR3_X1   g0772(.A1(new_n969), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n782), .A2(KEYINPUT46), .A3(G116), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n973), .B(new_n974), .C1(new_n850), .C2(new_n843), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n966), .A2(new_n975), .ZN(new_n976));
  XOR2_X1   g0776(.A(KEYINPUT114), .B(KEYINPUT47), .Z(new_n977));
  XNOR2_X1  g0777(.A(new_n976), .B(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n957), .B1(new_n978), .B2(new_n768), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n955), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT43), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n953), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n662), .B1(new_n614), .B2(new_n690), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n666), .A2(new_n682), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n613), .B(new_n628), .C1(new_n986), .C2(new_n489), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n987), .A2(KEYINPUT111), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(KEYINPUT111), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n988), .A2(new_n690), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n492), .A2(new_n695), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n986), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT42), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n982), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n953), .A2(new_n981), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n693), .A2(new_n986), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n994), .A2(new_n995), .ZN(new_n999));
  AND3_X1   g0799(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n998), .B1(new_n997), .B2(new_n999), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n991), .B1(new_n692), .B2(new_n695), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1003), .A2(new_n687), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT112), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AND2_X1   g0806(.A1(new_n758), .A2(new_n1003), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n756), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n696), .A2(new_n985), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT44), .Z(new_n1012));
  NAND2_X1  g0812(.A1(new_n696), .A2(new_n985), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT45), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(new_n693), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n756), .B1(new_n1010), .B2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n699), .B(KEYINPUT41), .Z(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n760), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(KEYINPUT113), .B1(new_n1002), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1020), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT113), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n980), .B1(new_n1021), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(G387));
  OR2_X1    g0827(.A1(new_n692), .A2(new_n767), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n233), .A2(new_n776), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n1029), .A2(new_n775), .B1(new_n701), .B2(new_n771), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n253), .A2(G50), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT50), .ZN(new_n1032));
  AOI21_X1  g0832(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1032), .A2(new_n701), .A3(new_n1033), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n1030), .A2(new_n1034), .B1(new_n414), .B2(new_n698), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n761), .B1(new_n1035), .B2(new_n770), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n786), .A2(new_n204), .B1(new_n788), .B2(new_n859), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n318), .B(new_n1037), .C1(G50), .C2(new_n792), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n964), .A2(G77), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n801), .A2(new_n427), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n254), .B2(new_n803), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n796), .A2(G159), .B1(new_n798), .B2(G97), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1038), .A2(new_n1039), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n274), .B1(new_n789), .B2(G326), .ZN(new_n1044));
  INV_X1    g0844(.A(G283), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n801), .A2(new_n1045), .B1(new_n781), .B2(new_n850), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT115), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n792), .A2(G317), .B1(new_n787), .B2(G303), .ZN(new_n1048));
  INV_X1    g0848(.A(G322), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1048), .B1(new_n1049), .B2(new_n857), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n844), .B2(G311), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1047), .B1(new_n1051), .B2(KEYINPUT48), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT116), .Z(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(KEYINPUT48), .B2(new_n1051), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT49), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1044), .B1(new_n542), .B2(new_n797), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1043), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1036), .B1(new_n1058), .B2(new_n768), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n1009), .A2(new_n760), .B1(new_n1028), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1010), .A2(new_n699), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1009), .A2(new_n756), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1060), .B1(new_n1061), .B2(new_n1062), .ZN(G393));
  OAI22_X1  g0863(.A1(new_n243), .A2(new_n775), .B1(new_n546), .B2(new_n209), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n761), .B1(new_n770), .B2(new_n1064), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(G317), .A2(new_n796), .B1(new_n792), .B2(G311), .ZN(new_n1066));
  XOR2_X1   g0866(.A(KEYINPUT117), .B(KEYINPUT52), .Z(new_n1067));
  AOI22_X1  g0867(.A1(new_n844), .A2(G303), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n318), .B1(new_n786), .B2(new_n850), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(G322), .B2(new_n789), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n809), .B1(G116), .B2(new_n802), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(new_n1045), .C2(new_n781), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G150), .A2(new_n796), .B1(new_n792), .B2(G159), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT51), .ZN(new_n1075));
  INV_X1    g0875(.A(G143), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n274), .B1(new_n788), .B2(new_n1076), .C1(new_n253), .C2(new_n786), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n801), .A2(new_n376), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n853), .B(new_n1079), .C1(G68), .C2(new_n964), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1078), .B(new_n1080), .C1(new_n843), .C2(new_n201), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n1069), .A2(new_n1073), .B1(new_n1075), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1065), .B1(new_n1082), .B2(new_n768), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n985), .B2(new_n767), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n1016), .B2(new_n759), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1010), .A2(new_n1016), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(KEYINPUT118), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT118), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1010), .A2(new_n1016), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1010), .A2(new_n1016), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1091), .A2(new_n700), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(KEYINPUT119), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT119), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1090), .A2(new_n1095), .A3(new_n1092), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1085), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(G390));
  INV_X1    g0898(.A(new_n922), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n835), .B(new_n1099), .C1(new_n754), .C2(new_n755), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n722), .A2(new_n690), .A3(new_n830), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n832), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n1099), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n918), .B1(new_n898), .B2(new_n908), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n916), .B1(new_n919), .B2(new_n923), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1100), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n930), .B1(new_n932), .B2(new_n751), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n1109), .A2(new_n936), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n836), .A2(new_n832), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n1099), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1112), .A2(new_n918), .B1(new_n909), .B2(new_n915), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1104), .B1(new_n1102), .B2(new_n1099), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1110), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AND2_X1   g0915(.A1(new_n1108), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n760), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n844), .A2(G107), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n791), .A2(new_n542), .B1(new_n786), .B2(new_n546), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n274), .B(new_n1119), .C1(G294), .C2(new_n789), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n865), .B(new_n1079), .C1(G283), .C2(new_n796), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n782), .A2(G87), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1118), .A2(new_n1120), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n844), .A2(G137), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT54), .B(G143), .ZN(new_n1125));
  INV_X1    g0925(.A(G125), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n786), .A2(new_n1125), .B1(new_n788), .B2(new_n1126), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n318), .B(new_n1127), .C1(G132), .C2(new_n792), .ZN(new_n1128));
  INV_X1    g0928(.A(G128), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n857), .A2(new_n1129), .B1(new_n333), .B2(new_n801), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n202), .B2(new_n798), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n781), .A2(new_n859), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT53), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1124), .A2(new_n1128), .A3(new_n1131), .A4(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n769), .B1(new_n1123), .B2(new_n1134), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n762), .B(new_n1135), .C1(new_n253), .C2(new_n872), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n917), .B2(new_n765), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1117), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(KEYINPUT120), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1109), .A2(new_n835), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1102), .B1(new_n1141), .B2(new_n922), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1100), .A2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n835), .B1(new_n754), .B2(new_n755), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1110), .B1(new_n1144), .B2(new_n922), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1111), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1143), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1109), .A2(new_n440), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n927), .A2(new_n648), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1116), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1116), .A2(new_n1147), .A3(new_n1150), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1153), .A2(new_n699), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT120), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1138), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1140), .A2(new_n1155), .A3(new_n1157), .ZN(G378));
  NAND2_X1  g0958(.A1(new_n942), .A2(G330), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1159), .A2(new_n920), .A3(new_n925), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n930), .B1(new_n939), .B2(new_n941), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n926), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n633), .A2(new_n412), .A3(new_n635), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n271), .A2(new_n680), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT122), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1164), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n633), .A2(new_n412), .A3(new_n635), .A4(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1165), .A2(new_n1166), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1166), .B1(new_n1165), .B2(new_n1168), .ZN(new_n1171));
  XOR2_X1   g0971(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(new_n1170), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1165), .A2(new_n1168), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(KEYINPUT122), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1172), .B1(new_n1176), .B2(new_n1169), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1174), .A2(new_n1177), .ZN(new_n1178));
  AND3_X1   g0978(.A1(new_n1160), .A2(new_n1162), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1178), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  OR2_X1    g0981(.A1(new_n1178), .A2(new_n765), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n872), .A2(new_n201), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(G33), .A2(G41), .ZN(new_n1184));
  INV_X1    g0984(.A(G41), .ZN(new_n1185));
  AOI211_X1 g0985(.A(G50), .B(new_n1184), .C1(new_n318), .C2(new_n1185), .ZN(new_n1186));
  AOI211_X1 g0986(.A(G41), .B(new_n274), .C1(new_n789), .C2(G283), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1187), .B(new_n1039), .C1(new_n203), .C2(new_n797), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT121), .Z(new_n1189));
  OAI22_X1  g0989(.A1(new_n791), .A2(new_n414), .B1(new_n786), .B2(new_n427), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n546), .A2(new_n840), .B1(new_n857), .B2(new_n542), .ZN(new_n1191));
  NOR4_X1   g0991(.A1(new_n1189), .A2(new_n961), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1186), .B1(new_n1192), .B2(KEYINPUT58), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n1126), .A2(new_n857), .B1(new_n840), .B2(new_n866), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n792), .A2(G128), .B1(new_n787), .B2(G137), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n781), .B2(new_n1125), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1194), .B(new_n1196), .C1(G150), .C2(new_n802), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1198), .A2(KEYINPUT59), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(KEYINPUT59), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n798), .A2(new_n813), .ZN(new_n1201));
  AOI211_X1 g1001(.A(G33), .B(G41), .C1(new_n789), .C2(G124), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1193), .B1(KEYINPUT58), .B2(new_n1192), .C1(new_n1199), .C2(new_n1203), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n762), .B(new_n1183), .C1(new_n1204), .C2(new_n768), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1181), .A2(new_n760), .B1(new_n1182), .B2(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1149), .B(KEYINPUT123), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1154), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT124), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1154), .A2(KEYINPUT124), .A3(new_n1207), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(KEYINPUT57), .B1(new_n1212), .B2(new_n1181), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT57), .ZN(new_n1214));
  NOR3_X1   g1014(.A1(new_n1179), .A2(new_n1180), .A3(new_n1214), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n1154), .A2(KEYINPUT124), .A3(new_n1207), .ZN(new_n1216));
  AOI21_X1  g1016(.A(KEYINPUT124), .B1(new_n1154), .B2(new_n1207), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1215), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n699), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1206), .B1(new_n1213), .B2(new_n1219), .ZN(G375));
  OR2_X1    g1020(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1221), .A2(new_n1019), .A3(new_n1151), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n922), .A2(new_n764), .ZN(new_n1223));
  NOR3_X1   g1023(.A1(new_n768), .A2(G68), .A3(new_n764), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n844), .A2(G116), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n791), .A2(new_n1045), .B1(new_n786), .B2(new_n414), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n274), .B(new_n1226), .C1(G303), .C2(new_n789), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n963), .B(new_n1040), .C1(G294), .C2(new_n796), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n782), .A2(G97), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1225), .A2(new_n1227), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(G132), .A2(new_n796), .B1(new_n792), .B2(G137), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n843), .B2(new_n1125), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT125), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n782), .A2(G159), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n797), .A2(new_n203), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n274), .B1(new_n788), .B2(new_n1129), .C1(new_n859), .C2(new_n786), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n1236), .B(new_n1237), .C1(G50), .C2(new_n802), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1234), .A2(new_n1235), .A3(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1230), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n762), .B(new_n1224), .C1(new_n1241), .C2(new_n768), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n1147), .A2(new_n760), .B1(new_n1223), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1222), .A2(new_n1243), .ZN(G381));
  OR2_X1    g1044(.A1(G393), .A2(G396), .ZN(new_n1245));
  NOR4_X1   g1045(.A1(G390), .A2(G384), .A3(G381), .A4(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(G375), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1155), .A2(new_n1139), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1246), .A2(new_n1026), .A3(new_n1247), .A4(new_n1248), .ZN(G407));
  NAND4_X1  g1049(.A1(new_n1247), .A2(G213), .A3(new_n681), .A4(new_n1248), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(G407), .A2(G213), .A3(new_n1250), .ZN(G409));
  NAND2_X1  g1051(.A1(G387), .A2(new_n1097), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G390), .A2(new_n1026), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(G393), .B(new_n824), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT61), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1252), .A2(new_n1255), .A3(new_n1253), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  OAI211_X1 g1060(.A(G378), .B(new_n1206), .C1(new_n1213), .C2(new_n1219), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1019), .B(new_n1181), .C1(new_n1216), .C2(new_n1217), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1206), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1248), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1261), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n681), .A2(G213), .ZN(new_n1266));
  AND2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1151), .A2(KEYINPUT60), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1268), .A2(new_n1221), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n699), .B1(new_n1268), .B2(new_n1221), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1243), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n875), .ZN(new_n1272));
  OAI211_X1 g1072(.A(G384), .B(new_n1243), .C1(new_n1269), .C2(new_n1270), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT63), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1260), .B1(new_n1267), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1265), .A2(KEYINPUT126), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1274), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT126), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1261), .A2(new_n1280), .A3(new_n1264), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1278), .A2(new_n1266), .A3(new_n1279), .A4(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1275), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1278), .A2(new_n1266), .A3(new_n1281), .ZN(new_n1284));
  AND3_X1   g1084(.A1(new_n681), .A2(G213), .A3(G2897), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1274), .B(new_n1285), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1277), .B(new_n1283), .C1(new_n1284), .C2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1258), .B1(new_n1267), .B2(new_n1286), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT62), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1282), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1267), .A2(KEYINPUT62), .A3(new_n1279), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1289), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT127), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1288), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  AOI211_X1 g1095(.A(KEYINPUT127), .B(new_n1289), .C1(new_n1291), .C2(new_n1292), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1287), .B1(new_n1295), .B2(new_n1296), .ZN(G405));
  INV_X1    g1097(.A(new_n1261), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1298), .B1(G375), .B2(new_n1248), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1299), .B(new_n1274), .ZN(new_n1300));
  XNOR2_X1  g1100(.A(new_n1300), .B(new_n1288), .ZN(G402));
endmodule


