//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 1 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 0 1 1 1 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n841, new_n842,
    new_n843, new_n844, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961;
  AND2_X1   g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT29), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G169gat), .ZN(new_n205));
  INV_X1    g004(.A(G176gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AND2_X1   g006(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n208));
  NOR2_X1   g007(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT66), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n207), .B(KEYINPUT66), .C1(new_n208), .C2(new_n209), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n215), .B(KEYINPUT24), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n216), .B1(G183gat), .B2(G190gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n218), .B(KEYINPUT67), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(KEYINPUT64), .B(G176gat), .Z(new_n221));
  NAND3_X1  g020(.A1(new_n221), .A2(KEYINPUT23), .A3(new_n205), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n214), .A2(new_n217), .A3(new_n220), .A4(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT25), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT68), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n207), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT68), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT23), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT69), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(new_n232), .A3(new_n220), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT23), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n234), .B1(new_n227), .B2(new_n229), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT69), .B1(new_n235), .B2(new_n219), .ZN(new_n236));
  OR2_X1    g035(.A1(KEYINPUT70), .A2(G183gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(KEYINPUT70), .A2(G183gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(G190gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n224), .B1(new_n241), .B2(new_n216), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n233), .A2(new_n236), .A3(new_n214), .A4(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n225), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n237), .A2(KEYINPUT27), .A3(new_n238), .ZN(new_n245));
  NOR2_X1   g044(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(G190gat), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(KEYINPUT71), .B1(new_n248), .B2(KEYINPUT28), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT71), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT28), .ZN(new_n251));
  AND2_X1   g050(.A1(KEYINPUT70), .A2(G183gat), .ZN(new_n252));
  NOR2_X1   g051(.A1(KEYINPUT70), .A2(G183gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n246), .B1(new_n254), .B2(KEYINPUT27), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n250), .B(new_n251), .C1(new_n255), .C2(G190gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT27), .B(G183gat), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n257), .A2(KEYINPUT28), .A3(new_n240), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n249), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n207), .A2(KEYINPUT26), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT26), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n261), .B1(new_n230), .B2(new_n262), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n263), .A2(new_n220), .B1(G183gat), .B2(G190gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n204), .B1(new_n244), .B2(new_n265), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n236), .A2(new_n214), .ZN(new_n267));
  NOR3_X1   g066(.A1(new_n235), .A2(KEYINPUT69), .A3(new_n219), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n241), .A2(new_n216), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT25), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n267), .A2(new_n271), .B1(new_n223), .B2(new_n224), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n265), .A2(KEYINPUT72), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT72), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n259), .A2(new_n274), .A3(new_n264), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n272), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n266), .B1(new_n276), .B2(new_n202), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT22), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT77), .B(G211gat), .ZN(new_n279));
  INV_X1    g078(.A(G218gat), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G197gat), .B(G204gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G211gat), .B(G218gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(KEYINPUT78), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n281), .B(new_n282), .C1(KEYINPUT78), .C2(new_n284), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n286), .A2(KEYINPUT79), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT79), .B1(new_n286), .B2(new_n287), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT80), .B1(new_n277), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n244), .A2(new_n265), .A3(new_n202), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n294), .B(new_n292), .C1(new_n276), .C2(new_n204), .ZN(new_n295));
  AND3_X1   g094(.A1(new_n259), .A2(new_n274), .A3(new_n264), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n274), .B1(new_n259), .B2(new_n264), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n244), .B(new_n202), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n244), .A2(new_n265), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(new_n203), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT80), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(new_n302), .A3(new_n291), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n293), .A2(new_n295), .A3(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G8gat), .B(G36gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(G64gat), .B(G92gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n307), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n293), .A2(new_n295), .A3(new_n303), .A4(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(KEYINPUT30), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n302), .B1(new_n301), .B2(new_n291), .ZN(new_n312));
  AOI211_X1 g111(.A(KEYINPUT80), .B(new_n292), .C1(new_n298), .C2(new_n300), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT30), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n314), .A2(new_n315), .A3(new_n295), .A4(new_n309), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G78gat), .B(G106gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n319), .B(G22gat), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(KEYINPUT31), .B(G50gat), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G228gat), .ZN(new_n324));
  INV_X1    g123(.A(G233gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n286), .A2(new_n287), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT79), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT29), .ZN(new_n331));
  XOR2_X1   g130(.A(G141gat), .B(G148gat), .Z(new_n332));
  INV_X1    g131(.A(G155gat), .ZN(new_n333));
  INV_X1    g132(.A(G162gat), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT2), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G155gat), .B(G162gat), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT3), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n332), .A2(new_n335), .A3(new_n337), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n330), .A2(new_n288), .B1(new_n331), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n339), .A2(new_n341), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT29), .B1(new_n283), .B2(new_n284), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n346), .B1(new_n284), .B2(new_n283), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n345), .B1(new_n347), .B2(new_n340), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n327), .B1(new_n343), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT85), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI211_X1 g150(.A(KEYINPUT85), .B(new_n327), .C1(new_n343), .C2(new_n348), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n342), .A2(new_n331), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n354), .B1(new_n289), .B2(new_n290), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT81), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n344), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n339), .A2(KEYINPUT81), .A3(new_n341), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT29), .B1(new_n286), .B2(new_n287), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n359), .B1(KEYINPUT3), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n355), .A2(new_n361), .A3(new_n326), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n323), .B1(new_n353), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n362), .ZN(new_n364));
  AOI211_X1 g163(.A(new_n322), .B(new_n364), .C1(new_n351), .C2(new_n352), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n321), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n347), .A2(new_n340), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n355), .B1(new_n367), .B2(new_n345), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT85), .B1(new_n368), .B2(new_n327), .ZN(new_n369));
  INV_X1    g168(.A(new_n352), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n362), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(new_n322), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n353), .A2(new_n323), .A3(new_n362), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n372), .A2(new_n320), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n366), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT73), .ZN(new_n376));
  INV_X1    g175(.A(G113gat), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n376), .B1(new_n377), .B2(G120gat), .ZN(new_n378));
  INV_X1    g177(.A(G120gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n379), .A2(KEYINPUT73), .A3(G113gat), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n378), .B(new_n380), .C1(G113gat), .C2(new_n379), .ZN(new_n381));
  XNOR2_X1  g180(.A(G127gat), .B(G134gat), .ZN(new_n382));
  XOR2_X1   g181(.A(KEYINPUT74), .B(KEYINPUT1), .Z(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n382), .ZN(new_n385));
  XNOR2_X1  g184(.A(G113gat), .B(G120gat), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n385), .B1(KEYINPUT1), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n273), .A2(new_n275), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n389), .B1(new_n390), .B2(new_n244), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n389), .B(new_n244), .C1(new_n296), .C2(new_n297), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G227gat), .A2(G233gat), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT33), .ZN(new_n396));
  OAI22_X1  g195(.A1(new_n394), .A2(new_n395), .B1(KEYINPUT32), .B2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G15gat), .B(G43gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(G71gat), .B(G99gat), .ZN(new_n399));
  XOR2_X1   g198(.A(new_n398), .B(new_n399), .Z(new_n400));
  NAND2_X1  g199(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n244), .B1(new_n296), .B2(new_n297), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n388), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n403), .A2(new_n395), .A3(new_n392), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT76), .B(KEYINPUT34), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n404), .B(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n395), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n408), .B1(new_n391), .B2(new_n393), .ZN(new_n409));
  INV_X1    g208(.A(new_n400), .ZN(new_n410));
  OR2_X1    g209(.A1(new_n410), .A2(KEYINPUT75), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(KEYINPUT75), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(KEYINPUT33), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n409), .A2(KEYINPUT32), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n401), .A2(new_n407), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n403), .A2(new_n392), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT32), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n416), .A2(new_n408), .B1(new_n417), .B2(KEYINPUT33), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n414), .B1(new_n418), .B2(new_n410), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n404), .B(new_n405), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n375), .A2(new_n415), .A3(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n318), .A2(new_n422), .ZN(new_n423));
  XOR2_X1   g222(.A(KEYINPUT91), .B(KEYINPUT35), .Z(new_n424));
  AND3_X1   g223(.A1(new_n339), .A2(KEYINPUT81), .A3(new_n341), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT81), .B1(new_n339), .B2(new_n341), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n388), .B(new_n342), .C1(new_n427), .C2(new_n340), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT5), .ZN(new_n429));
  NAND2_X1  g228(.A1(G225gat), .A2(G233gat), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n339), .A2(new_n384), .A3(new_n341), .A4(new_n387), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT4), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(KEYINPUT82), .B(KEYINPUT4), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT84), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n436), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT84), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(new_n439), .A3(new_n433), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n432), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT4), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(KEYINPUT83), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n432), .A2(new_n435), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT83), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n446), .B1(new_n432), .B2(KEYINPUT4), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n444), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n448), .A2(new_n428), .A3(new_n430), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n388), .B1(new_n425), .B2(new_n426), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n432), .ZN(new_n451));
  INV_X1    g250(.A(new_n430), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n429), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n431), .A2(new_n441), .B1(new_n449), .B2(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(G1gat), .B(G29gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n455), .B(G85gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(KEYINPUT0), .B(G57gat), .ZN(new_n457));
  XOR2_X1   g256(.A(new_n456), .B(new_n457), .Z(new_n458));
  AOI21_X1  g257(.A(KEYINPUT6), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n431), .A2(new_n441), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n449), .A2(new_n453), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  XOR2_X1   g261(.A(new_n458), .B(KEYINPUT87), .Z(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n458), .B1(new_n460), .B2(new_n461), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n459), .A2(new_n465), .B1(KEYINPUT6), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n423), .A2(new_n424), .A3(new_n468), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n375), .A2(new_n415), .A3(new_n421), .ZN(new_n470));
  INV_X1    g269(.A(new_n459), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n466), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n459), .B1(new_n458), .B2(new_n454), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n311), .A2(new_n316), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT92), .B1(new_n475), .B2(KEYINPUT35), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT92), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT35), .ZN(new_n478));
  AOI211_X1 g277(.A(new_n477), .B(new_n478), .C1(new_n470), .C2(new_n474), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n469), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n467), .A2(new_n310), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT37), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n293), .A2(new_n482), .A3(new_n295), .A4(new_n303), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n307), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n482), .B1(new_n314), .B2(new_n295), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT38), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n301), .A2(new_n292), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n294), .B1(new_n276), .B2(new_n204), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n487), .B(KEYINPUT37), .C1(new_n292), .C2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT38), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT89), .B1(new_n484), .B2(new_n491), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n489), .A2(new_n490), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT89), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n493), .A2(new_n494), .A3(new_n307), .A4(new_n483), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n481), .A2(new_n486), .A3(new_n492), .A4(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n439), .B1(new_n438), .B2(new_n433), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n434), .A2(KEYINPUT84), .A3(new_n436), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n428), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT39), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(new_n500), .A3(new_n452), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n389), .B1(new_n359), .B2(KEYINPUT3), .ZN(new_n502));
  AOI22_X1  g301(.A1(new_n437), .A2(new_n440), .B1(new_n502), .B2(new_n342), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n503), .A2(new_n430), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n450), .A2(new_n430), .A3(new_n432), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n500), .B1(new_n505), .B2(KEYINPUT88), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n506), .B1(KEYINPUT88), .B2(new_n505), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n501), .B(new_n463), .C1(new_n504), .C2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT40), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n465), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n464), .B1(new_n504), .B2(new_n500), .ZN(new_n511));
  OAI221_X1 g310(.A(new_n506), .B1(KEYINPUT88), .B2(new_n505), .C1(new_n503), .C2(new_n430), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT40), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n514), .A2(new_n311), .A3(new_n316), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n496), .A2(new_n375), .A3(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n516), .A2(KEYINPUT90), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT90), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n515), .A2(new_n375), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n518), .B1(new_n519), .B2(new_n496), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  AND3_X1   g320(.A1(new_n421), .A2(new_n415), .A3(KEYINPUT36), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT36), .B1(new_n421), .B2(new_n415), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n472), .A2(new_n473), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n375), .B1(new_n317), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT86), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n317), .A2(new_n525), .ZN(new_n528));
  INV_X1    g327(.A(new_n375), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT86), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT36), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n407), .B1(new_n401), .B2(new_n414), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n419), .A2(new_n420), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n421), .A2(new_n415), .A3(KEYINPUT36), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n530), .A2(new_n531), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n527), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n480), .B1(new_n521), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G15gat), .B(G22gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(KEYINPUT95), .ZN(new_n542));
  INV_X1    g341(.A(G1gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT16), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n545), .A2(G1gat), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n544), .B1(new_n546), .B2(new_n542), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n547), .A2(G8gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(G8gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT96), .ZN(new_n551));
  OR3_X1    g350(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n553));
  AOI22_X1  g352(.A1(new_n552), .A2(new_n553), .B1(G29gat), .B2(G36gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(G43gat), .B(G50gat), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n554), .B1(KEYINPUT15), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(KEYINPUT15), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n556), .B(new_n557), .Z(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT17), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n551), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT97), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n550), .A2(new_n558), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT98), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT97), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n551), .A2(new_n564), .A3(new_n559), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n561), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT18), .ZN(new_n567));
  NAND2_X1  g366(.A1(G229gat), .A2(G233gat), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  OR3_X1    g368(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n563), .B1(new_n550), .B2(new_n558), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n568), .B(KEYINPUT13), .Z(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n567), .B1(new_n566), .B2(new_n569), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n570), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT94), .ZN(new_n576));
  XNOR2_X1  g375(.A(G113gat), .B(G141gat), .ZN(new_n577));
  INV_X1    g376(.A(G197gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(KEYINPUT11), .B(G169gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT93), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT12), .ZN(new_n583));
  AND3_X1   g382(.A1(new_n575), .A2(new_n576), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n583), .B1(new_n575), .B2(new_n576), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G99gat), .A2(G106gat), .ZN(new_n588));
  INV_X1    g387(.A(G85gat), .ZN(new_n589));
  INV_X1    g388(.A(G92gat), .ZN(new_n590));
  AOI22_X1  g389(.A1(KEYINPUT8), .A2(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n592), .B1(new_n589), .B2(new_n590), .ZN(new_n593));
  NAND4_X1  g392(.A1(KEYINPUT100), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT101), .ZN(new_n596));
  XOR2_X1   g395(.A(G99gat), .B(G106gat), .Z(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT102), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT10), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G57gat), .B(G64gat), .ZN(new_n603));
  AOI21_X1  g402(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n604));
  OR2_X1    g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G71gat), .B(G78gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n598), .B(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(KEYINPUT103), .B(KEYINPUT10), .Z(new_n609));
  AOI22_X1  g408(.A1(new_n602), .A2(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AND2_X1   g409(.A1(G230gat), .A2(G233gat), .ZN(new_n611));
  MUX2_X1   g410(.A(new_n610), .B(new_n608), .S(new_n611), .Z(new_n612));
  XNOR2_X1  g411(.A(G176gat), .B(G204gat), .ZN(new_n613));
  INV_X1    g412(.A(G148gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(KEYINPUT104), .B(G120gat), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n615), .B(new_n616), .Z(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n612), .B(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT105), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n587), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n540), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n607), .A2(KEYINPUT21), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n548), .A2(new_n624), .A3(new_n549), .ZN(new_n625));
  INV_X1    g424(.A(G183gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n607), .A2(KEYINPUT21), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n627), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(G231gat), .A2(G233gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G127gat), .B(G155gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(G211gat), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n630), .A2(G231gat), .A3(G233gat), .A4(new_n631), .ZN(new_n638));
  AND3_X1   g437(.A1(new_n634), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n637), .B1(new_n634), .B2(new_n638), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  OR3_X1    g441(.A1(new_n639), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n642), .B1(new_n639), .B2(new_n640), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(G232gat), .A2(G233gat), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT41), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n648), .B(KEYINPUT99), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(G162gat), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n600), .A2(new_n559), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n598), .B(KEYINPUT102), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n558), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n651), .B(new_n653), .C1(new_n647), .C2(new_n646), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G134gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(G190gat), .B(G218gat), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n650), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n657), .A2(new_n650), .A3(new_n658), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n623), .A2(new_n645), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n525), .B(KEYINPUT106), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g465(.A1(new_n663), .A2(new_n318), .ZN(new_n667));
  NAND2_X1  g466(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n668));
  INV_X1    g467(.A(G8gat), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n545), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n667), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT42), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n673), .B(new_n674), .C1(new_n669), .C2(new_n667), .ZN(G1325gat));
  NOR2_X1   g474(.A1(new_n533), .A2(new_n534), .ZN(new_n676));
  AOI21_X1  g475(.A(G15gat), .B1(new_n663), .B2(new_n676), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n524), .A2(G15gat), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n677), .B1(new_n663), .B2(new_n678), .ZN(G1326gat));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n529), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(G22gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  NAND2_X1  g482(.A1(new_n622), .A2(new_n645), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT108), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n527), .A2(new_n538), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n516), .A2(KEYINPUT90), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n519), .A2(new_n518), .A3(new_n496), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(KEYINPUT35), .B1(new_n528), .B2(new_n422), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n477), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n475), .A2(KEYINPUT92), .A3(KEYINPUT35), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI22_X1  g493(.A1(new_n687), .A2(new_n690), .B1(new_n694), .B2(new_n469), .ZN(new_n695));
  INV_X1    g494(.A(new_n662), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT44), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n524), .A2(new_n526), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n698), .B1(new_n517), .B2(new_n520), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n696), .B1(new_n699), .B2(new_n480), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n686), .B1(new_n697), .B2(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n701), .B1(new_n540), .B2(new_n662), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n704), .A2(KEYINPUT108), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n664), .B(new_n685), .C1(new_n703), .C2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT109), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI211_X1 g507(.A(KEYINPUT44), .B(new_n696), .C1(new_n699), .C2(new_n480), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT108), .B1(new_n704), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n697), .A2(new_n686), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n712), .A2(KEYINPUT109), .A3(new_n664), .A4(new_n685), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n708), .A2(G29gat), .A3(new_n713), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n684), .A2(new_n695), .A3(new_n696), .ZN(new_n715));
  INV_X1    g514(.A(G29gat), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n715), .A2(new_n716), .A3(new_n664), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT45), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT110), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n714), .A2(KEYINPUT110), .A3(new_n718), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(G1328gat));
  INV_X1    g522(.A(G36gat), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n715), .A2(new_n724), .A3(new_n318), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n725), .B1(KEYINPUT111), .B2(KEYINPUT46), .ZN(new_n726));
  NAND2_X1  g525(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n727));
  XOR2_X1   g526(.A(new_n726), .B(new_n727), .Z(new_n728));
  AOI21_X1  g527(.A(new_n684), .B1(new_n710), .B2(new_n711), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n729), .A2(new_n318), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n728), .B1(new_n724), .B2(new_n730), .ZN(G1329gat));
  AOI21_X1  g530(.A(G43gat), .B1(new_n715), .B2(new_n676), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n524), .A2(G43gat), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n732), .B1(new_n729), .B2(new_n733), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n734), .B(KEYINPUT47), .Z(G1330gat));
  NAND3_X1  g534(.A1(new_n729), .A2(G50gat), .A3(new_n529), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n715), .A2(new_n529), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n736), .B1(G50gat), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g538(.A1(new_n699), .A2(new_n480), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n586), .A2(new_n645), .A3(new_n662), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n740), .A2(new_n621), .A3(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n664), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XOR2_X1   g543(.A(new_n744), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g544(.A1(new_n742), .A2(new_n317), .ZN(new_n746));
  NOR2_X1   g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  AND2_X1   g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n749), .B1(new_n746), .B2(new_n747), .ZN(G1333gat));
  INV_X1    g549(.A(new_n676), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n742), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n524), .A2(G71gat), .ZN(new_n753));
  OAI22_X1  g552(.A1(new_n752), .A2(G71gat), .B1(new_n742), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g554(.A1(new_n742), .A2(new_n375), .ZN(new_n756));
  XOR2_X1   g555(.A(KEYINPUT112), .B(G78gat), .Z(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1335gat));
  INV_X1    g557(.A(new_n645), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(new_n586), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n712), .A2(new_n621), .A3(new_n760), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n761), .A2(new_n589), .A3(new_n743), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n700), .A2(new_n760), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT51), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n700), .A2(KEYINPUT51), .A3(new_n760), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n621), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(G85gat), .B1(new_n769), .B2(new_n664), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n762), .A2(new_n770), .ZN(G1336gat));
  AND3_X1   g570(.A1(new_n712), .A2(new_n621), .A3(new_n760), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n590), .B1(new_n772), .B2(new_n318), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n318), .A2(new_n590), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n768), .B2(new_n775), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT113), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n765), .A2(new_n778), .A3(new_n766), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n763), .A2(KEYINPUT113), .A3(new_n764), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n621), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n781), .A2(new_n782), .A3(new_n775), .ZN(new_n783));
  OAI21_X1  g582(.A(KEYINPUT52), .B1(new_n773), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n777), .A2(new_n784), .ZN(G1337gat));
  NAND3_X1  g584(.A1(new_n772), .A2(KEYINPUT114), .A3(new_n524), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n787), .B1(new_n761), .B2(new_n537), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n786), .A2(G99gat), .A3(new_n788), .ZN(new_n789));
  OR2_X1    g588(.A1(new_n751), .A2(G99gat), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n789), .B1(new_n768), .B2(new_n790), .ZN(G1338gat));
  INV_X1    g590(.A(G106gat), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n792), .B1(new_n772), .B2(new_n529), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n782), .A2(G106gat), .A3(new_n375), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n767), .A2(new_n794), .ZN(new_n795));
  OR2_X1    g594(.A1(new_n795), .A2(KEYINPUT53), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n779), .A2(new_n780), .A3(new_n794), .ZN(new_n798));
  OAI21_X1  g597(.A(KEYINPUT53), .B1(new_n793), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(G1339gat));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(new_n610), .B2(new_n611), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n802), .B1(new_n611), .B2(new_n610), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n610), .A2(new_n611), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n801), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT115), .B1(new_n805), .B2(new_n618), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT115), .ZN(new_n807));
  AOI211_X1 g606(.A(new_n807), .B(new_n617), .C1(new_n804), .C2(new_n801), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n803), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n612), .A2(new_n617), .ZN(new_n812));
  OAI211_X1 g611(.A(KEYINPUT55), .B(new_n803), .C1(new_n806), .C2(new_n808), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n586), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n570), .A2(new_n574), .A3(new_n573), .A4(new_n583), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n566), .A2(new_n569), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n817), .B1(new_n571), .B2(new_n572), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n581), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n621), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n662), .B1(new_n815), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n820), .B1(new_n660), .B2(new_n661), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n814), .A2(new_n824), .A3(KEYINPUT116), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n657), .A2(new_n650), .A3(new_n658), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n816), .B(new_n819), .C1(new_n827), .C2(new_n659), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n826), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n825), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n645), .B1(new_n823), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n741), .A2(new_n782), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n835), .A2(new_n664), .A3(new_n423), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(new_n587), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(new_n377), .ZN(G1340gat));
  NOR2_X1   g637(.A1(new_n836), .A2(new_n782), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(new_n379), .ZN(G1341gat));
  INV_X1    g639(.A(new_n836), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n759), .ZN(new_n842));
  INV_X1    g641(.A(G127gat), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT117), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n842), .B(new_n844), .ZN(G1342gat));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n836), .A2(new_n696), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n846), .B1(new_n848), .B2(G134gat), .ZN(new_n849));
  INV_X1    g648(.A(G134gat), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n847), .A2(KEYINPUT118), .A3(new_n850), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n847), .A2(KEYINPUT56), .A3(new_n850), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT56), .B1(new_n847), .B2(new_n850), .ZN(new_n853));
  OAI22_X1  g652(.A1(new_n849), .A2(new_n851), .B1(new_n852), .B2(new_n853), .ZN(G1343gat));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT58), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n858));
  INV_X1    g657(.A(G141gat), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n524), .A2(new_n375), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(KEYINPUT119), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n835), .A2(new_n664), .A3(new_n317), .A4(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n859), .B1(new_n862), .B2(new_n587), .ZN(new_n863));
  AOI22_X1  g662(.A1(new_n814), .A2(new_n586), .B1(new_n621), .B2(new_n821), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n830), .B(new_n825), .C1(new_n864), .C2(new_n662), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n833), .B1(new_n865), .B2(new_n645), .ZN(new_n866));
  OAI21_X1  g665(.A(KEYINPUT57), .B1(new_n866), .B2(new_n375), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n835), .A2(new_n868), .A3(new_n529), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n664), .A2(new_n537), .A3(new_n317), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n587), .A2(new_n859), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n867), .A2(new_n869), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  AOI211_X1 g672(.A(new_n857), .B(new_n858), .C1(new_n863), .C2(new_n873), .ZN(new_n874));
  AND4_X1   g673(.A1(new_n855), .A2(new_n863), .A3(new_n873), .A4(new_n856), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n874), .A2(new_n875), .ZN(G1344gat));
  INV_X1    g675(.A(new_n862), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(new_n614), .A3(new_n621), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n867), .A2(new_n869), .A3(new_n871), .ZN(new_n879));
  AOI211_X1 g678(.A(KEYINPUT59), .B(new_n614), .C1(new_n879), .C2(new_n621), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n815), .A2(new_n822), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n696), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n814), .A2(new_n824), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n759), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n868), .B(new_n529), .C1(new_n885), .C2(new_n833), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n867), .A2(new_n886), .A3(new_n621), .A4(new_n871), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n881), .B1(new_n887), .B2(G148gat), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n878), .B1(new_n880), .B2(new_n888), .ZN(G1345gat));
  AOI21_X1  g688(.A(G155gat), .B1(new_n877), .B2(new_n759), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n645), .A2(new_n333), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n890), .B1(new_n879), .B2(new_n891), .ZN(G1346gat));
  NAND4_X1  g691(.A1(new_n867), .A2(new_n869), .A3(new_n662), .A4(new_n871), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n893), .A2(KEYINPUT121), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(KEYINPUT121), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n894), .A2(G162gat), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n877), .A2(new_n334), .A3(new_n662), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(G1347gat));
  NOR2_X1   g697(.A1(new_n664), .A2(new_n317), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n835), .A2(new_n470), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n900), .A2(new_n587), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(new_n205), .ZN(G1348gat));
  NOR2_X1   g701(.A1(new_n900), .A2(new_n782), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n221), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n904), .B1(new_n206), .B2(new_n903), .ZN(G1349gat));
  INV_X1    g704(.A(new_n899), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n866), .A2(new_n422), .A3(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(new_n257), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n907), .A2(new_n759), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n239), .B1(new_n900), .B2(new_n645), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT60), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(KEYINPUT122), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n909), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n911), .A2(KEYINPUT122), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n913), .B(new_n914), .ZN(G1350gat));
  OR2_X1    g714(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n916), .B1(new_n900), .B2(new_n696), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(KEYINPUT123), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n919), .B(new_n916), .C1(new_n900), .C2(new_n696), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n918), .A2(KEYINPUT61), .A3(G190gat), .A4(new_n920), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(G1351gat));
  NOR2_X1   g724(.A1(new_n906), .A2(new_n524), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n867), .A2(new_n886), .A3(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(G197gat), .B1(new_n927), .B2(new_n587), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n866), .A2(new_n375), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n929), .A2(new_n926), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n930), .A2(new_n578), .A3(new_n586), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n928), .A2(new_n931), .ZN(G1352gat));
  INV_X1    g731(.A(KEYINPUT125), .ZN(new_n933));
  INV_X1    g732(.A(G204gat), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n929), .A2(new_n934), .A3(new_n621), .A4(new_n926), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n933), .B1(new_n935), .B2(KEYINPUT62), .ZN(new_n936));
  AND4_X1   g735(.A1(new_n934), .A2(new_n835), .A3(new_n529), .A4(new_n926), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT62), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n937), .A2(KEYINPUT125), .A3(new_n938), .A4(new_n621), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n867), .A2(new_n886), .A3(new_n621), .A4(new_n926), .ZN(new_n940));
  AOI22_X1  g739(.A1(new_n936), .A2(new_n939), .B1(G204gat), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT124), .B1(new_n935), .B2(KEYINPUT62), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n935), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(G1353gat));
  NAND4_X1  g743(.A1(new_n867), .A2(new_n886), .A3(new_n759), .A4(new_n926), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT63), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(KEYINPUT126), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n945), .A2(G211gat), .A3(new_n947), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n946), .A2(KEYINPUT126), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n930), .A2(new_n759), .A3(new_n279), .ZN(new_n951));
  INV_X1    g750(.A(new_n949), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n945), .A2(G211gat), .A3(new_n947), .A4(new_n952), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n950), .A2(new_n951), .A3(new_n953), .ZN(G1354gat));
  NAND3_X1  g753(.A1(new_n930), .A2(new_n280), .A3(new_n662), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n867), .A2(new_n886), .A3(new_n662), .A4(new_n926), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(G218gat), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT127), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n955), .A2(new_n957), .A3(KEYINPUT127), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1355gat));
endmodule


