//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 1 1 1 1 0 1 0 1 0 0 0 0 1 1 0 1 1 1 0 1 0 0 0 1 0 0 1 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 0 0 0 0 1 1 1 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT64), .Z(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n211));
  AND2_X1   g0011(.A1(new_n211), .A2(KEYINPUT67), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(KEYINPUT67), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n210), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  OR2_X1    g0014(.A1(new_n214), .A2(KEYINPUT68), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G116), .A2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n217));
  AND2_X1   g0017(.A1(KEYINPUT66), .A2(G68), .ZN(new_n218));
  NOR2_X1   g0018(.A1(KEYINPUT66), .A2(G68), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n216), .B(new_n217), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(new_n214), .B2(KEYINPUT68), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n209), .B1(new_n215), .B2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT69), .ZN(new_n227));
  INV_X1    g0027(.A(G13), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n209), .A2(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT0), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n234), .A2(G20), .ZN(new_n235));
  INV_X1    g0035(.A(G58), .ZN(new_n236));
  INV_X1    g0036(.A(G68), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g0038(.A(KEYINPUT65), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g0040(.A1(new_n236), .A2(new_n237), .A3(KEYINPUT65), .ZN(new_n241));
  NAND3_X1  g0041(.A1(new_n240), .A2(G50), .A3(new_n241), .ZN(new_n242));
  OAI221_X1 g0042(.A(new_n232), .B1(new_n235), .B2(new_n242), .C1(new_n224), .C2(new_n225), .ZN(new_n243));
  NOR2_X1   g0043(.A1(new_n227), .A2(new_n243), .ZN(G361));
  XNOR2_X1  g0044(.A(G238), .B(G244), .ZN(new_n245));
  INV_X1    g0045(.A(G232), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(KEYINPUT2), .B(G226), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G264), .B(G270), .Z(new_n250));
  XNOR2_X1  g0050(.A(G250), .B(G257), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G358));
  XOR2_X1   g0053(.A(G68), .B(G77), .Z(new_n254));
  XNOR2_X1  g0054(.A(G50), .B(G58), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XOR2_X1   g0056(.A(G107), .B(G116), .Z(new_n257));
  XNOR2_X1  g0057(.A(G87), .B(G97), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n256), .B(new_n259), .ZN(G351));
  NAND3_X1  g0060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n233), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT71), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT71), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n261), .A2(new_n264), .A3(new_n233), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n228), .A2(G1), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G20), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n207), .A2(G20), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(G50), .A3(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT8), .B(G58), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n208), .A2(G33), .ZN(new_n274));
  INV_X1    g0074(.A(G150), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  OAI22_X1  g0077(.A1(new_n273), .A2(new_n274), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G50), .A2(G58), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n208), .B1(new_n279), .B2(new_n237), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n266), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n272), .B(new_n281), .C1(G50), .C2(new_n268), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT9), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n233), .B1(G33), .B2(G41), .ZN(new_n284));
  INV_X1    g0084(.A(G41), .ZN(new_n285));
  INV_X1    g0085(.A(G45), .ZN(new_n286));
  AOI21_X1  g0086(.A(G1), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G226), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(KEYINPUT70), .ZN(new_n290));
  INV_X1    g0090(.A(G33), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n234), .B1(new_n291), .B2(new_n285), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT70), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G41), .A2(G45), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n293), .B1(new_n294), .B2(G1), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n290), .A2(new_n292), .A3(new_n295), .A4(G274), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n289), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT3), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n291), .ZN(new_n299));
  NAND2_X1  g0099(.A1(KEYINPUT3), .A2(G33), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G1698), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n301), .A2(G222), .A3(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n301), .A2(G223), .A3(G1698), .ZN(new_n304));
  INV_X1    g0104(.A(G77), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n303), .B(new_n304), .C1(new_n305), .C2(new_n301), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n297), .B1(new_n306), .B2(new_n284), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n282), .A2(new_n283), .B1(new_n307), .B2(G190), .ZN(new_n308));
  INV_X1    g0108(.A(G200), .ZN(new_n309));
  OAI221_X1 g0109(.A(new_n308), .B1(new_n283), .B2(new_n282), .C1(new_n309), .C2(new_n307), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT10), .ZN(new_n311));
  INV_X1    g0111(.A(G179), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n313), .B(new_n282), .C1(G169), .C2(new_n307), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G50), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n277), .A2(new_n316), .B1(new_n274), .B2(new_n305), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n317), .B1(G20), .B2(new_n220), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n318), .B1(new_n263), .B2(new_n265), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n319), .A2(KEYINPUT11), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n269), .A2(new_n262), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n321), .A2(G68), .A3(new_n271), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n319), .A2(KEYINPUT11), .ZN(new_n323));
  INV_X1    g0123(.A(new_n220), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT12), .B1(new_n324), .B2(new_n268), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT73), .ZN(new_n326));
  OR2_X1    g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OR3_X1    g0127(.A1(new_n268), .A2(KEYINPUT12), .A3(G68), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n325), .A2(new_n326), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n320), .A2(new_n322), .A3(new_n323), .A4(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT14), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT13), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n246), .A2(G1698), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n301), .B(new_n334), .C1(G226), .C2(G1698), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G33), .A2(G97), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n292), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT72), .ZN(new_n338));
  OR2_X1    g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n337), .A2(new_n338), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n288), .A2(G238), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n296), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n333), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  AOI211_X1 g0145(.A(KEYINPUT13), .B(new_n343), .C1(new_n339), .C2(new_n340), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n332), .B(G169), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n340), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n337), .A2(new_n338), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n344), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT13), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n341), .A2(new_n333), .A3(new_n344), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(G179), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n347), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n351), .A2(new_n352), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n332), .B1(new_n355), .B2(G169), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n331), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(G200), .B1(new_n345), .B2(new_n346), .ZN(new_n358));
  INV_X1    g0158(.A(new_n331), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n351), .A2(G190), .A3(new_n352), .ZN(new_n360));
  AND3_X1   g0160(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n288), .A2(G232), .ZN(new_n364));
  NOR2_X1   g0164(.A1(G223), .A2(G1698), .ZN(new_n365));
  INV_X1    g0165(.A(G226), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n365), .B1(new_n366), .B2(G1698), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n367), .A2(new_n301), .B1(G33), .B2(G87), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n364), .B(new_n296), .C1(new_n368), .C2(new_n292), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n369), .A2(new_n312), .ZN(new_n370));
  INV_X1    g0170(.A(G169), .ZN(new_n371));
  NOR3_X1   g0171(.A1(new_n284), .A2(new_n287), .A3(new_n246), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n366), .A2(G1698), .ZN(new_n373));
  AND2_X1   g0173(.A1(KEYINPUT3), .A2(G33), .ZN(new_n374));
  NOR2_X1   g0174(.A1(KEYINPUT3), .A2(G33), .ZN(new_n375));
  OAI221_X1 g0175(.A(new_n373), .B1(G223), .B2(G1698), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G33), .A2(G87), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n372), .B1(new_n378), .B2(new_n284), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n371), .B1(new_n379), .B2(new_n296), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n370), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(G58), .B1(new_n218), .B2(new_n219), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT74), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI211_X1 g0184(.A(KEYINPUT74), .B(G58), .C1(new_n218), .C2(new_n219), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(new_n238), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(G20), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n276), .A2(G159), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n299), .A2(new_n208), .A3(new_n300), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT7), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n299), .A2(KEYINPUT7), .A3(new_n208), .A4(new_n300), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n324), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n387), .A2(new_n388), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT16), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n262), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n386), .A2(G20), .B1(G159), .B2(new_n276), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n396), .B1(new_n393), .B2(G68), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n273), .B1(new_n207), .B2(G20), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n270), .A2(new_n403), .B1(new_n269), .B2(new_n273), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n381), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT18), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n369), .A2(new_n309), .ZN(new_n408));
  INV_X1    g0208(.A(G190), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n379), .A2(new_n409), .A3(new_n296), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n402), .A2(new_n404), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT17), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n404), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n415), .B1(new_n397), .B2(new_n401), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT18), .B1(new_n416), .B2(new_n381), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n416), .A2(KEYINPUT17), .A3(new_n411), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n407), .A2(new_n414), .A3(new_n417), .A4(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(G232), .A2(G1698), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n302), .A2(G238), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n301), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n422), .B(new_n284), .C1(G107), .C2(new_n301), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n288), .A2(G244), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(new_n296), .A3(new_n424), .ZN(new_n425));
  OR2_X1    g0225(.A1(new_n425), .A2(G179), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n305), .B1(new_n207), .B2(G20), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n321), .A2(new_n427), .B1(new_n305), .B2(new_n269), .ZN(new_n428));
  XNOR2_X1  g0228(.A(KEYINPUT15), .B(G87), .ZN(new_n429));
  OAI22_X1  g0229(.A1(new_n429), .A2(new_n274), .B1(new_n208), .B2(new_n305), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n273), .A2(new_n277), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n262), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n425), .A2(new_n371), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n426), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n433), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n425), .A2(G200), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n436), .B(new_n437), .C1(new_n409), .C2(new_n425), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  NOR4_X1   g0239(.A1(new_n315), .A2(new_n363), .A3(new_n419), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n269), .A2(new_n203), .ZN(new_n441));
  XNOR2_X1  g0241(.A(new_n441), .B(KEYINPUT25), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n207), .A2(G33), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n263), .A2(new_n265), .A3(new_n268), .A4(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n444), .A2(new_n203), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n301), .A2(new_n208), .A3(G87), .ZN(new_n448));
  XNOR2_X1  g0248(.A(new_n448), .B(KEYINPUT22), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT23), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(new_n208), .B2(G107), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n203), .A2(KEYINPUT23), .A3(G20), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G33), .A2(G116), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n451), .A2(new_n452), .B1(new_n454), .B2(new_n208), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n449), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT24), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT24), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n449), .A2(new_n458), .A3(new_n455), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n447), .B1(new_n460), .B2(new_n262), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n286), .A2(G1), .ZN(new_n462));
  XNOR2_X1  g0262(.A(KEYINPUT5), .B(G41), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n284), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G264), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n462), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G274), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n284), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n301), .A2(G257), .A3(G1698), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n301), .A2(G250), .A3(new_n302), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G294), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n475), .A2(KEYINPUT80), .A3(new_n284), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT80), .B1(new_n475), .B2(new_n284), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n471), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G169), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n465), .A2(KEYINPUT82), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n475), .A2(new_n284), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT82), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n464), .A2(new_n482), .A3(G264), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n480), .A2(new_n481), .A3(new_n470), .A4(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n479), .A2(KEYINPUT81), .B1(G179), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT81), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n478), .A2(new_n487), .A3(G169), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n461), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  OAI22_X1  g0289(.A1(new_n485), .A2(G200), .B1(new_n478), .B2(G190), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n461), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n301), .A2(G250), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n302), .B1(new_n493), .B2(KEYINPUT4), .ZN(new_n494));
  AND2_X1   g0294(.A1(KEYINPUT4), .A2(G244), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n302), .B(new_n495), .C1(new_n374), .C2(new_n375), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G283), .ZN(new_n497));
  INV_X1    g0297(.A(G244), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n498), .B1(new_n299), .B2(new_n300), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n496), .B(new_n497), .C1(new_n499), .C2(KEYINPUT4), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n284), .B1(new_n494), .B2(new_n500), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n464), .A2(G257), .B1(new_n467), .B2(new_n469), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(new_n309), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n276), .A2(G77), .ZN(new_n505));
  OR2_X1    g0305(.A1(new_n505), .A2(KEYINPUT75), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(KEYINPUT75), .ZN(new_n507));
  XNOR2_X1  g0307(.A(KEYINPUT76), .B(G97), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT6), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n509), .A2(G107), .ZN(new_n510));
  XNOR2_X1  g0310(.A(G97), .B(G107), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n508), .A2(new_n510), .B1(new_n511), .B2(new_n509), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n506), .B(new_n507), .C1(new_n512), .C2(new_n208), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n203), .B1(new_n391), .B2(new_n392), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n262), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OR2_X1    g0315(.A1(new_n444), .A2(new_n202), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n268), .A2(G97), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n515), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n501), .A2(new_n502), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n520), .A2(new_n409), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n504), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n503), .A2(G179), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n371), .B1(new_n501), .B2(new_n502), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n393), .A2(G107), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n508), .A2(new_n510), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n511), .A2(new_n509), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G20), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n526), .A2(new_n530), .A3(new_n506), .A4(new_n507), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n517), .B1(new_n531), .B2(new_n262), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n523), .A2(new_n525), .B1(new_n532), .B2(new_n516), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n522), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT77), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(KEYINPUT77), .B1(new_n522), .B2(new_n533), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n464), .A2(G270), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n470), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n301), .A2(G264), .A3(G1698), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n301), .A2(G257), .A3(new_n302), .ZN(new_n542));
  INV_X1    g0342(.A(G303), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n541), .B(new_n542), .C1(new_n543), .C2(new_n301), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n284), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT79), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n544), .A2(KEYINPUT79), .A3(new_n284), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n540), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G190), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n497), .A2(new_n208), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n551), .B1(new_n508), .B2(new_n291), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT20), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n262), .B1(new_n208), .B2(G116), .ZN(new_n554));
  OR3_X1    g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n553), .B1(new_n552), .B2(new_n554), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(G116), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n558), .B1(new_n207), .B2(G33), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n208), .A2(G116), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n321), .A2(new_n559), .B1(new_n267), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n550), .B(new_n563), .C1(new_n309), .C2(new_n549), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n549), .A2(G179), .A3(new_n562), .ZN(new_n566));
  INV_X1    g0366(.A(new_n540), .ZN(new_n567));
  INV_X1    g0367(.A(new_n548), .ZN(new_n568));
  AOI21_X1  g0368(.A(KEYINPUT79), .B1(new_n544), .B2(new_n284), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n371), .B1(new_n557), .B2(new_n561), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT21), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n572), .B1(new_n570), .B2(new_n571), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n566), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT19), .ZN(new_n576));
  XOR2_X1   g0376(.A(KEYINPUT76), .B(G97), .Z(new_n577));
  OAI21_X1  g0377(.A(new_n576), .B1(new_n577), .B2(new_n274), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n208), .B1(new_n336), .B2(new_n576), .ZN(new_n579));
  INV_X1    g0379(.A(G87), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n203), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n579), .B1(new_n508), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n301), .A2(new_n208), .A3(G68), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n578), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n584), .A2(new_n262), .B1(new_n269), .B2(new_n429), .ZN(new_n585));
  OR2_X1    g0385(.A1(new_n444), .A2(new_n580), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n301), .A2(G244), .A3(G1698), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n301), .A2(G238), .A3(new_n302), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n588), .A2(new_n589), .A3(new_n453), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n284), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n462), .A2(new_n468), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n292), .B(new_n592), .C1(G250), .C2(new_n462), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(G190), .A3(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT78), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n591), .A2(KEYINPUT78), .A3(G190), .A4(new_n593), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n591), .A2(new_n593), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(G200), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n587), .A2(new_n596), .A3(new_n597), .A4(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(new_n371), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n584), .A2(new_n262), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n269), .A2(new_n429), .ZN(new_n603));
  OR2_X1    g0403(.A1(new_n444), .A2(new_n429), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n591), .A2(new_n312), .A3(new_n593), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n601), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n600), .A2(new_n607), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n565), .A2(new_n575), .A3(new_n608), .ZN(new_n609));
  AND4_X1   g0409(.A1(new_n440), .A2(new_n492), .A3(new_n538), .A4(new_n609), .ZN(new_n610));
  XNOR2_X1  g0410(.A(new_n610), .B(KEYINPUT83), .ZN(G372));
  AND2_X1   g0411(.A1(new_n414), .A2(new_n418), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n362), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n613), .B1(new_n357), .B2(new_n435), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n416), .A2(KEYINPUT18), .A3(new_n381), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n400), .A2(new_n387), .A3(new_n388), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n262), .ZN(new_n617));
  AOI21_X1  g0417(.A(KEYINPUT16), .B1(new_n399), .B2(new_n394), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n404), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n381), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n406), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n615), .A2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n311), .B1(new_n614), .B2(new_n623), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n624), .A2(new_n314), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n520), .A2(new_n312), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n519), .B1(new_n626), .B2(new_n524), .ZN(new_n627));
  OAI21_X1  g0427(.A(KEYINPUT26), .B1(new_n608), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT26), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n599), .A2(new_n585), .A3(new_n594), .A4(new_n586), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n533), .A2(new_n629), .A3(new_n607), .A4(new_n630), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n628), .A2(new_n607), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n630), .A2(new_n607), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n633), .B1(new_n461), .B2(new_n490), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n534), .B(new_n634), .C1(new_n489), .C2(new_n575), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n440), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n625), .A2(new_n637), .ZN(G369));
  INV_X1    g0438(.A(new_n575), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n267), .A2(new_n208), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n640), .A2(KEYINPUT27), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(KEYINPUT27), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(G213), .A3(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(G343), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n639), .B(new_n564), .C1(new_n563), .C2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n575), .A2(new_n562), .A3(new_n645), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(G330), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n492), .B1(new_n461), .B2(new_n646), .ZN(new_n652));
  INV_X1    g0452(.A(new_n489), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n652), .B1(new_n653), .B2(new_n646), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n639), .A2(new_n645), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n492), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n489), .A2(new_n646), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n655), .A2(new_n660), .ZN(G399));
  NOR3_X1   g0461(.A1(new_n508), .A2(G116), .A3(new_n581), .ZN(new_n662));
  XOR2_X1   g0462(.A(new_n662), .B(KEYINPUT84), .Z(new_n663));
  NOR2_X1   g0463(.A1(new_n229), .A2(G41), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n663), .A2(new_n207), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n242), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n665), .B1(new_n666), .B2(new_n664), .ZN(new_n667));
  XOR2_X1   g0467(.A(new_n667), .B(KEYINPUT28), .Z(new_n668));
  AOI21_X1  g0468(.A(new_n645), .B1(new_n632), .B2(new_n635), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT29), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n533), .A2(new_n629), .A3(new_n600), .A4(new_n607), .ZN(new_n672));
  OAI21_X1  g0472(.A(KEYINPUT26), .B1(new_n633), .B2(new_n627), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(new_n673), .A3(new_n607), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(KEYINPUT86), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT86), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n672), .A2(new_n673), .A3(new_n676), .A4(new_n607), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n675), .A2(new_n635), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n670), .B1(new_n678), .B2(new_n646), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n671), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n609), .A2(new_n538), .A3(new_n492), .A4(new_n646), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(new_n598), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n549), .A2(new_n683), .A3(new_n626), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT30), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n549), .A2(new_n683), .A3(new_n626), .A4(KEYINPUT30), .ZN(new_n687));
  AOI21_X1  g0487(.A(G179), .B1(new_n591), .B2(new_n593), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n570), .A2(new_n688), .A3(new_n484), .A4(new_n520), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n686), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n690), .A2(new_n645), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n691), .A2(KEYINPUT31), .ZN(new_n692));
  XOR2_X1   g0492(.A(KEYINPUT85), .B(KEYINPUT31), .Z(new_n693));
  NAND2_X1  g0493(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n681), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G330), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n680), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n668), .B1(new_n698), .B2(G1), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT87), .ZN(G364));
  NOR2_X1   g0500(.A1(new_n228), .A2(G20), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n207), .B1(new_n701), .B2(G45), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n664), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n651), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(G330), .B2(new_n649), .ZN(new_n706));
  INV_X1    g0506(.A(new_n704), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n233), .B1(G20), .B2(new_n371), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n301), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n208), .A2(G179), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n712), .A2(G190), .A3(new_n309), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(G283), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n710), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n409), .A2(G179), .A3(G200), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(new_n208), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n716), .B1(G294), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n208), .A2(new_n312), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n409), .A2(new_n309), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n721), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n725), .A2(new_n309), .A3(G190), .ZN(new_n726));
  XNOR2_X1  g0526(.A(KEYINPUT33), .B(G317), .ZN(new_n727));
  AOI22_X1  g0527(.A1(new_n724), .A2(G326), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(G190), .A2(G200), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n711), .A2(new_n729), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n730), .A2(KEYINPUT90), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(KEYINPUT90), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT89), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n721), .A2(new_n735), .A3(new_n729), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n735), .B1(new_n721), .B2(new_n729), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI22_X1  g0538(.A1(new_n734), .A2(G329), .B1(G311), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n721), .A2(G190), .A3(new_n309), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n722), .A2(new_n711), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n741), .A2(G322), .B1(new_n743), .B2(G303), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n720), .A2(new_n728), .A3(new_n739), .A4(new_n744), .ZN(new_n745));
  OAI22_X1  g0545(.A1(new_n714), .A2(new_n203), .B1(new_n236), .B2(new_n740), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n723), .A2(new_n316), .B1(new_n742), .B2(new_n580), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n718), .A2(new_n202), .ZN(new_n749));
  AOI211_X1 g0549(.A(new_n710), .B(new_n749), .C1(G68), .C2(new_n726), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n738), .A2(G77), .ZN(new_n751));
  INV_X1    g0551(.A(G159), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n730), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT32), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n748), .A2(new_n750), .A3(new_n751), .A4(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n709), .B1(new_n745), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G13), .A2(G33), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n708), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n230), .A2(new_n710), .ZN(new_n761));
  XOR2_X1   g0561(.A(new_n761), .B(KEYINPUT88), .Z(new_n762));
  NAND2_X1  g0562(.A1(new_n666), .A2(new_n286), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n762), .B(new_n763), .C1(new_n286), .C2(new_n256), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n710), .A2(new_n229), .ZN(new_n765));
  AOI22_X1  g0565(.A1(G355), .A2(new_n765), .B1(new_n558), .B2(new_n229), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n707), .B(new_n756), .C1(new_n760), .C2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n759), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n768), .B1(new_n649), .B2(new_n769), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n706), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(G396));
  OR2_X1    g0572(.A1(new_n435), .A2(KEYINPUT93), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n435), .A2(KEYINPUT93), .ZN(new_n774));
  AND2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n775), .A2(new_n438), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n669), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n433), .A2(new_n645), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n773), .A2(new_n438), .A3(new_n778), .A4(new_n774), .ZN(new_n779));
  INV_X1    g0579(.A(new_n435), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(new_n645), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n777), .B1(new_n669), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n696), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n784), .B(KEYINPUT94), .Z(new_n785));
  AOI21_X1  g0585(.A(new_n704), .B1(new_n783), .B2(new_n696), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n734), .A2(G311), .B1(G116), .B2(new_n738), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n301), .B(new_n749), .C1(G87), .C2(new_n713), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n726), .A2(G283), .B1(new_n724), .B2(G303), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n741), .A2(G294), .B1(new_n743), .B2(G107), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n788), .A2(new_n789), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n714), .A2(new_n237), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n710), .B(new_n793), .C1(G50), .C2(new_n743), .ZN(new_n794));
  INV_X1    g0594(.A(G132), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n794), .B1(new_n236), .B2(new_n718), .C1(new_n795), .C2(new_n733), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT91), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n726), .A2(G150), .B1(new_n724), .B2(G137), .ZN(new_n799));
  INV_X1    g0599(.A(G143), .ZN(new_n800));
  INV_X1    g0600(.A(new_n738), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n799), .B1(new_n800), .B2(new_n740), .C1(new_n801), .C2(new_n752), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT34), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n798), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n796), .A2(new_n797), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n792), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n709), .B1(new_n806), .B2(KEYINPUT92), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(KEYINPUT92), .B2(new_n806), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n708), .A2(new_n757), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n707), .B1(new_n305), .B2(new_n809), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n808), .B(new_n810), .C1(new_n758), .C2(new_n782), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n787), .A2(new_n811), .ZN(G384));
  AOI211_X1 g0612(.A(new_n558), .B(new_n235), .C1(new_n529), .C2(KEYINPUT35), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(KEYINPUT35), .B2(new_n529), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT36), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n666), .A2(G77), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n384), .A2(new_n385), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n816), .A2(new_n817), .B1(G50), .B2(new_n237), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n818), .A2(G1), .A3(new_n228), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT95), .ZN(new_n821));
  INV_X1    g0621(.A(new_n782), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n331), .A2(new_n645), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n357), .A2(new_n362), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(G169), .B1(new_n345), .B2(new_n346), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(KEYINPUT14), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n826), .A2(new_n353), .A3(new_n347), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n331), .B(new_n645), .C1(new_n827), .C2(new_n361), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n822), .B1(new_n824), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n693), .B1(new_n690), .B2(new_n645), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(KEYINPUT31), .B2(new_n691), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n681), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT40), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n399), .A2(new_n400), .B1(new_n263), .B2(new_n265), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n393), .A2(G68), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n387), .A2(new_n388), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n396), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n415), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(new_n643), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(new_n612), .B2(new_n622), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n412), .B1(new_n381), .B2(new_n840), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT96), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n412), .B(KEYINPUT96), .C1(new_n381), .C2(new_n840), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n846), .A2(new_n847), .A3(new_n842), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(KEYINPUT37), .ZN(new_n849));
  OAI21_X1  g0649(.A(KEYINPUT97), .B1(new_n416), .B2(new_n643), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT97), .ZN(new_n851));
  INV_X1    g0651(.A(new_n643), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n619), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  AOI221_X4 g0654(.A(new_n415), .B1(new_n408), .B2(new_n410), .C1(new_n397), .C2(new_n401), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n855), .A2(new_n405), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT37), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n843), .B1(new_n849), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT38), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT100), .ZN(new_n861));
  INV_X1    g0661(.A(new_n854), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n419), .A2(new_n862), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n857), .B1(new_n854), .B2(new_n856), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n866), .A2(KEYINPUT98), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT98), .B1(new_n866), .B2(new_n867), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n860), .B(new_n861), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT98), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n854), .A2(new_n856), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT37), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n874), .A2(new_n858), .B1(new_n419), .B2(new_n862), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n872), .B1(new_n875), .B2(KEYINPUT38), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n866), .A2(KEYINPUT98), .A3(new_n867), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n861), .B1(new_n878), .B2(new_n860), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n835), .B1(new_n871), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n864), .B1(KEYINPUT37), .B2(new_n848), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n867), .B1(new_n881), .B2(new_n843), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n833), .B1(new_n860), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n880), .B1(KEYINPUT40), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n440), .A2(new_n832), .ZN(new_n885));
  OAI21_X1  g0685(.A(G330), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n886), .B1(new_n884), .B2(new_n885), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n860), .A2(new_n882), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n824), .A2(new_n828), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n775), .A2(new_n645), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n890), .B1(new_n669), .B2(new_n776), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n888), .A2(new_n889), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n622), .B2(new_n852), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT39), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n860), .B(new_n895), .C1(new_n868), .C2(new_n869), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT99), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n878), .A2(KEYINPUT99), .A3(new_n895), .A4(new_n860), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n888), .A2(KEYINPUT39), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n827), .A2(new_n331), .A3(new_n646), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n894), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n440), .B1(new_n671), .B2(new_n679), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n625), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n904), .B(new_n906), .ZN(new_n907));
  OAI22_X1  g0707(.A1(new_n887), .A2(new_n907), .B1(new_n207), .B2(new_n701), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n887), .A2(new_n907), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n821), .B1(new_n908), .B2(new_n909), .ZN(G367));
  NAND2_X1  g0710(.A1(new_n519), .A2(new_n645), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n534), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n533), .A2(new_n645), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT101), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n489), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n645), .B1(new_n917), .B2(new_n627), .ZN(new_n918));
  INV_X1    g0718(.A(new_n914), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n657), .A2(new_n919), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n920), .B(KEYINPUT42), .Z(new_n921));
  INV_X1    g0721(.A(KEYINPUT43), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n587), .A2(new_n646), .ZN(new_n923));
  MUX2_X1   g0723(.A(new_n633), .B(new_n607), .S(new_n923), .Z(new_n924));
  OAI22_X1  g0724(.A1(new_n918), .A2(new_n921), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n922), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n925), .B(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n655), .A2(new_n915), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n927), .B(new_n928), .Z(new_n929));
  XOR2_X1   g0729(.A(new_n664), .B(KEYINPUT41), .Z(new_n930));
  INV_X1    g0730(.A(KEYINPUT44), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n660), .B2(new_n914), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT103), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n932), .A2(new_n933), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n659), .A2(KEYINPUT44), .A3(new_n919), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT102), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n936), .A2(new_n937), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n934), .A2(new_n935), .A3(new_n938), .A4(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n659), .A2(new_n919), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT45), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n655), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n657), .B1(new_n654), .B2(new_n656), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(new_n650), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n946), .A2(new_n697), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n940), .A2(new_n655), .A3(new_n942), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n944), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n930), .B1(new_n949), .B2(new_n698), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n702), .B(KEYINPUT104), .Z(new_n951));
  OAI21_X1  g0751(.A(new_n929), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n714), .A2(new_n305), .B1(new_n800), .B2(new_n723), .ZN(new_n953));
  INV_X1    g0753(.A(new_n730), .ZN(new_n954));
  AOI211_X1 g0754(.A(new_n710), .B(new_n953), .C1(G137), .C2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n718), .A2(new_n237), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n738), .A2(G50), .ZN(new_n958));
  INV_X1    g0758(.A(new_n726), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n959), .A2(new_n752), .B1(new_n740), .B2(new_n275), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(G58), .B2(new_n743), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n955), .A2(new_n957), .A3(new_n958), .A4(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n710), .B1(new_n740), .B2(new_n543), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT46), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n743), .A2(G116), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n966), .B1(new_n964), .B2(new_n965), .C1(new_n203), .C2(new_n718), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n726), .A2(G294), .B1(new_n724), .B2(G311), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n713), .A2(new_n508), .B1(G317), .B2(new_n954), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n968), .B(new_n969), .C1(new_n801), .C2(new_n715), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n962), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT47), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n708), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n924), .A2(new_n759), .ZN(new_n974));
  INV_X1    g0774(.A(new_n762), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n760), .B1(new_n230), .B2(new_n429), .C1(new_n975), .C2(new_n252), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n973), .A2(new_n704), .A3(new_n974), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n952), .A2(new_n977), .ZN(G387));
  INV_X1    g0778(.A(new_n664), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n947), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n946), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n980), .B1(new_n698), .B2(new_n981), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n249), .A2(new_n286), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n983), .A2(new_n762), .B1(new_n663), .B2(new_n765), .ZN(new_n984));
  INV_X1    g0784(.A(new_n273), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n316), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT50), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n286), .B1(new_n237), .B2(new_n305), .ZN(new_n988));
  NOR3_X1   g0788(.A1(new_n663), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n984), .A2(new_n989), .B1(G107), .B2(new_n230), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n760), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n704), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n742), .A2(new_n305), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n994), .B1(new_n275), .B2(new_n730), .C1(new_n959), .C2(new_n273), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(G68), .B2(new_n738), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n718), .A2(new_n429), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n710), .B1(new_n741), .B2(G50), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n713), .A2(G97), .B1(new_n724), .B2(G159), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n996), .A2(new_n997), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n301), .B1(new_n954), .B2(G326), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n719), .A2(G283), .B1(new_n743), .B2(G294), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n724), .A2(G322), .ZN(new_n1003));
  INV_X1    g0803(.A(G317), .ZN(new_n1004));
  INV_X1    g0804(.A(G311), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1003), .B1(new_n740), .B2(new_n1004), .C1(new_n1005), .C2(new_n959), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(G303), .B2(new_n738), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT105), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1002), .B1(new_n1010), .B2(KEYINPUT48), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(KEYINPUT48), .B2(new_n1010), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT106), .Z(new_n1013));
  INV_X1    g0813(.A(KEYINPUT49), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1001), .B1(new_n558), .B2(new_n714), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  AND2_X1   g0815(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1000), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n992), .B1(new_n1017), .B2(new_n708), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n654), .B2(new_n769), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n951), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n982), .B(new_n1019), .C1(new_n946), .C2(new_n1020), .ZN(G393));
  NAND3_X1  g0821(.A1(new_n944), .A2(new_n948), .A3(new_n951), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n710), .B1(new_n714), .B2(new_n203), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n726), .A2(G303), .B1(G322), .B2(new_n954), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n715), .B2(new_n742), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1023), .B(new_n1025), .C1(G116), .C2(new_n719), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n740), .A2(new_n1005), .B1(new_n723), .B2(new_n1004), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT108), .Z(new_n1028));
  OR2_X1    g0828(.A1(new_n1028), .A2(KEYINPUT52), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(KEYINPUT52), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n738), .A2(G294), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1026), .A2(new_n1029), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n959), .A2(new_n316), .B1(new_n742), .B2(new_n220), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(G143), .B2(new_n954), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n740), .A2(new_n752), .B1(new_n723), .B2(new_n275), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT51), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n738), .A2(new_n985), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n718), .A2(new_n305), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n710), .B(new_n1038), .C1(G87), .C2(new_n713), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1034), .A2(new_n1036), .A3(new_n1037), .A4(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n709), .B1(new_n1032), .B2(new_n1040), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n760), .B1(new_n230), .B2(new_n577), .C1(new_n975), .C2(new_n259), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n704), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT107), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1041), .B(new_n1044), .C1(new_n915), .C2(new_n759), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1022), .A2(new_n1046), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n949), .A2(new_n664), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n948), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n1049), .A2(new_n943), .B1(new_n697), .B2(new_n946), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1047), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(G390));
  NAND3_X1  g0852(.A1(new_n678), .A2(new_n646), .A3(new_n776), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n890), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT109), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1053), .A2(KEYINPUT109), .A3(new_n1054), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1057), .A2(new_n889), .A3(new_n1058), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1059), .B(new_n902), .C1(new_n871), .C2(new_n879), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n889), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n902), .B1(new_n891), .B2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n898), .A2(new_n899), .A3(new_n900), .A4(new_n1062), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n695), .A2(G330), .A3(new_n782), .A4(new_n889), .ZN(new_n1064));
  AND3_X1   g0864(.A1(new_n1060), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(G330), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n681), .B2(new_n831), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n829), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1065), .A2(new_n1069), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n901), .A2(new_n758), .ZN(new_n1071));
  INV_X1    g0871(.A(G125), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n301), .B1(new_n714), .B2(new_n316), .C1(new_n733), .C2(new_n1072), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT110), .Z(new_n1074));
  OR3_X1    g0874(.A1(new_n742), .A2(KEYINPUT53), .A3(new_n275), .ZN(new_n1075));
  OAI21_X1  g0875(.A(KEYINPUT53), .B1(new_n742), .B2(new_n275), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1075), .B(new_n1076), .C1(new_n752), .C2(new_n718), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n726), .A2(G137), .B1(new_n741), .B2(G132), .ZN(new_n1078));
  INV_X1    g0878(.A(G128), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(KEYINPUT54), .B(G143), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1078), .B1(new_n1079), .B2(new_n723), .C1(new_n801), .C2(new_n1080), .ZN(new_n1081));
  OR3_X1    g0881(.A1(new_n1074), .A2(new_n1077), .A3(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n793), .B1(G116), .B2(new_n741), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n734), .A2(G294), .B1(new_n508), .B2(new_n738), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n726), .A2(G107), .B1(new_n724), .B2(G283), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n301), .B(new_n1038), .C1(G87), .C2(new_n743), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .A4(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n709), .B1(new_n1082), .B2(new_n1087), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n707), .B(new_n1088), .C1(new_n273), .C2(new_n809), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n1070), .A2(new_n951), .B1(new_n1071), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n440), .A2(new_n1067), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n625), .A2(new_n905), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1066), .B(new_n822), .C1(new_n681), .C2(new_n831), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1064), .B1(new_n1094), .B2(new_n889), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1061), .B1(new_n696), .B2(new_n822), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n891), .B1(new_n1097), .B2(new_n1068), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1093), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n1065), .B2(new_n1069), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1068), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1060), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1098), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1106), .B(new_n1064), .C1(new_n889), .C2(new_n1094), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1092), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1103), .A2(new_n1104), .A3(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1100), .A2(new_n1109), .A3(new_n664), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1090), .A2(new_n1110), .ZN(G378));
  AND2_X1   g0911(.A1(new_n829), .A2(new_n832), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(KEYINPUT40), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n860), .B1(new_n868), .B2(new_n869), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(KEYINPUT100), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1113), .B1(new_n1115), .B2(new_n870), .ZN(new_n1116));
  OAI21_X1  g0916(.A(G330), .B1(new_n883), .B2(KEYINPUT40), .ZN(new_n1117));
  OAI21_X1  g0917(.A(KEYINPUT114), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT114), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1112), .A2(new_n888), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1066), .B1(new_n1120), .B2(new_n834), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n880), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n282), .A2(new_n852), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT112), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n315), .B(new_n1124), .ZN(new_n1125));
  XOR2_X1   g0925(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1126));
  XOR2_X1   g0926(.A(new_n1125), .B(new_n1126), .Z(new_n1127));
  NAND3_X1  g0927(.A1(new_n1118), .A2(new_n1122), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1127), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1129), .A2(new_n1119), .A3(new_n880), .A4(new_n1121), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n904), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1128), .A2(new_n904), .A3(new_n1130), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1133), .A2(new_n951), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n809), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n704), .B1(G50), .B2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n714), .A2(new_n236), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G116), .B2(new_n724), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1139), .B1(new_n202), .B2(new_n959), .C1(new_n203), .C2(new_n740), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n957), .A2(new_n285), .A3(new_n710), .A4(new_n994), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n801), .A2(new_n429), .B1(new_n733), .B2(new_n715), .ZN(new_n1142));
  NOR3_X1   g0942(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(KEYINPUT58), .ZN(new_n1144));
  AOI21_X1  g0944(.A(G50), .B1(new_n291), .B2(new_n285), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n301), .B2(G41), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT111), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n723), .A2(new_n1072), .B1(new_n742), .B2(new_n1080), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n959), .A2(new_n795), .B1(new_n740), .B2(new_n1079), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1149), .B(new_n1150), .C1(G150), .C2(new_n719), .ZN(new_n1151));
  INV_X1    g0951(.A(G137), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1151), .B1(new_n1152), .B2(new_n801), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1153), .A2(KEYINPUT59), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(KEYINPUT59), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n713), .A2(G159), .ZN(new_n1156));
  AOI211_X1 g0956(.A(G33), .B(G41), .C1(new_n954), .C2(G124), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n1148), .B1(KEYINPUT58), .B2(new_n1143), .C1(new_n1154), .C2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1137), .B1(new_n1159), .B2(new_n708), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n1127), .B2(new_n758), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n1161), .B(KEYINPUT113), .Z(new_n1162));
  NAND2_X1  g0962(.A1(new_n1135), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT115), .ZN(new_n1165));
  NOR3_X1   g0965(.A1(new_n1065), .A2(new_n1069), .A3(new_n1099), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1165), .B1(new_n1166), .B2(new_n1092), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1109), .A2(KEYINPUT115), .A3(new_n1093), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n1128), .A2(new_n904), .A3(new_n1130), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n904), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT57), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1169), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n664), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1176));
  AOI21_X1  g0976(.A(KEYINPUT57), .B1(new_n1169), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1164), .B1(new_n1175), .B2(new_n1177), .ZN(G375));
  NOR2_X1   g0978(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n1092), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n930), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(new_n1181), .A3(new_n1099), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n707), .B1(new_n237), .B2(new_n809), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n710), .B(new_n1138), .C1(G50), .C2(new_n719), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n741), .A2(G137), .B1(new_n724), .B2(G132), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1080), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n726), .A2(new_n1186), .B1(G159), .B2(new_n743), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1184), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n801), .A2(new_n275), .B1(new_n733), .B2(new_n1079), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n726), .A2(G116), .B1(new_n741), .B2(G283), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(G294), .A2(new_n724), .B1(new_n743), .B2(G97), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n301), .B1(new_n713), .B2(G77), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .A4(new_n997), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n801), .A2(new_n203), .B1(new_n733), .B2(new_n543), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n1188), .A2(new_n1189), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1195), .A2(KEYINPUT116), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(KEYINPUT116), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n708), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1183), .B1(new_n1196), .B2(new_n1198), .C1(new_n889), .C2(new_n758), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n1179), .B2(new_n1020), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1182), .A2(new_n1201), .ZN(G381));
  XOR2_X1   g1002(.A(G375), .B(KEYINPUT118), .Z(new_n1203));
  NAND2_X1  g1003(.A1(G378), .A2(KEYINPUT117), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT117), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1090), .A2(new_n1110), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n952), .A2(new_n977), .A3(new_n1051), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NOR4_X1   g1010(.A1(G393), .A2(G396), .A3(G384), .A4(G381), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1203), .A2(new_n1208), .A3(new_n1210), .A4(new_n1211), .ZN(G407));
  NAND2_X1  g1012(.A1(new_n644), .A2(G213), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1203), .A2(new_n1208), .A3(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(G407), .A2(G213), .A3(new_n1215), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT119), .ZN(G409));
  NAND2_X1  g1017(.A1(new_n1180), .A2(KEYINPUT60), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT60), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1179), .A2(new_n1219), .A3(new_n1092), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1108), .A2(new_n979), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1223), .A2(G384), .A3(new_n1201), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(G384), .B1(new_n1223), .B2(new_n1201), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(G378), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1109), .A2(KEYINPUT115), .A3(new_n1093), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT115), .B1(new_n1109), .B2(new_n1093), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1176), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n1172), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n979), .B1(new_n1169), .B2(new_n1173), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1228), .B(new_n1163), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1135), .A2(new_n1161), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1170), .A2(new_n1171), .A3(new_n930), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1169), .A2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1235), .B1(new_n1237), .B2(KEYINPUT120), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT120), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1169), .A2(new_n1236), .A3(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1207), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1213), .B(new_n1227), .C1(new_n1234), .C2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT121), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT63), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1243), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(G393), .B(new_n771), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1051), .B1(new_n952), .B2(new_n977), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1248), .B1(new_n1210), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1249), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1248), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1251), .A2(new_n1209), .A3(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT61), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1250), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT122), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1223), .A2(new_n1201), .ZN(new_n1257));
  INV_X1    g1057(.A(G384), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(G2897), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1213), .A2(new_n1260), .ZN(new_n1261));
  AND3_X1   g1061(.A1(new_n1259), .A2(new_n1224), .A3(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1261), .B1(new_n1259), .B2(new_n1224), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1256), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n1225), .A2(new_n1226), .B1(new_n1260), .B2(new_n1213), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1259), .A2(new_n1224), .A3(new_n1261), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1265), .A2(new_n1266), .A3(KEYINPUT122), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1264), .A2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1213), .B1(new_n1234), .B2(new_n1241), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1255), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT123), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1133), .A2(new_n1181), .A3(new_n1134), .ZN(new_n1273));
  OAI21_X1  g1073(.A(KEYINPUT120), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1235), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1274), .A2(new_n1240), .A3(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1208), .ZN(new_n1277));
  OAI211_X1 g1077(.A(G378), .B(new_n1164), .C1(new_n1175), .C2(new_n1177), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1227), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1280), .A2(new_n1244), .ZN(new_n1281));
  AND4_X1   g1081(.A1(new_n1271), .A2(new_n1279), .A3(new_n1213), .A4(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1214), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1271), .B1(new_n1283), .B2(new_n1281), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1270), .B1(new_n1282), .B2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(KEYINPUT124), .B1(new_n1247), .B2(new_n1285), .ZN(new_n1286));
  AOI211_X1 g1086(.A(new_n1214), .B(new_n1280), .C1(new_n1277), .C2(new_n1278), .ZN(new_n1287));
  OAI21_X1  g1087(.A(KEYINPUT121), .B1(new_n1287), .B2(KEYINPUT63), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT124), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1281), .ZN(new_n1292));
  OAI21_X1  g1092(.A(KEYINPUT123), .B1(new_n1269), .B2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1283), .A2(new_n1271), .A3(new_n1281), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1290), .A2(new_n1291), .A3(new_n1295), .A4(new_n1270), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1286), .A2(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(KEYINPUT125), .B1(new_n1287), .B2(KEYINPUT62), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT126), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1287), .A2(new_n1299), .A3(KEYINPUT62), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT62), .ZN(new_n1301));
  OAI21_X1  g1101(.A(KEYINPUT126), .B1(new_n1242), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT125), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1242), .A2(new_n1303), .A3(new_n1301), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1298), .A2(new_n1300), .A3(new_n1302), .A4(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1306));
  AOI21_X1  g1106(.A(KEYINPUT61), .B1(new_n1269), .B2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1305), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1250), .A2(new_n1253), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1297), .A2(new_n1310), .ZN(G405));
  AOI21_X1  g1111(.A(new_n1234), .B1(G375), .B2(new_n1208), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT127), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1227), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1316), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1318), .A2(new_n1280), .A3(new_n1314), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1309), .ZN(new_n1320));
  AND3_X1   g1120(.A1(new_n1317), .A2(new_n1319), .A3(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1320), .B1(new_n1317), .B2(new_n1319), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1321), .A2(new_n1322), .ZN(G402));
endmodule


