

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584;

  XOR2_X1 U326 ( .A(G29GAT), .B(G43GAT), .Z(n294) );
  XOR2_X1 U327 ( .A(n428), .B(n427), .Z(n295) );
  XOR2_X1 U328 ( .A(KEYINPUT58), .B(n565), .Z(n296) );
  INV_X1 U329 ( .A(G176GAT), .ZN(n352) );
  NOR2_X1 U330 ( .A1(n529), .A2(n507), .ZN(n508) );
  XNOR2_X1 U331 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U332 ( .A(n355), .B(n354), .ZN(n356) );
  INV_X1 U333 ( .A(KEYINPUT48), .ZN(n514) );
  NOR2_X1 U334 ( .A1(n463), .A2(n582), .ZN(n464) );
  NOR2_X1 U335 ( .A1(n414), .A2(n413), .ZN(n415) );
  XNOR2_X1 U336 ( .A(n515), .B(n514), .ZN(n546) );
  XOR2_X1 U337 ( .A(n435), .B(n434), .Z(n568) );
  XNOR2_X1 U338 ( .A(n371), .B(n370), .ZN(n552) );
  XOR2_X1 U339 ( .A(KEYINPUT16), .B(KEYINPUT82), .Z(n328) );
  XOR2_X1 U340 ( .A(KEYINPUT80), .B(KEYINPUT15), .Z(n298) );
  XNOR2_X1 U341 ( .A(G64GAT), .B(KEYINPUT14), .ZN(n297) );
  XNOR2_X1 U342 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U343 ( .A(G22GAT), .B(G155GAT), .Z(n396) );
  XOR2_X1 U344 ( .A(G78GAT), .B(n396), .Z(n300) );
  XOR2_X1 U345 ( .A(G15GAT), .B(G127GAT), .Z(n355) );
  XNOR2_X1 U346 ( .A(G1GAT), .B(n355), .ZN(n299) );
  XNOR2_X1 U347 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U348 ( .A(n302), .B(n301), .Z(n304) );
  NAND2_X1 U349 ( .A1(G231GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U351 ( .A(n305), .B(KEYINPUT81), .Z(n308) );
  XNOR2_X1 U352 ( .A(G8GAT), .B(G183GAT), .ZN(n306) );
  XNOR2_X1 U353 ( .A(n306), .B(G211GAT), .ZN(n373) );
  XNOR2_X1 U354 ( .A(n373), .B(KEYINPUT12), .ZN(n307) );
  XNOR2_X1 U355 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U356 ( .A(KEYINPUT72), .B(KEYINPUT73), .Z(n310) );
  XNOR2_X1 U357 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n309) );
  XNOR2_X1 U358 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U359 ( .A(G57GAT), .B(n311), .ZN(n448) );
  XNOR2_X1 U360 ( .A(n312), .B(n448), .ZN(n578) );
  XOR2_X1 U361 ( .A(G36GAT), .B(G190GAT), .Z(n377) );
  XOR2_X1 U362 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n314) );
  XNOR2_X1 U363 ( .A(G92GAT), .B(KEYINPUT9), .ZN(n313) );
  XNOR2_X1 U364 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U365 ( .A(n377), .B(n315), .Z(n318) );
  XNOR2_X1 U366 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n316) );
  XNOR2_X1 U367 ( .A(n294), .B(n316), .ZN(n428) );
  XOR2_X1 U368 ( .A(G50GAT), .B(G162GAT), .Z(n397) );
  XNOR2_X1 U369 ( .A(n428), .B(n397), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U371 ( .A(n319), .B(KEYINPUT79), .Z(n321) );
  XOR2_X1 U372 ( .A(G99GAT), .B(G85GAT), .Z(n439) );
  XNOR2_X1 U373 ( .A(G218GAT), .B(n439), .ZN(n320) );
  XNOR2_X1 U374 ( .A(n321), .B(n320), .ZN(n326) );
  XOR2_X1 U375 ( .A(G106GAT), .B(KEYINPUT64), .Z(n323) );
  NAND2_X1 U376 ( .A1(G232GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U377 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U378 ( .A(G134GAT), .B(n324), .Z(n325) );
  XNOR2_X1 U379 ( .A(n326), .B(n325), .ZN(n529) );
  INV_X1 U380 ( .A(n529), .ZN(n564) );
  NAND2_X1 U381 ( .A1(n578), .A2(n564), .ZN(n327) );
  XNOR2_X1 U382 ( .A(n328), .B(n327), .ZN(n416) );
  XOR2_X1 U383 ( .A(KEYINPUT84), .B(G134GAT), .Z(n330) );
  XNOR2_X1 U384 ( .A(KEYINPUT83), .B(G120GAT), .ZN(n329) );
  XNOR2_X1 U385 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U386 ( .A(KEYINPUT0), .B(n331), .Z(n369) );
  XOR2_X1 U387 ( .A(KEYINPUT95), .B(KEYINPUT93), .Z(n333) );
  XNOR2_X1 U388 ( .A(G57GAT), .B(KEYINPUT94), .ZN(n332) );
  XNOR2_X1 U389 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U390 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n335) );
  XNOR2_X1 U391 ( .A(KEYINPUT92), .B(KEYINPUT6), .ZN(n334) );
  XNOR2_X1 U392 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U393 ( .A(n337), .B(n336), .Z(n350) );
  XOR2_X1 U394 ( .A(KEYINPUT2), .B(KEYINPUT89), .Z(n339) );
  XNOR2_X1 U395 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n338) );
  XNOR2_X1 U396 ( .A(n339), .B(n338), .ZN(n390) );
  XOR2_X1 U397 ( .A(n390), .B(KEYINPUT4), .Z(n341) );
  NAND2_X1 U398 ( .A1(G225GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U399 ( .A(n341), .B(n340), .ZN(n348) );
  XOR2_X1 U400 ( .A(G85GAT), .B(G148GAT), .Z(n343) );
  XNOR2_X1 U401 ( .A(G127GAT), .B(G155GAT), .ZN(n342) );
  XNOR2_X1 U402 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U403 ( .A(n344), .B(G162GAT), .Z(n346) );
  XOR2_X1 U404 ( .A(G113GAT), .B(G1GAT), .Z(n427) );
  XNOR2_X1 U405 ( .A(G29GAT), .B(n427), .ZN(n345) );
  XNOR2_X1 U406 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U407 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U408 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U409 ( .A(n369), .B(n351), .ZN(n549) );
  NAND2_X1 U410 ( .A1(G227GAT), .A2(G233GAT), .ZN(n353) );
  XOR2_X1 U411 ( .A(n356), .B(G190GAT), .Z(n361) );
  XOR2_X1 U412 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n358) );
  XNOR2_X1 U413 ( .A(KEYINPUT86), .B(KEYINPUT18), .ZN(n357) );
  XNOR2_X1 U414 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U415 ( .A(G169GAT), .B(n359), .Z(n383) );
  XNOR2_X1 U416 ( .A(G43GAT), .B(n383), .ZN(n360) );
  XNOR2_X1 U417 ( .A(n361), .B(n360), .ZN(n365) );
  XOR2_X1 U418 ( .A(KEYINPUT85), .B(KEYINPUT20), .Z(n363) );
  XNOR2_X1 U419 ( .A(G99GAT), .B(KEYINPUT87), .ZN(n362) );
  XNOR2_X1 U420 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U421 ( .A(n365), .B(n364), .Z(n371) );
  XOR2_X1 U422 ( .A(KEYINPUT88), .B(G71GAT), .Z(n367) );
  XNOR2_X1 U423 ( .A(G113GAT), .B(G183GAT), .ZN(n366) );
  XNOR2_X1 U424 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U425 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U426 ( .A(G197GAT), .B(G218GAT), .ZN(n372) );
  XNOR2_X1 U427 ( .A(n372), .B(KEYINPUT21), .ZN(n391) );
  XNOR2_X1 U428 ( .A(n391), .B(n373), .ZN(n381) );
  XOR2_X1 U429 ( .A(G92GAT), .B(G64GAT), .Z(n375) );
  XNOR2_X1 U430 ( .A(G176GAT), .B(KEYINPUT75), .ZN(n374) );
  XNOR2_X1 U431 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U432 ( .A(G204GAT), .B(n376), .Z(n447) );
  XOR2_X1 U433 ( .A(n377), .B(n447), .Z(n379) );
  NAND2_X1 U434 ( .A1(G226GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U435 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U436 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U437 ( .A(n383), .B(n382), .ZN(n545) );
  INV_X1 U438 ( .A(n545), .ZN(n497) );
  AND2_X1 U439 ( .A1(n552), .A2(n497), .ZN(n384) );
  XNOR2_X1 U440 ( .A(n384), .B(KEYINPUT97), .ZN(n402) );
  XOR2_X1 U441 ( .A(KEYINPUT22), .B(KEYINPUT91), .Z(n386) );
  XNOR2_X1 U442 ( .A(G204GAT), .B(KEYINPUT23), .ZN(n385) );
  XNOR2_X1 U443 ( .A(n386), .B(n385), .ZN(n401) );
  XOR2_X1 U444 ( .A(KEYINPUT24), .B(KEYINPUT90), .Z(n388) );
  NAND2_X1 U445 ( .A1(G228GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U446 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U447 ( .A(n389), .B(G211GAT), .Z(n393) );
  XNOR2_X1 U448 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U449 ( .A(n393), .B(n392), .ZN(n395) );
  XNOR2_X1 U450 ( .A(G106GAT), .B(G78GAT), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n394), .B(G148GAT), .ZN(n442) );
  XOR2_X1 U452 ( .A(n395), .B(n442), .Z(n399) );
  XNOR2_X1 U453 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U454 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n401), .B(n400), .ZN(n550) );
  NAND2_X1 U456 ( .A1(n402), .A2(n550), .ZN(n404) );
  XNOR2_X1 U457 ( .A(KEYINPUT98), .B(KEYINPUT25), .ZN(n403) );
  XNOR2_X1 U458 ( .A(n404), .B(n403), .ZN(n407) );
  NOR2_X1 U459 ( .A1(n552), .A2(n550), .ZN(n405) );
  XNOR2_X1 U460 ( .A(KEYINPUT26), .B(n405), .ZN(n566) );
  XNOR2_X1 U461 ( .A(KEYINPUT27), .B(n497), .ZN(n409) );
  AND2_X1 U462 ( .A1(n566), .A2(n409), .ZN(n406) );
  NOR2_X1 U463 ( .A1(n407), .A2(n406), .ZN(n408) );
  NOR2_X1 U464 ( .A1(n549), .A2(n408), .ZN(n414) );
  NAND2_X1 U465 ( .A1(n549), .A2(n409), .ZN(n516) );
  XNOR2_X1 U466 ( .A(KEYINPUT28), .B(KEYINPUT65), .ZN(n410) );
  XNOR2_X1 U467 ( .A(n410), .B(n550), .ZN(n519) );
  NOR2_X1 U468 ( .A1(n516), .A2(n519), .ZN(n411) );
  XOR2_X1 U469 ( .A(KEYINPUT96), .B(n411), .Z(n412) );
  NOR2_X1 U470 ( .A1(n552), .A2(n412), .ZN(n413) );
  XNOR2_X1 U471 ( .A(n415), .B(KEYINPUT99), .ZN(n462) );
  NAND2_X1 U472 ( .A1(n416), .A2(n462), .ZN(n482) );
  XOR2_X1 U473 ( .A(G8GAT), .B(KEYINPUT68), .Z(n418) );
  XNOR2_X1 U474 ( .A(KEYINPUT67), .B(KEYINPUT30), .ZN(n417) );
  XNOR2_X1 U475 ( .A(n418), .B(n417), .ZN(n435) );
  XOR2_X1 U476 ( .A(G15GAT), .B(G36GAT), .Z(n420) );
  XNOR2_X1 U477 ( .A(G169GAT), .B(G50GAT), .ZN(n419) );
  XNOR2_X1 U478 ( .A(n420), .B(n419), .ZN(n424) );
  XOR2_X1 U479 ( .A(KEYINPUT29), .B(G141GAT), .Z(n422) );
  XNOR2_X1 U480 ( .A(G197GAT), .B(G22GAT), .ZN(n421) );
  XNOR2_X1 U481 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U482 ( .A(n424), .B(n423), .Z(n433) );
  XOR2_X1 U483 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n426) );
  XNOR2_X1 U484 ( .A(KEYINPUT71), .B(KEYINPUT66), .ZN(n425) );
  XNOR2_X1 U485 ( .A(n426), .B(n425), .ZN(n431) );
  NAND2_X1 U486 ( .A1(G229GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U487 ( .A(n295), .B(n429), .ZN(n430) );
  XNOR2_X1 U488 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U490 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n437) );
  XNOR2_X1 U491 ( .A(KEYINPUT33), .B(KEYINPUT32), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U493 ( .A(n438), .B(KEYINPUT31), .Z(n441) );
  XNOR2_X1 U494 ( .A(G120GAT), .B(n439), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n446) );
  XOR2_X1 U496 ( .A(n442), .B(KEYINPUT74), .Z(n444) );
  NAND2_X1 U497 ( .A1(G230GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U499 ( .A(n446), .B(n445), .Z(n450) );
  XOR2_X1 U500 ( .A(n448), .B(n447), .Z(n449) );
  XNOR2_X1 U501 ( .A(n450), .B(n449), .ZN(n574) );
  NOR2_X1 U502 ( .A1(n568), .A2(n574), .ZN(n451) );
  XOR2_X1 U503 ( .A(KEYINPUT78), .B(n451), .Z(n465) );
  NOR2_X1 U504 ( .A1(n482), .A2(n465), .ZN(n452) );
  XNOR2_X1 U505 ( .A(n452), .B(KEYINPUT100), .ZN(n459) );
  NAND2_X1 U506 ( .A1(n459), .A2(n549), .ZN(n453) );
  XNOR2_X1 U507 ( .A(n453), .B(KEYINPUT34), .ZN(n454) );
  XNOR2_X1 U508 ( .A(G1GAT), .B(n454), .ZN(G1324GAT) );
  NAND2_X1 U509 ( .A1(n459), .A2(n497), .ZN(n455) );
  XNOR2_X1 U510 ( .A(n455), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U511 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n457) );
  NAND2_X1 U512 ( .A1(n552), .A2(n459), .ZN(n456) );
  XNOR2_X1 U513 ( .A(n457), .B(n456), .ZN(n458) );
  XOR2_X1 U514 ( .A(G15GAT), .B(n458), .Z(G1326GAT) );
  NAND2_X1 U515 ( .A1(n459), .A2(n519), .ZN(n460) );
  XNOR2_X1 U516 ( .A(n460), .B(KEYINPUT102), .ZN(n461) );
  XNOR2_X1 U517 ( .A(G22GAT), .B(n461), .ZN(G1327GAT) );
  XOR2_X1 U518 ( .A(KEYINPUT103), .B(KEYINPUT39), .Z(n469) );
  INV_X1 U519 ( .A(n578), .ZN(n541) );
  NAND2_X1 U520 ( .A1(n541), .A2(n462), .ZN(n463) );
  XNOR2_X1 U521 ( .A(KEYINPUT36), .B(n564), .ZN(n582) );
  XNOR2_X1 U522 ( .A(n464), .B(KEYINPUT37), .ZN(n492) );
  NOR2_X1 U523 ( .A1(n492), .A2(n465), .ZN(n466) );
  XNOR2_X1 U524 ( .A(n466), .B(KEYINPUT38), .ZN(n467) );
  XNOR2_X2 U525 ( .A(KEYINPUT104), .B(n467), .ZN(n478) );
  NAND2_X1 U526 ( .A1(n478), .A2(n549), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n469), .B(n468), .ZN(n470) );
  XOR2_X1 U528 ( .A(n470), .B(G29GAT), .Z(G1328GAT) );
  XOR2_X1 U529 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n472) );
  NAND2_X1 U530 ( .A1(n478), .A2(n497), .ZN(n471) );
  XNOR2_X1 U531 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U532 ( .A(G36GAT), .B(n473), .ZN(G1329GAT) );
  XNOR2_X1 U533 ( .A(G43GAT), .B(KEYINPUT108), .ZN(n477) );
  XOR2_X1 U534 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n475) );
  NAND2_X1 U535 ( .A1(n478), .A2(n552), .ZN(n474) );
  XNOR2_X1 U536 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U537 ( .A(n477), .B(n476), .ZN(G1330GAT) );
  XOR2_X1 U538 ( .A(G50GAT), .B(KEYINPUT109), .Z(n480) );
  NAND2_X1 U539 ( .A1(n478), .A2(n519), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n480), .B(n479), .ZN(G1331GAT) );
  XNOR2_X1 U541 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n484) );
  XOR2_X1 U542 ( .A(n574), .B(KEYINPUT41), .Z(n535) );
  NAND2_X1 U543 ( .A1(n535), .A2(n568), .ZN(n481) );
  XNOR2_X1 U544 ( .A(n481), .B(KEYINPUT110), .ZN(n493) );
  NOR2_X1 U545 ( .A1(n493), .A2(n482), .ZN(n487) );
  NAND2_X1 U546 ( .A1(n487), .A2(n549), .ZN(n483) );
  XNOR2_X1 U547 ( .A(n484), .B(n483), .ZN(G1332GAT) );
  NAND2_X1 U548 ( .A1(n487), .A2(n497), .ZN(n485) );
  XNOR2_X1 U549 ( .A(n485), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U550 ( .A1(n487), .A2(n552), .ZN(n486) );
  XNOR2_X1 U551 ( .A(n486), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U552 ( .A(KEYINPUT112), .B(KEYINPUT43), .Z(n489) );
  NAND2_X1 U553 ( .A1(n487), .A2(n519), .ZN(n488) );
  XNOR2_X1 U554 ( .A(n489), .B(n488), .ZN(n491) );
  XOR2_X1 U555 ( .A(G78GAT), .B(KEYINPUT111), .Z(n490) );
  XNOR2_X1 U556 ( .A(n491), .B(n490), .ZN(G1335GAT) );
  NOR2_X1 U557 ( .A1(n493), .A2(n492), .ZN(n494) );
  XOR2_X1 U558 ( .A(KEYINPUT113), .B(n494), .Z(n500) );
  NAND2_X1 U559 ( .A1(n549), .A2(n500), .ZN(n495) );
  XNOR2_X1 U560 ( .A(n495), .B(KEYINPUT114), .ZN(n496) );
  XNOR2_X1 U561 ( .A(G85GAT), .B(n496), .ZN(G1336GAT) );
  NAND2_X1 U562 ( .A1(n500), .A2(n497), .ZN(n498) );
  XNOR2_X1 U563 ( .A(n498), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U564 ( .A1(n500), .A2(n552), .ZN(n499) );
  XNOR2_X1 U565 ( .A(n499), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U566 ( .A1(n519), .A2(n500), .ZN(n501) );
  XNOR2_X1 U567 ( .A(n501), .B(KEYINPUT44), .ZN(n502) );
  XNOR2_X1 U568 ( .A(G106GAT), .B(n502), .ZN(G1339GAT) );
  INV_X1 U569 ( .A(n568), .ZN(n520) );
  NAND2_X1 U570 ( .A1(n520), .A2(n535), .ZN(n505) );
  XOR2_X1 U571 ( .A(KEYINPUT46), .B(KEYINPUT117), .Z(n503) );
  XNOR2_X1 U572 ( .A(KEYINPUT116), .B(n503), .ZN(n504) );
  XNOR2_X1 U573 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U574 ( .A(n578), .B(KEYINPUT115), .ZN(n560) );
  NAND2_X1 U575 ( .A1(n506), .A2(n560), .ZN(n507) );
  XNOR2_X1 U576 ( .A(n508), .B(KEYINPUT47), .ZN(n513) );
  NOR2_X1 U577 ( .A1(n582), .A2(n541), .ZN(n509) );
  XOR2_X1 U578 ( .A(KEYINPUT45), .B(n509), .Z(n510) );
  NOR2_X1 U579 ( .A1(n574), .A2(n510), .ZN(n511) );
  NAND2_X1 U580 ( .A1(n511), .A2(n568), .ZN(n512) );
  NAND2_X1 U581 ( .A1(n513), .A2(n512), .ZN(n515) );
  NOR2_X1 U582 ( .A1(n546), .A2(n516), .ZN(n533) );
  NAND2_X1 U583 ( .A1(n552), .A2(n533), .ZN(n517) );
  XNOR2_X1 U584 ( .A(KEYINPUT118), .B(n517), .ZN(n518) );
  NOR2_X1 U585 ( .A1(n519), .A2(n518), .ZN(n530) );
  NAND2_X1 U586 ( .A1(n530), .A2(n520), .ZN(n521) );
  XNOR2_X1 U587 ( .A(G113GAT), .B(n521), .ZN(G1340GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT119), .B(KEYINPUT49), .Z(n523) );
  NAND2_X1 U589 ( .A1(n530), .A2(n535), .ZN(n522) );
  XNOR2_X1 U590 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U591 ( .A(G120GAT), .B(n524), .Z(G1341GAT) );
  INV_X1 U592 ( .A(n530), .ZN(n525) );
  NOR2_X1 U593 ( .A1(n560), .A2(n525), .ZN(n527) );
  XNOR2_X1 U594 ( .A(KEYINPUT50), .B(KEYINPUT120), .ZN(n526) );
  XNOR2_X1 U595 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U596 ( .A(G127GAT), .B(n528), .Z(G1342GAT) );
  XOR2_X1 U597 ( .A(G134GAT), .B(KEYINPUT51), .Z(n532) );
  NAND2_X1 U598 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n532), .B(n531), .ZN(G1343GAT) );
  NAND2_X1 U600 ( .A1(n533), .A2(n566), .ZN(n543) );
  NOR2_X1 U601 ( .A1(n568), .A2(n543), .ZN(n534) );
  XOR2_X1 U602 ( .A(G141GAT), .B(n534), .Z(G1344GAT) );
  INV_X1 U603 ( .A(n535), .ZN(n555) );
  NOR2_X1 U604 ( .A1(n555), .A2(n543), .ZN(n540) );
  XOR2_X1 U605 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n537) );
  XNOR2_X1 U606 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n536) );
  XNOR2_X1 U607 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U608 ( .A(KEYINPUT53), .B(n538), .ZN(n539) );
  XNOR2_X1 U609 ( .A(n540), .B(n539), .ZN(G1345GAT) );
  NOR2_X1 U610 ( .A1(n541), .A2(n543), .ZN(n542) );
  XOR2_X1 U611 ( .A(G155GAT), .B(n542), .Z(G1346GAT) );
  NOR2_X1 U612 ( .A1(n564), .A2(n543), .ZN(n544) );
  XOR2_X1 U613 ( .A(G162GAT), .B(n544), .Z(G1347GAT) );
  NOR2_X1 U614 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U615 ( .A(KEYINPUT54), .B(n547), .Z(n548) );
  NOR2_X1 U616 ( .A1(n549), .A2(n548), .ZN(n567) );
  NAND2_X1 U617 ( .A1(n567), .A2(n550), .ZN(n551) );
  XNOR2_X1 U618 ( .A(KEYINPUT55), .B(n551), .ZN(n553) );
  NAND2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n563) );
  NOR2_X1 U620 ( .A1(n568), .A2(n563), .ZN(n554) );
  XOR2_X1 U621 ( .A(G169GAT), .B(n554), .Z(G1348GAT) );
  NOR2_X1 U622 ( .A1(n563), .A2(n555), .ZN(n559) );
  XOR2_X1 U623 ( .A(KEYINPUT56), .B(KEYINPUT123), .Z(n557) );
  XNOR2_X1 U624 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  NOR2_X1 U627 ( .A1(n563), .A2(n560), .ZN(n561) );
  XOR2_X1 U628 ( .A(KEYINPUT124), .B(n561), .Z(n562) );
  XNOR2_X1 U629 ( .A(G183GAT), .B(n562), .ZN(G1350GAT) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(G190GAT), .B(n296), .ZN(G1351GAT) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n581) );
  NOR2_X1 U633 ( .A1(n568), .A2(n581), .ZN(n573) );
  XOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n570) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(KEYINPUT125), .B(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n576) );
  INV_X1 U640 ( .A(n581), .ZN(n579) );
  NAND2_X1 U641 ( .A1(n579), .A2(n574), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U643 ( .A(G204GAT), .B(n577), .Z(G1353GAT) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U647 ( .A(KEYINPUT62), .B(n583), .Z(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

