

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n594, n595, n596, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765;

  BUF_X1 U371 ( .A(G101), .Z(n349) );
  XNOR2_X1 U372 ( .A(n465), .B(G472), .ZN(n538) );
  XNOR2_X1 U373 ( .A(n442), .B(n358), .ZN(n524) );
  AND2_X2 U374 ( .A1(n663), .A2(n632), .ZN(n701) );
  XNOR2_X2 U375 ( .A(n630), .B(n604), .ZN(n663) );
  XNOR2_X1 U376 ( .A(n350), .B(n363), .ZN(n362) );
  XNOR2_X1 U377 ( .A(n461), .B(n482), .ZN(n350) );
  XNOR2_X2 U378 ( .A(n351), .B(KEYINPUT108), .ZN(n760) );
  NAND2_X2 U379 ( .A1(n397), .A2(n396), .ZN(n351) );
  XNOR2_X2 U380 ( .A(n352), .B(KEYINPUT105), .ZN(n599) );
  NAND2_X2 U381 ( .A1(n591), .A2(n592), .ZN(n352) );
  AND2_X2 U382 ( .A1(n676), .A2(G478), .ZN(n652) );
  NOR2_X1 U383 ( .A1(G953), .A2(G237), .ZN(n496) );
  NOR2_X1 U384 ( .A1(n574), .A2(n573), .ZN(n691) );
  XOR2_X1 U385 ( .A(n434), .B(n447), .Z(n353) );
  AND2_X2 U386 ( .A1(n390), .A2(n388), .ZN(n387) );
  AND2_X2 U387 ( .A1(n524), .A2(n710), .ZN(n454) );
  NOR2_X1 U388 ( .A1(n468), .A2(n374), .ZN(n585) );
  OR2_X1 U389 ( .A1(n638), .A2(n621), .ZN(n486) );
  AND2_X2 U390 ( .A1(n635), .A2(n634), .ZN(n676) );
  XNOR2_X1 U391 ( .A(n381), .B(KEYINPUT40), .ZN(n568) );
  NOR2_X1 U392 ( .A1(n393), .A2(KEYINPUT47), .ZN(n571) );
  XNOR2_X1 U393 ( .A(n726), .B(KEYINPUT77), .ZN(n393) );
  XNOR2_X1 U394 ( .A(n509), .B(n508), .ZN(n694) );
  NAND2_X1 U395 ( .A1(n590), .A2(n716), .ZN(n403) );
  NAND2_X1 U396 ( .A1(n454), .A2(n564), .ZN(n529) );
  XNOR2_X1 U397 ( .A(n448), .B(G104), .ZN(n481) );
  NOR2_X1 U398 ( .A1(n747), .A2(n633), .ZN(n703) );
  AND2_X1 U399 ( .A1(n606), .A2(n605), .ZN(n608) );
  NAND2_X1 U400 ( .A1(n545), .A2(n544), .ZN(n548) );
  AND2_X1 U401 ( .A1(n400), .A2(n398), .ZN(n397) );
  BUF_X1 U402 ( .A(n592), .Z(n567) );
  AND2_X1 U403 ( .A1(n368), .A2(n590), .ZN(n591) );
  NOR2_X1 U404 ( .A1(n529), .A2(n560), .ZN(n383) );
  XNOR2_X1 U405 ( .A(n453), .B(G469), .ZN(n564) );
  XNOR2_X1 U406 ( .A(n395), .B(n507), .ZN(n554) );
  XNOR2_X1 U407 ( .A(n429), .B(n428), .ZN(n674) );
  XNOR2_X1 U408 ( .A(n481), .B(n480), .ZN(n371) );
  XNOR2_X1 U409 ( .A(n470), .B(n511), .ZN(n493) );
  XNOR2_X1 U410 ( .A(KEYINPUT70), .B(KEYINPUT16), .ZN(n479) );
  XNOR2_X1 U411 ( .A(KEYINPUT68), .B(G101), .ZN(n471) );
  INV_X1 U412 ( .A(KEYINPUT64), .ZN(n430) );
  XNOR2_X1 U413 ( .A(G110), .B(G107), .ZN(n448) );
  XNOR2_X1 U414 ( .A(n371), .B(n482), .ZN(n754) );
  NOR2_X1 U415 ( .A1(n674), .A2(G902), .ZN(n442) );
  XNOR2_X1 U416 ( .A(n499), .B(G137), .ZN(n447) );
  XNOR2_X1 U417 ( .A(n431), .B(KEYINPUT8), .ZN(n489) );
  INV_X1 U418 ( .A(n703), .ZN(n634) );
  AND2_X1 U419 ( .A1(n760), .A2(n419), .ZN(n418) );
  NOR2_X1 U420 ( .A1(n588), .A2(n587), .ZN(n419) );
  INV_X1 U421 ( .A(KEYINPUT44), .ZN(n380) );
  NOR2_X1 U422 ( .A1(n389), .A2(n603), .ZN(n388) );
  NOR2_X1 U423 ( .A1(n699), .A2(KEYINPUT81), .ZN(n389) );
  XNOR2_X1 U424 ( .A(G116), .B(G107), .ZN(n491) );
  XNOR2_X1 U425 ( .A(G131), .B(G122), .ZN(n500) );
  XNOR2_X1 U426 ( .A(n414), .B(n413), .ZN(n412) );
  XNOR2_X1 U427 ( .A(KEYINPUT94), .B(KEYINPUT12), .ZN(n414) );
  XNOR2_X1 U428 ( .A(G113), .B(G104), .ZN(n413) );
  XOR2_X1 U429 ( .A(G143), .B(KEYINPUT11), .Z(n498) );
  XNOR2_X1 U430 ( .A(n493), .B(n446), .ZN(n462) );
  XNOR2_X1 U431 ( .A(KEYINPUT4), .B(G131), .ZN(n446) );
  NOR2_X1 U432 ( .A1(n524), .A2(n562), .ZN(n590) );
  NAND2_X1 U433 ( .A1(n646), .A2(n504), .ZN(n395) );
  OR2_X1 U434 ( .A1(n678), .A2(G902), .ZN(n453) );
  XNOR2_X1 U435 ( .A(G110), .B(G128), .ZN(n433) );
  XNOR2_X1 U436 ( .A(n664), .B(n437), .ZN(n373) );
  XNOR2_X1 U437 ( .A(G119), .B(KEYINPUT23), .ZN(n436) );
  XNOR2_X1 U438 ( .A(KEYINPUT24), .B(KEYINPUT69), .ZN(n435) );
  XNOR2_X1 U439 ( .A(n462), .B(n447), .ZN(n665) );
  NAND2_X1 U440 ( .A1(n405), .A2(n408), .ZN(n404) );
  INV_X1 U441 ( .A(KEYINPUT78), .ZN(n408) );
  AND2_X1 U442 ( .A1(n399), .A2(n596), .ZN(n398) );
  NAND2_X1 U443 ( .A1(n595), .A2(KEYINPUT36), .ZN(n399) );
  NOR2_X1 U444 ( .A1(n552), .A2(n741), .ZN(n377) );
  XNOR2_X1 U445 ( .A(n467), .B(n375), .ZN(n374) );
  INV_X1 U446 ( .A(KEYINPUT30), .ZN(n375) );
  XNOR2_X1 U447 ( .A(n611), .B(n528), .ZN(n552) );
  INV_X1 U448 ( .A(KEYINPUT88), .ZN(n528) );
  XNOR2_X1 U449 ( .A(n427), .B(n426), .ZN(n653) );
  NOR2_X1 U450 ( .A1(n489), .A2(n488), .ZN(n426) );
  XNOR2_X1 U451 ( .A(n493), .B(n376), .ZN(n427) );
  AND2_X1 U452 ( .A1(n580), .A2(n579), .ZN(n581) );
  INV_X1 U453 ( .A(KEYINPUT46), .ZN(n417) );
  XNOR2_X1 U454 ( .A(G902), .B(KEYINPUT15), .ZN(n626) );
  XNOR2_X1 U455 ( .A(n463), .B(n421), .ZN(n420) );
  XNOR2_X1 U456 ( .A(KEYINPUT93), .B(KEYINPUT92), .ZN(n463) );
  XNOR2_X1 U457 ( .A(G137), .B(KEYINPUT5), .ZN(n421) );
  XNOR2_X1 U458 ( .A(n423), .B(n422), .ZN(n482) );
  XNOR2_X1 U459 ( .A(G116), .B(G113), .ZN(n422) );
  XNOR2_X1 U460 ( .A(n424), .B(KEYINPUT3), .ZN(n423) );
  INV_X1 U461 ( .A(G119), .ZN(n424) );
  NAND2_X1 U462 ( .A1(n379), .A2(n355), .ZN(n618) );
  XNOR2_X1 U463 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n474) );
  XNOR2_X1 U464 ( .A(KEYINPUT18), .B(KEYINPUT73), .ZN(n473) );
  NAND2_X1 U465 ( .A1(n386), .A2(n385), .ZN(n384) );
  INV_X1 U466 ( .A(KEYINPUT81), .ZN(n385) );
  NAND2_X1 U467 ( .A1(G234), .A2(G237), .ZN(n455) );
  INV_X1 U468 ( .A(G237), .ZN(n466) );
  INV_X1 U469 ( .A(KEYINPUT72), .ZN(n382) );
  AND2_X1 U470 ( .A1(n716), .A2(n720), .ZN(n467) );
  INV_X1 U471 ( .A(G902), .ZN(n504) );
  XNOR2_X1 U472 ( .A(n362), .B(n462), .ZN(n655) );
  XNOR2_X1 U473 ( .A(n420), .B(n464), .ZN(n363) );
  XNOR2_X1 U474 ( .A(n492), .B(n356), .ZN(n376) );
  XNOR2_X1 U475 ( .A(n491), .B(n490), .ZN(n492) );
  INV_X1 U476 ( .A(G122), .ZN(n490) );
  XNOR2_X1 U477 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U478 ( .A(n664), .B(n412), .ZN(n411) );
  XNOR2_X1 U479 ( .A(n500), .B(n499), .ZN(n501) );
  INV_X1 U480 ( .A(KEYINPUT28), .ZN(n402) );
  XNOR2_X1 U481 ( .A(n523), .B(n522), .ZN(n539) );
  INV_X1 U482 ( .A(KEYINPUT97), .ZN(n394) );
  AND2_X1 U483 ( .A1(n589), .A2(n539), .ZN(n545) );
  XNOR2_X1 U484 ( .A(n563), .B(KEYINPUT1), .ZN(n707) );
  AND2_X1 U485 ( .A1(n634), .A2(G472), .ZN(n365) );
  XNOR2_X1 U486 ( .A(n655), .B(KEYINPUT62), .ZN(n656) );
  XNOR2_X1 U487 ( .A(n373), .B(n353), .ZN(n429) );
  AND2_X1 U488 ( .A1(n634), .A2(G475), .ZN(n367) );
  XOR2_X1 U489 ( .A(n646), .B(KEYINPUT59), .Z(n647) );
  XNOR2_X1 U490 ( .A(n665), .B(n452), .ZN(n678) );
  AND2_X1 U491 ( .A1(n634), .A2(G210), .ZN(n366) );
  XNOR2_X1 U492 ( .A(n638), .B(n637), .ZN(n639) );
  INV_X1 U493 ( .A(G140), .ZN(n499) );
  INV_X1 U494 ( .A(G134), .ZN(n511) );
  XNOR2_X1 U495 ( .A(n557), .B(n556), .ZN(n607) );
  XNOR2_X1 U496 ( .A(n586), .B(KEYINPUT106), .ZN(n765) );
  NAND2_X1 U497 ( .A1(n357), .A2(n585), .ZN(n586) );
  NOR2_X1 U498 ( .A1(n707), .A2(n610), .ZN(n354) );
  AND2_X1 U499 ( .A1(n617), .A2(n616), .ZN(n355) );
  XNOR2_X1 U500 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n356) );
  AND2_X1 U501 ( .A1(n584), .A2(n583), .ZN(n357) );
  XOR2_X1 U502 ( .A(n441), .B(n440), .Z(n358) );
  XNOR2_X1 U503 ( .A(n495), .B(n494), .ZN(n532) );
  AND2_X1 U504 ( .A1(n594), .A2(n409), .ZN(n359) );
  XOR2_X1 U505 ( .A(n518), .B(KEYINPUT0), .Z(n360) );
  XOR2_X1 U506 ( .A(n553), .B(KEYINPUT34), .Z(n361) );
  INV_X1 U507 ( .A(KEYINPUT36), .ZN(n409) );
  XNOR2_X1 U508 ( .A(n411), .B(n503), .ZN(n646) );
  INV_X1 U509 ( .A(KEYINPUT76), .ZN(n369) );
  NAND2_X1 U510 ( .A1(n365), .A2(n635), .ZN(n657) );
  NAND2_X1 U511 ( .A1(n366), .A2(n635), .ZN(n640) );
  NAND2_X1 U512 ( .A1(n367), .A2(n635), .ZN(n648) );
  XNOR2_X1 U513 ( .A(n599), .B(n410), .ZN(n401) );
  XNOR2_X2 U514 ( .A(n618), .B(KEYINPUT45), .ZN(n632) );
  INV_X1 U515 ( .A(n564), .ZN(n563) );
  XNOR2_X1 U516 ( .A(n383), .B(n382), .ZN(n468) );
  XNOR2_X1 U517 ( .A(n538), .B(KEYINPUT6), .ZN(n589) );
  INV_X1 U518 ( .A(n589), .ZN(n368) );
  XNOR2_X1 U519 ( .A(n403), .B(n402), .ZN(n565) );
  OR2_X1 U520 ( .A1(n691), .A2(n369), .ZN(n576) );
  BUF_X1 U521 ( .A(n524), .Z(n370) );
  XNOR2_X2 U522 ( .A(n594), .B(KEYINPUT19), .ZN(n573) );
  XNOR2_X2 U523 ( .A(n372), .B(n360), .ZN(n611) );
  NOR2_X2 U524 ( .A1(n573), .A2(n517), .ZN(n372) );
  XNOR2_X1 U525 ( .A(n570), .B(n417), .ZN(n416) );
  NAND2_X2 U526 ( .A1(n387), .A2(n384), .ZN(n630) );
  XNOR2_X1 U527 ( .A(n554), .B(n394), .ZN(n534) );
  XNOR2_X2 U528 ( .A(n536), .B(KEYINPUT99), .ZN(n592) );
  XNOR2_X1 U529 ( .A(n377), .B(n361), .ZN(n555) );
  XNOR2_X2 U530 ( .A(n378), .B(KEYINPUT84), .ZN(n594) );
  NOR2_X2 U531 ( .A1(n601), .A2(n512), .ZN(n378) );
  XNOR2_X1 U532 ( .A(n609), .B(n380), .ZN(n379) );
  NAND2_X1 U533 ( .A1(n568), .A2(n569), .ZN(n570) );
  NAND2_X1 U534 ( .A1(n510), .A2(n567), .ZN(n381) );
  XNOR2_X1 U535 ( .A(n487), .B(KEYINPUT39), .ZN(n510) );
  INV_X1 U536 ( .A(n392), .ZN(n386) );
  NAND2_X1 U537 ( .A1(n392), .A2(n391), .ZN(n390) );
  AND2_X1 U538 ( .A1(n699), .A2(KEYINPUT81), .ZN(n391) );
  XNOR2_X2 U539 ( .A(n415), .B(n425), .ZN(n392) );
  OR2_X1 U540 ( .A1(n613), .A2(n393), .ZN(n615) );
  INV_X1 U541 ( .A(n534), .ZN(n533) );
  NAND2_X1 U542 ( .A1(n401), .A2(n359), .ZN(n400) );
  OR2_X1 U543 ( .A1(n401), .A2(n409), .ZN(n396) );
  NAND2_X2 U544 ( .A1(n406), .A2(n404), .ZN(n635) );
  INV_X1 U545 ( .A(n701), .ZN(n405) );
  AND2_X2 U546 ( .A1(n407), .A2(n629), .ZN(n406) );
  NAND2_X1 U547 ( .A1(n701), .A2(n623), .ZN(n407) );
  INV_X1 U548 ( .A(KEYINPUT107), .ZN(n410) );
  XNOR2_X2 U549 ( .A(n472), .B(KEYINPUT10), .ZN(n664) );
  XNOR2_X2 U550 ( .A(G125), .B(G146), .ZN(n472) );
  NAND2_X1 U551 ( .A1(n418), .A2(n416), .ZN(n415) );
  INV_X1 U552 ( .A(KEYINPUT48), .ZN(n425) );
  INV_X1 U553 ( .A(n568), .ZN(n662) );
  NOR2_X1 U554 ( .A1(n489), .A2(n432), .ZN(n428) );
  XNOR2_X2 U555 ( .A(n430), .B(G953), .ZN(n666) );
  INV_X1 U556 ( .A(n454), .ZN(n706) );
  NAND2_X1 U557 ( .A1(n666), .A2(G234), .ZN(n431) );
  INV_X1 U558 ( .A(G221), .ZN(n432) );
  XNOR2_X1 U559 ( .A(n433), .B(KEYINPUT90), .ZN(n434) );
  XNOR2_X1 U560 ( .A(n436), .B(n435), .ZN(n437) );
  NAND2_X1 U561 ( .A1(n626), .A2(G234), .ZN(n439) );
  XOR2_X1 U562 ( .A(KEYINPUT20), .B(KEYINPUT91), .Z(n438) );
  XNOR2_X1 U563 ( .A(n439), .B(n438), .ZN(n443) );
  NAND2_X1 U564 ( .A1(n443), .A2(G217), .ZN(n441) );
  INV_X1 U565 ( .A(KEYINPUT25), .ZN(n440) );
  NAND2_X1 U566 ( .A1(n443), .A2(G221), .ZN(n445) );
  INV_X1 U567 ( .A(KEYINPUT21), .ZN(n444) );
  XNOR2_X1 U568 ( .A(n445), .B(n444), .ZN(n710) );
  XNOR2_X2 U569 ( .A(G143), .B(G128), .ZN(n470) );
  XNOR2_X1 U570 ( .A(n471), .B(G146), .ZN(n461) );
  XNOR2_X1 U571 ( .A(n481), .B(n461), .ZN(n451) );
  NAND2_X1 U572 ( .A1(n666), .A2(G227), .ZN(n449) );
  XNOR2_X1 U573 ( .A(n449), .B(KEYINPUT89), .ZN(n450) );
  XNOR2_X1 U574 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U575 ( .A(n455), .B(KEYINPUT14), .ZN(n459) );
  NAND2_X1 U576 ( .A1(G902), .A2(n459), .ZN(n513) );
  NOR2_X1 U577 ( .A1(G900), .A2(n513), .ZN(n456) );
  INV_X1 U578 ( .A(n666), .ZN(n642) );
  AND2_X1 U579 ( .A1(n456), .A2(n642), .ZN(n458) );
  INV_X1 U580 ( .A(KEYINPUT104), .ZN(n457) );
  XNOR2_X1 U581 ( .A(n458), .B(n457), .ZN(n460) );
  NAND2_X1 U582 ( .A1(G952), .A2(n459), .ZN(n739) );
  OR2_X1 U583 ( .A1(n739), .A2(G953), .ZN(n515) );
  AND2_X1 U584 ( .A1(n460), .A2(n515), .ZN(n560) );
  NAND2_X1 U585 ( .A1(n496), .A2(G210), .ZN(n464) );
  NAND2_X1 U586 ( .A1(n655), .A2(n504), .ZN(n465) );
  BUF_X2 U587 ( .A(n538), .Z(n716) );
  NAND2_X1 U588 ( .A1(n504), .A2(n466), .ZN(n484) );
  AND2_X1 U589 ( .A1(n484), .A2(G214), .ZN(n512) );
  INV_X1 U590 ( .A(n512), .ZN(n720) );
  NAND2_X1 U591 ( .A1(n666), .A2(G224), .ZN(n469) );
  XNOR2_X1 U592 ( .A(n470), .B(n469), .ZN(n478) );
  XNOR2_X1 U593 ( .A(n472), .B(n471), .ZN(n476) );
  XNOR2_X1 U594 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U595 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U596 ( .A(n477), .B(n478), .ZN(n483) );
  XNOR2_X1 U597 ( .A(n479), .B(G122), .ZN(n480) );
  XNOR2_X1 U598 ( .A(n754), .B(n483), .ZN(n638) );
  INV_X1 U599 ( .A(n626), .ZN(n621) );
  NAND2_X1 U600 ( .A1(n484), .A2(G210), .ZN(n485) );
  XNOR2_X2 U601 ( .A(n486), .B(n485), .ZN(n601) );
  XNOR2_X1 U602 ( .A(n601), .B(KEYINPUT38), .ZN(n721) );
  NAND2_X1 U603 ( .A1(n585), .A2(n721), .ZN(n487) );
  INV_X1 U604 ( .A(G217), .ZN(n488) );
  NAND2_X1 U605 ( .A1(n653), .A2(n504), .ZN(n495) );
  XNOR2_X1 U606 ( .A(KEYINPUT98), .B(G478), .ZN(n494) );
  NAND2_X1 U607 ( .A1(G214), .A2(n496), .ZN(n497) );
  XNOR2_X1 U608 ( .A(n498), .B(n497), .ZN(n502) );
  XOR2_X1 U609 ( .A(KEYINPUT13), .B(KEYINPUT96), .Z(n506) );
  XNOR2_X1 U610 ( .A(KEYINPUT95), .B(G475), .ZN(n505) );
  XOR2_X1 U611 ( .A(n506), .B(n505), .Z(n507) );
  NAND2_X1 U612 ( .A1(n532), .A2(n533), .ZN(n509) );
  INV_X1 U613 ( .A(KEYINPUT100), .ZN(n508) );
  AND2_X1 U614 ( .A1(n510), .A2(n694), .ZN(n603) );
  XNOR2_X1 U615 ( .A(n603), .B(n511), .ZN(G36) );
  INV_X1 U616 ( .A(G898), .ZN(n751) );
  NAND2_X1 U617 ( .A1(G953), .A2(n751), .ZN(n755) );
  OR2_X1 U618 ( .A1(n513), .A2(n755), .ZN(n514) );
  NAND2_X1 U619 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X1 U620 ( .A(n516), .B(KEYINPUT87), .ZN(n517) );
  INV_X1 U621 ( .A(KEYINPUT86), .ZN(n518) );
  OR2_X1 U622 ( .A1(n532), .A2(n554), .ZN(n724) );
  INV_X1 U623 ( .A(n710), .ZN(n561) );
  NOR2_X1 U624 ( .A1(n724), .A2(n561), .ZN(n519) );
  XNOR2_X1 U625 ( .A(n519), .B(KEYINPUT102), .ZN(n520) );
  NAND2_X1 U626 ( .A1(n611), .A2(n520), .ZN(n523) );
  INV_X1 U627 ( .A(KEYINPUT66), .ZN(n521) );
  XNOR2_X1 U628 ( .A(n521), .B(KEYINPUT22), .ZN(n522) );
  INV_X1 U629 ( .A(n539), .ZN(n527) );
  NOR2_X1 U630 ( .A1(n716), .A2(n370), .ZN(n525) );
  NAND2_X1 U631 ( .A1(n707), .A2(n525), .ZN(n526) );
  OR2_X1 U632 ( .A1(n527), .A2(n526), .ZN(n605) );
  XNOR2_X1 U633 ( .A(n605), .B(G110), .ZN(G12) );
  INV_X1 U634 ( .A(n552), .ZN(n531) );
  NOR2_X1 U635 ( .A1(n716), .A2(n529), .ZN(n530) );
  AND2_X1 U636 ( .A1(n531), .A2(n530), .ZN(n683) );
  INV_X1 U637 ( .A(n532), .ZN(n535) );
  NAND2_X1 U638 ( .A1(n535), .A2(n534), .ZN(n536) );
  NAND2_X1 U639 ( .A1(n683), .A2(n592), .ZN(n537) );
  XNOR2_X1 U640 ( .A(n537), .B(G104), .ZN(G6) );
  INV_X1 U641 ( .A(n545), .ZN(n540) );
  XNOR2_X1 U642 ( .A(n540), .B(KEYINPUT83), .ZN(n542) );
  AND2_X1 U643 ( .A1(n707), .A2(n370), .ZN(n541) );
  NAND2_X1 U644 ( .A1(n542), .A2(n541), .ZN(n616) );
  XNOR2_X1 U645 ( .A(n616), .B(n349), .ZN(G3) );
  OR2_X1 U646 ( .A1(n707), .A2(n370), .ZN(n543) );
  XNOR2_X1 U647 ( .A(n543), .B(KEYINPUT103), .ZN(n544) );
  INV_X1 U648 ( .A(KEYINPUT65), .ZN(n546) );
  XNOR2_X1 U649 ( .A(n546), .B(KEYINPUT32), .ZN(n547) );
  XNOR2_X2 U650 ( .A(n548), .B(n547), .ZN(n606) );
  XNOR2_X1 U651 ( .A(n606), .B(G119), .ZN(G21) );
  OR2_X1 U652 ( .A1(n589), .A2(n706), .ZN(n549) );
  OR2_X1 U653 ( .A1(n549), .A2(n707), .ZN(n551) );
  INV_X1 U654 ( .A(KEYINPUT33), .ZN(n550) );
  XNOR2_X1 U655 ( .A(n551), .B(n550), .ZN(n741) );
  INV_X1 U656 ( .A(KEYINPUT74), .ZN(n553) );
  AND2_X1 U657 ( .A1(n554), .A2(n532), .ZN(n584) );
  NAND2_X1 U658 ( .A1(n555), .A2(n584), .ZN(n557) );
  INV_X1 U659 ( .A(KEYINPUT35), .ZN(n556) );
  XOR2_X1 U660 ( .A(G122), .B(KEYINPUT125), .Z(n558) );
  XNOR2_X1 U661 ( .A(n607), .B(n558), .ZN(G24) );
  NAND2_X1 U662 ( .A1(n721), .A2(n720), .ZN(n727) );
  NOR2_X1 U663 ( .A1(n727), .A2(n724), .ZN(n559) );
  XNOR2_X1 U664 ( .A(n559), .B(KEYINPUT41), .ZN(n740) );
  OR2_X1 U665 ( .A1(n561), .A2(n560), .ZN(n562) );
  NAND2_X1 U666 ( .A1(n565), .A2(n564), .ZN(n574) );
  NOR2_X1 U667 ( .A1(n740), .A2(n574), .ZN(n566) );
  XNOR2_X1 U668 ( .A(n566), .B(KEYINPUT42), .ZN(n764) );
  INV_X1 U669 ( .A(n764), .ZN(n569) );
  OR2_X2 U670 ( .A1(n592), .A2(n694), .ZN(n726) );
  XNOR2_X1 U671 ( .A(n571), .B(KEYINPUT71), .ZN(n572) );
  NAND2_X1 U672 ( .A1(n572), .A2(KEYINPUT76), .ZN(n575) );
  NAND2_X1 U673 ( .A1(n575), .A2(n691), .ZN(n582) );
  NAND2_X1 U674 ( .A1(n576), .A2(n726), .ZN(n577) );
  NAND2_X1 U675 ( .A1(n577), .A2(KEYINPUT47), .ZN(n580) );
  INV_X1 U676 ( .A(KEYINPUT47), .ZN(n578) );
  NAND2_X1 U677 ( .A1(n578), .A2(n369), .ZN(n579) );
  NAND2_X1 U678 ( .A1(n582), .A2(n581), .ZN(n588) );
  INV_X1 U679 ( .A(n601), .ZN(n583) );
  INV_X1 U680 ( .A(n765), .ZN(n587) );
  INV_X1 U681 ( .A(n594), .ZN(n595) );
  INV_X1 U682 ( .A(n707), .ZN(n596) );
  AND2_X1 U683 ( .A1(n707), .A2(n720), .ZN(n598) );
  NAND2_X1 U684 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U685 ( .A(n600), .B(KEYINPUT43), .ZN(n602) );
  NAND2_X1 U686 ( .A1(n602), .A2(n601), .ZN(n699) );
  INV_X1 U687 ( .A(KEYINPUT80), .ZN(n604) );
  NAND2_X1 U688 ( .A1(n608), .A2(n607), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n716), .A2(n454), .ZN(n610) );
  NAND2_X1 U690 ( .A1(n611), .A2(n354), .ZN(n612) );
  XNOR2_X1 U691 ( .A(n612), .B(KEYINPUT31), .ZN(n695) );
  NOR2_X1 U692 ( .A1(n695), .A2(n683), .ZN(n613) );
  INV_X1 U693 ( .A(KEYINPUT101), .ZN(n614) );
  XNOR2_X1 U694 ( .A(n615), .B(n614), .ZN(n617) );
  NAND2_X1 U695 ( .A1(KEYINPUT2), .A2(KEYINPUT79), .ZN(n619) );
  NAND2_X1 U696 ( .A1(n619), .A2(KEYINPUT78), .ZN(n620) );
  NOR2_X1 U697 ( .A1(n621), .A2(n620), .ZN(n628) );
  INV_X1 U698 ( .A(n628), .ZN(n622) );
  AND2_X1 U699 ( .A1(KEYINPUT78), .A2(n622), .ZN(n623) );
  INV_X1 U700 ( .A(KEYINPUT2), .ZN(n624) );
  NOR2_X1 U701 ( .A1(n624), .A2(KEYINPUT79), .ZN(n625) );
  NOR2_X1 U702 ( .A1(n626), .A2(n625), .ZN(n627) );
  OR2_X1 U703 ( .A1(n628), .A2(n627), .ZN(n629) );
  INV_X1 U704 ( .A(n630), .ZN(n631) );
  NAND2_X1 U705 ( .A1(n631), .A2(KEYINPUT2), .ZN(n633) );
  INV_X1 U706 ( .A(n632), .ZN(n747) );
  XNOR2_X1 U707 ( .A(KEYINPUT85), .B(KEYINPUT54), .ZN(n636) );
  XOR2_X1 U708 ( .A(n636), .B(KEYINPUT55), .Z(n637) );
  XNOR2_X1 U709 ( .A(n640), .B(n639), .ZN(n643) );
  INV_X1 U710 ( .A(G952), .ZN(n641) );
  NAND2_X1 U711 ( .A1(n642), .A2(n641), .ZN(n658) );
  NAND2_X1 U712 ( .A1(n643), .A2(n658), .ZN(n645) );
  XOR2_X1 U713 ( .A(KEYINPUT82), .B(KEYINPUT56), .Z(n644) );
  XNOR2_X1 U714 ( .A(n645), .B(n644), .ZN(G51) );
  XNOR2_X1 U715 ( .A(n648), .B(n647), .ZN(n649) );
  NAND2_X1 U716 ( .A1(n649), .A2(n658), .ZN(n651) );
  XNOR2_X1 U717 ( .A(KEYINPUT67), .B(KEYINPUT60), .ZN(n650) );
  XNOR2_X1 U718 ( .A(n651), .B(n650), .ZN(G60) );
  XNOR2_X1 U719 ( .A(n652), .B(n653), .ZN(n654) );
  INV_X1 U720 ( .A(n658), .ZN(n681) );
  NOR2_X1 U721 ( .A1(n654), .A2(n681), .ZN(G63) );
  XNOR2_X1 U722 ( .A(n657), .B(n656), .ZN(n659) );
  NAND2_X1 U723 ( .A1(n659), .A2(n658), .ZN(n661) );
  XOR2_X1 U724 ( .A(KEYINPUT109), .B(KEYINPUT63), .Z(n660) );
  XNOR2_X1 U725 ( .A(n661), .B(n660), .ZN(G57) );
  XOR2_X1 U726 ( .A(n662), .B(G131), .Z(G33) );
  XNOR2_X1 U727 ( .A(n665), .B(n664), .ZN(n668) );
  XNOR2_X1 U728 ( .A(n663), .B(n668), .ZN(n667) );
  NAND2_X1 U729 ( .A1(n667), .A2(n666), .ZN(n672) );
  XOR2_X1 U730 ( .A(G227), .B(n668), .Z(n669) );
  NAND2_X1 U731 ( .A1(n669), .A2(G900), .ZN(n670) );
  NAND2_X1 U732 ( .A1(n670), .A2(G953), .ZN(n671) );
  NAND2_X1 U733 ( .A1(n672), .A2(n671), .ZN(G72) );
  NAND2_X1 U734 ( .A1(n676), .A2(G217), .ZN(n673) );
  XNOR2_X1 U735 ( .A(n674), .B(n673), .ZN(n675) );
  NOR2_X1 U736 ( .A1(n675), .A2(n681), .ZN(G66) );
  NAND2_X1 U737 ( .A1(n676), .A2(G469), .ZN(n680) );
  XOR2_X1 U738 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n677) );
  XNOR2_X1 U739 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U740 ( .A(n680), .B(n679), .ZN(n682) );
  NOR2_X1 U741 ( .A1(n682), .A2(n681), .ZN(G54) );
  XNOR2_X1 U742 ( .A(KEYINPUT110), .B(KEYINPUT26), .ZN(n687) );
  NAND2_X1 U743 ( .A1(n683), .A2(n694), .ZN(n685) );
  XOR2_X1 U744 ( .A(G107), .B(KEYINPUT27), .Z(n684) );
  XNOR2_X1 U745 ( .A(n685), .B(n684), .ZN(n686) );
  XNOR2_X1 U746 ( .A(n687), .B(n686), .ZN(G9) );
  XOR2_X1 U747 ( .A(KEYINPUT111), .B(KEYINPUT29), .Z(n689) );
  NAND2_X1 U748 ( .A1(n691), .A2(n694), .ZN(n688) );
  XNOR2_X1 U749 ( .A(n689), .B(n688), .ZN(n690) );
  XOR2_X1 U750 ( .A(G128), .B(n690), .Z(G30) );
  NAND2_X1 U751 ( .A1(n691), .A2(n567), .ZN(n692) );
  XNOR2_X1 U752 ( .A(n692), .B(G146), .ZN(G48) );
  NAND2_X1 U753 ( .A1(n695), .A2(n567), .ZN(n693) );
  XNOR2_X1 U754 ( .A(n693), .B(G113), .ZN(G15) );
  XOR2_X1 U755 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n697) );
  NAND2_X1 U756 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U757 ( .A(n697), .B(n696), .ZN(n698) );
  XNOR2_X1 U758 ( .A(G116), .B(n698), .ZN(G18) );
  XNOR2_X1 U759 ( .A(n699), .B(n499), .ZN(n700) );
  XNOR2_X1 U760 ( .A(n700), .B(KEYINPUT115), .ZN(G42) );
  XNOR2_X1 U761 ( .A(KEYINPUT2), .B(KEYINPUT75), .ZN(n702) );
  AND2_X1 U762 ( .A1(n405), .A2(n702), .ZN(n704) );
  NOR2_X1 U763 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U764 ( .A1(n705), .A2(G953), .ZN(n745) );
  NAND2_X1 U765 ( .A1(n707), .A2(n706), .ZN(n709) );
  XOR2_X1 U766 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n708) );
  XNOR2_X1 U767 ( .A(n709), .B(n708), .ZN(n714) );
  XOR2_X1 U768 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n712) );
  NOR2_X1 U769 ( .A1(n370), .A2(n710), .ZN(n711) );
  XOR2_X1 U770 ( .A(n712), .B(n711), .Z(n713) );
  NAND2_X1 U771 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U772 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U773 ( .A1(n354), .A2(n717), .ZN(n718) );
  XOR2_X1 U774 ( .A(KEYINPUT51), .B(n718), .Z(n719) );
  NOR2_X1 U775 ( .A1(n740), .A2(n719), .ZN(n735) );
  NOR2_X1 U776 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U777 ( .A(n722), .B(KEYINPUT118), .ZN(n723) );
  NOR2_X1 U778 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U779 ( .A(KEYINPUT119), .B(n725), .Z(n731) );
  INV_X1 U780 ( .A(n726), .ZN(n728) );
  NOR2_X1 U781 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U782 ( .A(KEYINPUT120), .B(n729), .ZN(n730) );
  NOR2_X1 U783 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U784 ( .A1(n732), .A2(n741), .ZN(n733) );
  XOR2_X1 U785 ( .A(KEYINPUT121), .B(n733), .Z(n734) );
  NOR2_X1 U786 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U787 ( .A(KEYINPUT122), .B(n736), .Z(n737) );
  XOR2_X1 U788 ( .A(KEYINPUT52), .B(n737), .Z(n738) );
  NOR2_X1 U789 ( .A1(n739), .A2(n738), .ZN(n743) );
  NOR2_X1 U790 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U791 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U792 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U793 ( .A(KEYINPUT53), .B(n746), .Z(G75) );
  NOR2_X1 U794 ( .A1(n747), .A2(G953), .ZN(n753) );
  NAND2_X1 U795 ( .A1(G224), .A2(G953), .ZN(n748) );
  XNOR2_X1 U796 ( .A(n748), .B(KEYINPUT123), .ZN(n749) );
  XNOR2_X1 U797 ( .A(n749), .B(KEYINPUT61), .ZN(n750) );
  NOR2_X1 U798 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U799 ( .A1(n753), .A2(n752), .ZN(n759) );
  XNOR2_X1 U800 ( .A(n754), .B(n349), .ZN(n756) );
  NAND2_X1 U801 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U802 ( .A(n757), .B(KEYINPUT124), .ZN(n758) );
  XNOR2_X1 U803 ( .A(n759), .B(n758), .ZN(G69) );
  XOR2_X1 U804 ( .A(KEYINPUT114), .B(KEYINPUT37), .Z(n762) );
  XNOR2_X1 U805 ( .A(n760), .B(G125), .ZN(n761) );
  XNOR2_X1 U806 ( .A(n762), .B(n761), .ZN(G27) );
  XOR2_X1 U807 ( .A(G137), .B(KEYINPUT126), .Z(n763) );
  XNOR2_X1 U808 ( .A(n764), .B(n763), .ZN(G39) );
  XNOR2_X1 U809 ( .A(G143), .B(n765), .ZN(G45) );
endmodule

