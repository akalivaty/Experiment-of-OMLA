//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 1 0 1 1 1 0 1 0 0 0 0 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT31), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT67), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT2), .ZN(new_n190));
  INV_X1    g004(.A(G113), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n189), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  NAND3_X1  g006(.A1(KEYINPUT67), .A2(KEYINPUT2), .A3(G113), .ZN(new_n193));
  AOI22_X1  g007(.A1(new_n192), .A2(new_n193), .B1(new_n190), .B2(new_n191), .ZN(new_n194));
  INV_X1    g008(.A(G116), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT68), .B1(new_n195), .B2(G119), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT68), .ZN(new_n197));
  INV_X1    g011(.A(G119), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G116), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n195), .A2(G119), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n196), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(new_n194), .B(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(G143), .B(G146), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT1), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(G128), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G143), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n210), .B(G146), .C1(new_n207), .C2(KEYINPUT1), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n206), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n213));
  INV_X1    g027(.A(G137), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n213), .B1(new_n214), .B2(G134), .ZN(new_n215));
  INV_X1    g029(.A(G134), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(KEYINPUT65), .A3(G137), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G131), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT11), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n220), .B1(new_n216), .B2(G137), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n214), .A2(KEYINPUT11), .A3(G134), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n218), .A2(new_n219), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n216), .A2(G137), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n214), .A2(G134), .ZN(new_n225));
  OAI21_X1  g039(.A(G131), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n212), .A2(new_n223), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n208), .A2(G143), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n210), .A2(G146), .ZN(new_n230));
  OR2_X1    g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  NAND2_X1  g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  AOI22_X1  g046(.A1(new_n229), .A2(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n229), .A2(new_n230), .A3(new_n232), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n216), .A2(KEYINPUT65), .A3(G137), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT65), .B1(new_n216), .B2(G137), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n221), .A2(new_n222), .ZN(new_n239));
  OAI21_X1  g053(.A(G131), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n235), .B1(new_n240), .B2(new_n223), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT30), .ZN(new_n242));
  NOR3_X1   g056(.A1(new_n228), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT64), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n245), .B1(new_n233), .B2(new_n234), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n229), .A2(new_n230), .A3(new_n232), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n231), .A2(new_n232), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n247), .B(KEYINPUT64), .C1(new_n248), .C2(new_n204), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n240), .A2(new_n223), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT66), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n252), .B1(new_n250), .B2(new_n251), .ZN(new_n254));
  NOR3_X1   g068(.A1(new_n253), .A2(new_n254), .A3(new_n228), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n203), .B(new_n244), .C1(new_n255), .C2(KEYINPUT30), .ZN(new_n256));
  INV_X1    g070(.A(new_n235), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n251), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(new_n202), .A3(new_n227), .ZN(new_n259));
  NOR2_X1   g073(.A1(G237), .A2(G953), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G210), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n261), .B(G101), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n262), .B(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n256), .A2(new_n259), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT69), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n256), .A2(new_n267), .A3(new_n259), .A4(new_n264), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n188), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n259), .ZN(new_n270));
  INV_X1    g084(.A(new_n254), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n227), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n243), .B1(new_n273), .B2(new_n242), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n270), .B1(new_n274), .B2(new_n203), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(new_n188), .A3(new_n264), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n270), .A2(KEYINPUT28), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT28), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n259), .A2(new_n278), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n277), .B(new_n279), .C1(new_n255), .C2(new_n202), .ZN(new_n280));
  XOR2_X1   g094(.A(new_n264), .B(KEYINPUT70), .Z(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n276), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n187), .B1(new_n269), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT32), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NOR3_X1   g100(.A1(new_n280), .A2(KEYINPUT29), .A3(new_n281), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n203), .B1(new_n228), .B2(new_n241), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT71), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n259), .A3(new_n289), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n258), .A2(KEYINPUT71), .A3(new_n202), .A4(new_n227), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(KEYINPUT28), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT72), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n290), .A2(new_n294), .A3(KEYINPUT28), .A4(new_n291), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n279), .B(KEYINPUT73), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(new_n264), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT29), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n299), .B1(new_n275), .B2(new_n264), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n287), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(G472), .B1(new_n301), .B2(G902), .ZN(new_n302));
  OAI211_X1 g116(.A(KEYINPUT32), .B(new_n187), .C1(new_n269), .C2(new_n283), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n286), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n286), .A2(new_n302), .A3(KEYINPUT74), .A4(new_n303), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G902), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT22), .B(G137), .ZN(new_n310));
  INV_X1    g124(.A(G221), .ZN(new_n311));
  INV_X1    g125(.A(G234), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n311), .A2(new_n312), .A3(G953), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n310), .B(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G140), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G125), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT16), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT76), .B1(new_n315), .B2(G125), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT76), .ZN(new_n321));
  INV_X1    g135(.A(G125), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n322), .A3(G140), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n316), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n319), .B1(new_n325), .B2(KEYINPUT16), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n208), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n320), .A2(new_n323), .B1(G125), .B2(new_n315), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n318), .B1(new_n328), .B2(new_n317), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G146), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n198), .A2(G128), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT23), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT23), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n333), .B1(new_n198), .B2(G128), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n332), .B1(new_n334), .B2(new_n331), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n327), .A2(new_n330), .B1(G110), .B2(new_n335), .ZN(new_n336));
  XOR2_X1   g150(.A(G119), .B(G128), .Z(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT24), .B(G110), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n338), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n340), .B1(new_n335), .B2(G110), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT77), .ZN(new_n342));
  OR2_X1    g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n322), .A2(G140), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n316), .A2(new_n344), .A3(new_n208), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n341), .A2(new_n342), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n343), .A2(new_n345), .A3(new_n330), .A4(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n339), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT78), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n314), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT78), .B1(new_n339), .B2(new_n347), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI211_X1 g166(.A(KEYINPUT78), .B(new_n314), .C1(new_n339), .C2(new_n347), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n309), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT25), .ZN(new_n355));
  OAI21_X1  g169(.A(G217), .B1(new_n312), .B2(G902), .ZN(new_n356));
  XOR2_X1   g170(.A(new_n356), .B(KEYINPUT75), .Z(new_n357));
  INV_X1    g171(.A(KEYINPUT25), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n358), .B(new_n309), .C1(new_n352), .C2(new_n353), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n355), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n357), .A2(G902), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n361), .B1(new_n352), .B2(new_n353), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n308), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT79), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT91), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT20), .ZN(new_n368));
  NOR2_X1   g182(.A1(G475), .A2(G902), .ZN(new_n369));
  XNOR2_X1  g183(.A(G113), .B(G122), .ZN(new_n370));
  INV_X1    g184(.A(G104), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n370), .B(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT19), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n316), .A2(new_n344), .A3(new_n373), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n208), .B(new_n374), .C1(new_n328), .C2(new_n373), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n375), .B1(new_n326), .B2(new_n208), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT88), .ZN(new_n377));
  INV_X1    g191(.A(G237), .ZN(new_n378));
  INV_X1    g192(.A(G953), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(G214), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n210), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n260), .A2(G143), .A3(G214), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G131), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n381), .A2(new_n219), .A3(new_n382), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT88), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n330), .A2(new_n387), .A3(new_n375), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n377), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT86), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n381), .A2(new_n390), .A3(new_n382), .ZN(new_n391));
  NAND2_X1  g205(.A1(KEYINPUT18), .A2(G131), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n392), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n381), .A2(new_n390), .A3(new_n394), .A4(new_n382), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n345), .B1(new_n328), .B2(new_n208), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT87), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n396), .A2(KEYINPUT87), .A3(new_n397), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n372), .B1(new_n389), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n383), .A2(KEYINPUT17), .A3(G131), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT17), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n384), .A2(new_n405), .A3(new_n385), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n327), .A2(new_n404), .A3(new_n330), .A4(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT89), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n372), .B(new_n408), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n396), .A2(KEYINPUT87), .A3(new_n397), .ZN(new_n410));
  AOI21_X1  g224(.A(KEYINPUT87), .B1(new_n396), .B2(new_n397), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n407), .B(new_n409), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n368), .B(new_n369), .C1(new_n403), .C2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n386), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n415), .B1(new_n376), .B2(KEYINPUT88), .ZN(new_n416));
  AOI22_X1  g230(.A1(new_n416), .A2(new_n388), .B1(new_n400), .B2(new_n401), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n412), .B1(new_n417), .B2(new_n372), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n368), .B1(new_n418), .B2(new_n369), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT90), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n414), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n418), .A2(KEYINPUT90), .A3(new_n368), .A4(new_n369), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G475), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n402), .A2(new_n407), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n412), .B1(new_n425), .B2(new_n372), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n424), .B1(new_n426), .B2(new_n309), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n367), .B1(new_n423), .B2(new_n428), .ZN(new_n429));
  AOI211_X1 g243(.A(KEYINPUT91), .B(new_n427), .C1(new_n421), .C2(new_n422), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  XOR2_X1   g245(.A(G116), .B(G122), .Z(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G107), .ZN(new_n433));
  XNOR2_X1  g247(.A(G116), .B(G122), .ZN(new_n434));
  INV_X1    g248(.A(G107), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT92), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(G128), .B(G143), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n216), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(KEYINPUT13), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n210), .A2(G128), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n442), .B(G134), .C1(KEYINPUT13), .C2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n433), .A2(new_n436), .A3(KEYINPUT92), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n439), .A2(new_n441), .A3(new_n444), .A4(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n440), .B(new_n216), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n195), .A2(KEYINPUT14), .A3(G122), .ZN(new_n448));
  OAI211_X1 g262(.A(G107), .B(new_n448), .C1(new_n432), .C2(KEYINPUT14), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n447), .A2(new_n449), .A3(new_n436), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT9), .B(G234), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n452), .A2(G217), .A3(new_n379), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n446), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT93), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT93), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n446), .A2(new_n456), .A3(new_n450), .A4(new_n453), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n453), .B1(new_n446), .B2(new_n450), .ZN(new_n459));
  OR2_X1    g273(.A1(new_n459), .A2(KEYINPUT94), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(KEYINPUT94), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n309), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT95), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n462), .A2(KEYINPUT95), .A3(new_n309), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT15), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(G478), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n463), .A2(new_n470), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n431), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(G214), .B1(G237), .B2(G902), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(G110), .B(G122), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n435), .A2(G104), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n435), .A2(G104), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n479), .B1(KEYINPUT3), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT3), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n482), .A2(new_n435), .A3(G104), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n481), .A2(KEYINPUT80), .A3(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(KEYINPUT3), .B1(new_n371), .B2(G107), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n371), .A2(G107), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n483), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT80), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n484), .A2(G101), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT81), .ZN(new_n491));
  INV_X1    g305(.A(G101), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n481), .A2(new_n491), .A3(new_n492), .A4(new_n483), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n485), .A2(new_n483), .A3(new_n492), .A4(new_n486), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT81), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n490), .A2(new_n496), .A3(KEYINPUT4), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n484), .A2(new_n498), .A3(G101), .A4(new_n489), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n497), .A2(new_n203), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n194), .A2(new_n199), .A3(new_n200), .A4(new_n196), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT5), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(new_n198), .A3(G116), .ZN(new_n504));
  OAI211_X1 g318(.A(G113), .B(new_n504), .C1(new_n201), .C2(new_n503), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n492), .B1(new_n480), .B2(new_n486), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n494), .A2(KEYINPUT81), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n494), .A2(KEYINPUT81), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT82), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT82), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n496), .A2(new_n513), .A3(new_n508), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n506), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n478), .B1(new_n501), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n506), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n513), .B1(new_n496), .B2(new_n508), .ZN(new_n518));
  AOI211_X1 g332(.A(KEYINPUT82), .B(new_n507), .C1(new_n493), .C2(new_n495), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n477), .A3(new_n500), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n516), .A2(KEYINPUT6), .A3(new_n521), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n206), .A2(new_n322), .A3(new_n209), .A4(new_n211), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT84), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n235), .A2(G125), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n379), .A2(G224), .ZN(new_n528));
  XOR2_X1   g342(.A(new_n527), .B(new_n528), .Z(new_n529));
  INV_X1    g343(.A(KEYINPUT6), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n530), .B(new_n478), .C1(new_n501), .C2(new_n515), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n522), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n517), .A2(new_n511), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n477), .B(KEYINPUT8), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n506), .A2(new_n496), .A3(new_n508), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n537), .B1(new_n525), .B2(new_n526), .ZN(new_n538));
  OR2_X1    g352(.A1(new_n523), .A2(KEYINPUT84), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n523), .A2(KEYINPUT84), .ZN(new_n540));
  AND4_X1   g354(.A1(new_n537), .A2(new_n539), .A3(new_n526), .A4(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n536), .B1(new_n538), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT85), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(KEYINPUT85), .B(new_n536), .C1(new_n538), .C2(new_n541), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n545), .A3(new_n521), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n532), .A2(new_n546), .A3(new_n309), .ZN(new_n547));
  OAI21_X1  g361(.A(G210), .B1(G237), .B2(G902), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n532), .A2(new_n546), .A3(new_n309), .A4(new_n548), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n476), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(G234), .A2(G237), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n554), .A2(G952), .A3(new_n379), .ZN(new_n555));
  XOR2_X1   g369(.A(new_n555), .B(KEYINPUT96), .Z(new_n556));
  AND3_X1   g370(.A1(new_n554), .A2(G902), .A3(G953), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT21), .B(G898), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n474), .A2(new_n553), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n363), .B1(new_n306), .B2(new_n307), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT79), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n311), .B1(new_n452), .B2(new_n309), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(G469), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n212), .B(new_n508), .C1(new_n509), .C2(new_n510), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n212), .B1(new_n496), .B2(new_n508), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n251), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT12), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g387(.A(KEYINPUT12), .B(new_n251), .C1(new_n569), .C2(new_n570), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OR2_X1    g389(.A1(new_n569), .A2(KEYINPUT10), .ZN(new_n576));
  OAI211_X1 g390(.A(KEYINPUT10), .B(new_n212), .C1(new_n518), .C2(new_n519), .ZN(new_n577));
  INV_X1    g391(.A(new_n251), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n497), .A2(new_n257), .A3(new_n499), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n576), .A2(new_n577), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(G110), .B(G140), .ZN(new_n582));
  INV_X1    g396(.A(G227), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n583), .A2(G953), .ZN(new_n584));
  XOR2_X1   g398(.A(new_n582), .B(new_n584), .Z(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n251), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n589), .A2(new_n580), .A3(new_n585), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  OR2_X1    g405(.A1(new_n591), .A2(KEYINPUT83), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(KEYINPUT83), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n567), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n585), .B1(new_n589), .B2(new_n580), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n575), .A2(new_n580), .A3(new_n585), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n567), .B(new_n309), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n567), .A2(new_n309), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n566), .B1(new_n594), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n366), .A2(new_n561), .A3(new_n564), .A4(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(G3));
  OAI21_X1  g418(.A(new_n309), .B1(new_n269), .B2(new_n283), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(G472), .ZN(new_n606));
  OR2_X1    g420(.A1(new_n606), .A2(KEYINPUT97), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(KEYINPUT97), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n607), .A2(new_n284), .A3(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(new_n601), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT33), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n462), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n446), .A2(new_n450), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT98), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n453), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(new_n613), .B(new_n615), .Z(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT33), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n618), .A2(G478), .A3(new_n309), .ZN(new_n619));
  INV_X1    g433(.A(new_n467), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n619), .B1(new_n620), .B2(G478), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n621), .B1(new_n429), .B2(new_n430), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT99), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n553), .A2(new_n560), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n621), .B(KEYINPUT99), .C1(new_n429), .C2(new_n430), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n610), .A2(new_n364), .A3(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT34), .B(G104), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G6));
  NAND2_X1  g444(.A1(new_n471), .A2(new_n473), .ZN(new_n631));
  INV_X1    g445(.A(new_n419), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n427), .B1(new_n632), .B2(new_n414), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n625), .A2(new_n634), .A3(new_n364), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n610), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT35), .B(G107), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G9));
  NOR2_X1   g452(.A1(new_n314), .A2(KEYINPUT36), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT100), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n348), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n361), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n360), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n553), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n474), .A2(new_n560), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n610), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT37), .B(G110), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G12));
  AOI21_X1  g462(.A(new_n601), .B1(new_n306), .B2(new_n307), .ZN(new_n649));
  INV_X1    g463(.A(G900), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n557), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n556), .A2(new_n651), .ZN(new_n652));
  AND3_X1   g466(.A1(new_n631), .A2(new_n633), .A3(new_n652), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n644), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n649), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G128), .ZN(G30));
  NAND2_X1  g470(.A1(new_n550), .A2(new_n551), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT38), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n286), .A2(new_n303), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n266), .A2(new_n268), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n281), .A2(new_n291), .A3(new_n290), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g477(.A(G472), .B1(new_n663), .B2(G902), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n652), .B(KEYINPUT39), .Z(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n602), .A2(new_n668), .ZN(new_n669));
  AOI211_X1 g483(.A(new_n659), .B(new_n666), .C1(KEYINPUT40), .C2(new_n669), .ZN(new_n670));
  OR2_X1    g484(.A1(new_n669), .A2(KEYINPUT40), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n631), .B(new_n475), .C1(new_n429), .C2(new_n430), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n670), .A2(new_n643), .A3(new_n671), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G143), .ZN(G45));
  OAI211_X1 g489(.A(new_n621), .B(new_n652), .C1(new_n429), .C2(new_n430), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(KEYINPUT101), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n369), .B1(new_n403), .B2(new_n413), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n420), .B1(new_n678), .B2(KEYINPUT20), .ZN(new_n679));
  INV_X1    g493(.A(new_n414), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n422), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n428), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(KEYINPUT91), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n423), .A2(new_n367), .A3(new_n428), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT101), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n686), .A2(new_n687), .A3(new_n621), .A4(new_n652), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n677), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n689), .A2(new_n649), .A3(new_n644), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT102), .B(G146), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G48));
  NOR2_X1   g506(.A1(new_n595), .A2(new_n596), .ZN(new_n693));
  OAI21_X1  g507(.A(G469), .B1(new_n693), .B2(G902), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n566), .A3(new_n597), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n627), .A2(new_n562), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT41), .B(G113), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G15));
  NAND2_X1  g513(.A1(new_n696), .A2(new_n552), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n700), .B1(new_n306), .B2(new_n307), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n635), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G116), .ZN(G18));
  NAND2_X1  g517(.A1(new_n360), .A2(new_n642), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n701), .A2(new_n704), .A3(new_n645), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G119), .ZN(G21));
  INV_X1    g520(.A(new_n657), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n672), .A2(new_n695), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n661), .A2(KEYINPUT31), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n296), .A2(new_n297), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n281), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n709), .A2(new_n276), .A3(new_n711), .ZN(new_n712));
  XOR2_X1   g526(.A(new_n187), .B(KEYINPUT103), .Z(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n606), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n715), .A2(new_n560), .A3(new_n363), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n708), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G122), .ZN(G24));
  NOR3_X1   g532(.A1(new_n715), .A2(new_n700), .A3(new_n643), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n689), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT104), .B(G125), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G27));
  AND3_X1   g536(.A1(new_n550), .A2(new_n475), .A3(new_n551), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n587), .A2(new_n590), .A3(G469), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n597), .A2(new_n599), .A3(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n723), .A2(KEYINPUT105), .A3(new_n566), .A4(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT105), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n725), .A2(new_n566), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n550), .A2(new_n475), .A3(new_n551), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n677), .A2(new_n688), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n304), .A2(KEYINPUT42), .A3(new_n364), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n689), .A2(new_n562), .A3(new_n731), .ZN(new_n735));
  XOR2_X1   g549(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n736));
  AOI21_X1  g550(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(new_n219), .ZN(G33));
  NAND3_X1  g552(.A1(new_n562), .A2(new_n653), .A3(new_n731), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G134), .ZN(G36));
  NAND2_X1  g554(.A1(new_n431), .A2(new_n621), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n741), .A2(KEYINPUT43), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(KEYINPUT43), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n744), .A2(new_n609), .A3(new_n704), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT44), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n591), .A2(KEYINPUT45), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n591), .B(KEYINPUT83), .ZN(new_n749));
  OAI211_X1 g563(.A(G469), .B(new_n748), .C1(new_n749), .C2(KEYINPUT45), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n599), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT46), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n750), .A2(KEYINPUT46), .A3(new_n599), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(new_n597), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(new_n566), .A3(new_n668), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n745), .A2(new_n746), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n747), .A2(new_n723), .A3(new_n757), .A4(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G137), .ZN(G39));
  INV_X1    g574(.A(KEYINPUT47), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n755), .A2(new_n761), .A3(new_n566), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n761), .B1(new_n755), .B2(new_n566), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n763), .A2(new_n308), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n364), .A2(new_n729), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(new_n689), .A3(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G140), .ZN(G42));
  NOR4_X1   g582(.A1(new_n741), .A2(new_n476), .A3(new_n363), .A4(new_n565), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT107), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n658), .B1(new_n769), .B2(new_n770), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n694), .A2(new_n597), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT49), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(KEYINPUT49), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n665), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n771), .A2(new_n772), .A3(new_n774), .A4(new_n776), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n695), .A2(new_n729), .A3(new_n556), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n744), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n304), .A2(new_n364), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n779), .A2(KEYINPUT48), .A3(new_n781), .ZN(new_n782));
  AOI22_X1  g596(.A1(new_n701), .A2(new_n635), .B1(new_n716), .B2(new_n708), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n697), .A3(new_n705), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n737), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n360), .A2(new_n642), .A3(new_n652), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT109), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT109), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n360), .A2(new_n788), .A3(new_n642), .A4(new_n652), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n728), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n672), .A2(new_n707), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n790), .A2(new_n665), .A3(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n690), .A2(new_n720), .A3(new_n655), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT52), .ZN(new_n794));
  AOI22_X1  g608(.A1(new_n689), .A2(new_n719), .B1(new_n649), .B2(new_n654), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n795), .A2(new_n796), .A3(new_n690), .A4(new_n792), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n785), .A2(new_n739), .A3(new_n794), .A4(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT108), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n471), .A2(new_n799), .A3(new_n473), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n469), .B1(new_n465), .B2(new_n466), .ZN(new_n801));
  OAI21_X1  g615(.A(KEYINPUT108), .B1(new_n801), .B2(new_n472), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n803), .A2(new_n633), .A3(new_n652), .A4(new_n723), .ZN(new_n804));
  AOI211_X1 g618(.A(new_n601), .B(new_n804), .C1(new_n306), .C2(new_n307), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n732), .A2(new_n715), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n704), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n622), .B1(new_n686), .B2(new_n803), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n610), .A2(new_n625), .A3(new_n364), .A4(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n603), .A2(new_n807), .A3(new_n646), .A4(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n798), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT111), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n785), .A2(new_n812), .A3(new_n794), .A4(new_n797), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(KEYINPUT53), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  OAI211_X1 g629(.A(KEYINPUT53), .B(new_n813), .C1(new_n798), .C2(new_n810), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT54), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT110), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n794), .A2(new_n797), .ZN(new_n819));
  AND4_X1   g633(.A1(new_n603), .A2(new_n807), .A3(new_n646), .A4(new_n809), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n819), .A2(new_n739), .A3(new_n820), .A4(new_n785), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n818), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n811), .A2(KEYINPUT110), .A3(KEYINPUT53), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n823), .B(new_n824), .C1(KEYINPUT53), .C2(new_n811), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n817), .B1(new_n825), .B2(KEYINPUT54), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n715), .A2(new_n556), .A3(new_n363), .ZN(new_n827));
  AND4_X1   g641(.A1(new_n696), .A2(new_n742), .A3(new_n743), .A4(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n828), .A2(new_n476), .A3(new_n659), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(KEYINPUT112), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT112), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n828), .A2(new_n831), .A3(new_n476), .A4(new_n659), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT50), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n830), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n828), .A2(KEYINPUT50), .A3(new_n476), .A4(new_n659), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n830), .A2(new_n832), .A3(KEYINPUT113), .A4(new_n833), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  OAI22_X1  g653(.A1(new_n763), .A2(new_n764), .B1(new_n566), .B2(new_n773), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n840), .A2(new_n723), .A3(new_n744), .A4(new_n827), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n779), .A2(new_n606), .A3(new_n704), .A4(new_n714), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n666), .A2(new_n364), .A3(new_n778), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n686), .A2(new_n621), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n839), .A2(new_n843), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT51), .ZN(new_n848));
  INV_X1    g662(.A(new_n841), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n848), .B1(new_n849), .B2(KEYINPUT114), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n847), .B(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n844), .A2(new_n624), .A3(new_n626), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n379), .A2(G952), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(KEYINPUT115), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n744), .A2(new_n827), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n852), .B(new_n854), .C1(new_n855), .C2(new_n700), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(KEYINPUT116), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT48), .B1(new_n779), .B2(new_n781), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AND4_X1   g673(.A1(new_n782), .A2(new_n826), .A3(new_n851), .A4(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(G952), .A2(G953), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n777), .B1(new_n860), .B2(new_n861), .ZN(G75));
  NAND4_X1  g676(.A1(new_n815), .A2(G210), .A3(G902), .A4(new_n816), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT56), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n529), .B(KEYINPUT55), .Z(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n866), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n863), .A2(new_n864), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n522), .A2(new_n531), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(KEYINPUT117), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n379), .A2(G952), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n867), .A2(new_n872), .A3(new_n869), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n874), .A2(new_n876), .A3(new_n877), .ZN(G51));
  XNOR2_X1  g692(.A(new_n598), .B(KEYINPUT57), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n815), .A2(KEYINPUT54), .A3(new_n816), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n879), .B1(new_n881), .B2(new_n817), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT118), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n815), .A2(new_n816), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n880), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n888), .A2(KEYINPUT118), .A3(new_n879), .ZN(new_n889));
  INV_X1    g703(.A(new_n693), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n884), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  OR3_X1    g705(.A1(new_n885), .A2(new_n309), .A3(new_n750), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n875), .B1(new_n891), .B2(new_n892), .ZN(G54));
  INV_X1    g707(.A(KEYINPUT119), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n821), .B(new_n814), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n895), .A2(KEYINPUT58), .A3(G902), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(new_n424), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n894), .B1(new_n897), .B2(new_n418), .ZN(new_n898));
  INV_X1    g712(.A(new_n418), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n899), .B1(new_n896), .B2(new_n424), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n876), .ZN(new_n901));
  NOR4_X1   g715(.A1(new_n896), .A2(KEYINPUT119), .A3(new_n424), .A4(new_n899), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n898), .A2(new_n901), .A3(new_n902), .ZN(G60));
  INV_X1    g717(.A(new_n618), .ZN(new_n904));
  NAND2_X1  g718(.A1(G478), .A2(G902), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT59), .Z(new_n906));
  OAI21_X1  g720(.A(new_n904), .B1(new_n826), .B2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n906), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n618), .B(new_n908), .C1(new_n881), .C2(new_n817), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT120), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n888), .A2(KEYINPUT120), .A3(new_n618), .A4(new_n908), .ZN(new_n912));
  AND4_X1   g726(.A1(new_n876), .A2(new_n907), .A3(new_n911), .A4(new_n912), .ZN(G63));
  NAND2_X1  g727(.A1(G217), .A2(G902), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT60), .Z(new_n915));
  NAND4_X1  g729(.A1(new_n895), .A2(KEYINPUT122), .A3(new_n641), .A4(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n815), .A2(new_n816), .A3(new_n915), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n352), .A2(new_n353), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n875), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n815), .A2(new_n641), .A3(new_n816), .A4(new_n915), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT122), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n916), .A2(new_n919), .A3(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT121), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT61), .ZN(new_n925));
  AOI21_X1  g739(.A(KEYINPUT61), .B1(new_n923), .B2(new_n924), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(G66));
  INV_X1    g741(.A(G224), .ZN(new_n928));
  OAI21_X1  g742(.A(G953), .B1(new_n558), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n603), .A2(new_n646), .A3(new_n809), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n930), .A2(new_n784), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n929), .B1(new_n931), .B2(G953), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n873), .B1(G898), .B2(new_n379), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT123), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n932), .B(new_n934), .ZN(G69));
  AND2_X1   g749(.A1(new_n795), .A2(new_n690), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n674), .A2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT62), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n674), .A2(KEYINPUT62), .A3(new_n936), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n941), .A2(new_n767), .ZN(new_n942));
  AOI211_X1 g756(.A(new_n729), .B(new_n669), .C1(KEYINPUT124), .C2(new_n808), .ZN(new_n943));
  OR2_X1    g757(.A1(new_n808), .A2(KEYINPUT124), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n943), .A2(new_n366), .A3(new_n564), .A4(new_n944), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n759), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(G953), .B1(new_n942), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n374), .B1(new_n328), .B2(new_n373), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n274), .B(new_n948), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n739), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n747), .A2(new_n723), .A3(new_n758), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n781), .A2(new_n791), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n951), .B1(new_n954), .B2(new_n757), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n767), .A2(new_n936), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n956), .A2(new_n737), .ZN(new_n957));
  AOI21_X1  g771(.A(G953), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n379), .A2(G900), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n958), .A2(new_n959), .A3(new_n949), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n961));
  OAI21_X1  g775(.A(G953), .B1(new_n583), .B2(new_n650), .ZN(new_n962));
  OAI22_X1  g776(.A1(new_n950), .A2(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n961), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT126), .Z(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  OAI221_X1 g781(.A(new_n965), .B1(new_n961), .B2(new_n962), .C1(new_n950), .C2(new_n960), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(G72));
  NAND2_X1  g783(.A1(G472), .A2(G902), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT63), .Z(new_n971));
  OAI21_X1  g785(.A(new_n661), .B1(new_n275), .B2(new_n264), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n825), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n275), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n955), .A2(new_n957), .A3(new_n931), .ZN(new_n975));
  AOI211_X1 g789(.A(new_n974), .B(new_n264), .C1(new_n975), .C2(new_n971), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n974), .A2(new_n264), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n942), .A2(new_n931), .A3(new_n946), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n977), .B1(new_n978), .B2(new_n971), .ZN(new_n979));
  NOR4_X1   g793(.A1(new_n973), .A2(new_n976), .A3(new_n979), .A4(new_n875), .ZN(G57));
endmodule


