//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n530, new_n531, new_n532, new_n533, new_n534, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n552,
    new_n553, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n604,
    new_n605, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1160,
    new_n1161, new_n1162;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT64), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT65), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n451), .A2(new_n456), .B1(new_n457), .B2(new_n452), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT66), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n460), .A2(new_n461), .A3(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  OAI21_X1  g041(.A(KEYINPUT67), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n467));
  AND3_X1   g042(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G137), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n463), .A2(G2105), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n471), .B1(new_n476), .B2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n469), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n481));
  NAND4_X1  g056(.A1(new_n467), .A2(new_n462), .A3(G2105), .A4(new_n464), .ZN(new_n482));
  INV_X1    g057(.A(G124), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n484), .B1(new_n468), .B2(G136), .ZN(G162));
  OAI21_X1  g060(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n487), .B1(G114), .B2(new_n466), .ZN(new_n488));
  INV_X1    g063(.A(G126), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n488), .B1(new_n482), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n467), .A2(new_n462), .A3(new_n464), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  NOR3_X1   g070(.A1(new_n492), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n473), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n491), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(G50), .ZN(new_n501));
  AND2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  OR2_X1    g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT5), .B(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n501), .A2(new_n505), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n509), .A2(new_n512), .ZN(G303));
  INV_X1    g088(.A(G303), .ZN(G166));
  XNOR2_X1  g089(.A(KEYINPUT70), .B(KEYINPUT7), .ZN(new_n515));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n515), .B(new_n516), .ZN(new_n517));
  AND3_X1   g092(.A1(new_n504), .A2(G89), .A3(new_n506), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n519), .A2(KEYINPUT71), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(KEYINPUT71), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n522));
  XOR2_X1   g097(.A(KEYINPUT68), .B(G51), .Z(new_n523));
  OAI21_X1  g098(.A(new_n522), .B1(new_n505), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT69), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n524), .A2(new_n525), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n520), .A2(new_n521), .A3(new_n526), .A4(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  INV_X1    g104(.A(G52), .ZN(new_n530));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n530), .A2(new_n505), .B1(new_n507), .B2(new_n531), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n511), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n532), .A2(new_n534), .ZN(G171));
  NAND2_X1  g110(.A1(G68), .A2(G543), .ZN(new_n536));
  XOR2_X1   g111(.A(KEYINPUT5), .B(G543), .Z(new_n537));
  INV_X1    g112(.A(G56), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n511), .B1(new_n539), .B2(KEYINPUT72), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n540), .B1(KEYINPUT72), .B2(new_n539), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n502), .A2(new_n503), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n543), .A2(G81), .B1(new_n545), .B2(G43), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(G860), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT73), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  INV_X1    g129(.A(KEYINPUT74), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G53), .ZN(new_n556));
  OR3_X1    g131(.A1(new_n505), .A2(KEYINPUT9), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT9), .B1(new_n505), .B2(new_n556), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT75), .ZN(new_n559));
  INV_X1    g134(.A(G91), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n507), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n543), .A2(KEYINPUT75), .A3(G91), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n557), .A2(new_n558), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT76), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n511), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n566), .B1(new_n565), .B2(new_n564), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(G299));
  INV_X1    g143(.A(G171), .ZN(G301));
  INV_X1    g144(.A(G49), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT77), .B1(new_n505), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n545), .A2(new_n572), .A3(G49), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  OR2_X1    g149(.A1(new_n506), .A2(G74), .ZN(new_n575));
  AOI22_X1  g150(.A1(G651), .A2(new_n575), .B1(new_n543), .B2(G87), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(G288));
  INV_X1    g152(.A(G48), .ZN(new_n578));
  INV_X1    g153(.A(G86), .ZN(new_n579));
  OAI22_X1  g154(.A1(new_n578), .A2(new_n505), .B1(new_n507), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n506), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n511), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G305));
  AOI22_X1  g159(.A1(new_n543), .A2(G85), .B1(new_n545), .B2(G47), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n511), .B2(new_n586), .ZN(G290));
  INV_X1    g162(.A(G92), .ZN(new_n588));
  XNOR2_X1  g163(.A(KEYINPUT78), .B(KEYINPUT10), .ZN(new_n589));
  OR3_X1    g164(.A1(new_n507), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(G79), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G66), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n537), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n593), .A2(G651), .B1(new_n545), .B2(G54), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n589), .B1(new_n507), .B2(new_n588), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n590), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(G868), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n598), .B1(new_n597), .B2(G171), .ZN(G284));
  OAI21_X1  g174(.A(new_n598), .B1(new_n597), .B2(G171), .ZN(G321));
  NAND2_X1  g175(.A1(G299), .A2(new_n597), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(G168), .B2(new_n597), .ZN(G297));
  OAI21_X1  g177(.A(new_n601), .B1(G168), .B2(new_n597), .ZN(G280));
  INV_X1    g178(.A(new_n596), .ZN(new_n604));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(G860), .ZN(G148));
  NAND2_X1  g181(.A1(new_n547), .A2(new_n597), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n596), .A2(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n597), .B2(new_n608), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g185(.A(new_n482), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G123), .ZN(new_n612));
  OAI21_X1  g187(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n613));
  INV_X1    g188(.A(G111), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n613), .A2(KEYINPUT80), .B1(new_n614), .B2(G2105), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(KEYINPUT80), .B2(new_n613), .ZN(new_n616));
  INV_X1    g191(.A(G135), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n612), .B(new_n616), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n619), .A2(KEYINPUT81), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(KEYINPUT81), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(G2096), .Z(new_n623));
  NAND2_X1  g198(.A1(new_n473), .A2(new_n470), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT12), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2100), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT79), .B(KEYINPUT13), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n623), .A2(new_n628), .ZN(G156));
  XOR2_X1   g204(.A(G1341), .B(G1348), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT83), .ZN(new_n631));
  XOR2_X1   g206(.A(G2451), .B(G2454), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT16), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n631), .B(new_n633), .Z(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT82), .B(KEYINPUT14), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT15), .B(G2435), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2438), .ZN(new_n637));
  XOR2_X1   g212(.A(G2427), .B(G2430), .Z(new_n638));
  AOI21_X1  g213(.A(new_n635), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(new_n637), .B2(new_n638), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n634), .B(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g219(.A(G14), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n645), .B1(new_n644), .B2(new_n642), .ZN(G401));
  XOR2_X1   g221(.A(G2072), .B(G2078), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT17), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  INV_X1    g226(.A(new_n650), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n651), .B1(new_n652), .B2(new_n647), .ZN(new_n653));
  AOI22_X1  g228(.A1(new_n649), .A2(new_n650), .B1(new_n653), .B2(KEYINPUT84), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(KEYINPUT84), .B2(new_n653), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT85), .Z(new_n656));
  INV_X1    g231(.A(new_n647), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n657), .A2(new_n651), .A3(new_n650), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT18), .Z(new_n659));
  NAND3_X1  g234(.A1(new_n648), .A2(new_n651), .A3(new_n652), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n656), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2096), .B(G2100), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XOR2_X1   g238(.A(G1971), .B(G1976), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  XOR2_X1   g241(.A(G1961), .B(G1966), .Z(new_n667));
  AND2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT20), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n666), .A2(new_n667), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n665), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(new_n665), .B2(new_n671), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1991), .B(G1996), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1981), .B(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G229));
  MUX2_X1   g255(.A(G24), .B(G290), .S(G16), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(G1986), .ZN(new_n682));
  INV_X1    g257(.A(G29), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G25), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n468), .A2(KEYINPUT86), .A3(G131), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT86), .ZN(new_n686));
  INV_X1    g261(.A(G131), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(new_n618), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g264(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n690));
  INV_X1    g265(.A(G107), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(G2105), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(new_n611), .B2(G119), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT87), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n684), .B1(new_n695), .B2(new_n683), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT35), .B(G1991), .Z(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n682), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(G16), .A2(G23), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT88), .ZN(new_n701));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n701), .B1(G288), .B2(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT89), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT33), .B(G1976), .Z(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n704), .A2(new_n706), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n702), .A2(G22), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G166), .B2(new_n702), .ZN(new_n710));
  INV_X1    g285(.A(G1971), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(G6), .A2(G16), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n583), .B2(G16), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT32), .B(G1981), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NAND4_X1  g291(.A1(new_n707), .A2(new_n708), .A3(new_n712), .A4(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT34), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n717), .A2(new_n718), .ZN(new_n720));
  OAI221_X1 g295(.A(new_n699), .B1(new_n696), .B2(new_n698), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT36), .ZN(new_n722));
  INV_X1    g297(.A(G2078), .ZN(new_n723));
  NOR2_X1   g298(.A1(G164), .A2(new_n683), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G27), .B2(new_n683), .ZN(new_n725));
  INV_X1    g300(.A(new_n622), .ZN(new_n726));
  AOI22_X1  g301(.A1(new_n723), .A2(new_n725), .B1(new_n726), .B2(G29), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT25), .Z(new_n729));
  INV_X1    g304(.A(G139), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n618), .B2(new_n730), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT91), .Z(new_n732));
  AOI22_X1  g307(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(new_n466), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n735), .A2(new_n683), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n683), .B2(G33), .ZN(new_n737));
  INV_X1    g312(.A(G2072), .ZN(new_n738));
  OAI221_X1 g313(.A(new_n727), .B1(new_n723), .B2(new_n725), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n702), .A2(G21), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G168), .B2(new_n702), .ZN(new_n741));
  INV_X1    g316(.A(G1966), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT24), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n744), .A2(G34), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(G34), .ZN(new_n746));
  AOI21_X1  g321(.A(G29), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n478), .B2(G29), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT92), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n743), .B1(G2084), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(G4), .A2(G16), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n604), .B2(G16), .ZN(new_n752));
  INV_X1    g327(.A(G1348), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT31), .B(G11), .ZN(new_n755));
  INV_X1    g330(.A(G28), .ZN(new_n756));
  AOI21_X1  g331(.A(G29), .B1(new_n756), .B2(KEYINPUT30), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(KEYINPUT95), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(KEYINPUT30), .B2(new_n756), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n757), .A2(KEYINPUT95), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n755), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(G171), .A2(new_n702), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G5), .B2(new_n702), .ZN(new_n763));
  INV_X1    g338(.A(G1961), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n761), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n754), .B(new_n765), .C1(new_n764), .C2(new_n763), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n702), .A2(G19), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n541), .A2(new_n546), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n768), .B2(new_n702), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1341), .ZN(new_n770));
  NOR4_X1   g345(.A1(new_n739), .A2(new_n750), .A3(new_n766), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n702), .A2(G20), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT23), .Z(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G299), .B2(G16), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT98), .B(G1956), .Z(new_n775));
  XOR2_X1   g350(.A(new_n774), .B(new_n775), .Z(new_n776));
  NAND2_X1  g351(.A1(new_n683), .A2(G26), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT28), .ZN(new_n778));
  OAI21_X1  g353(.A(KEYINPUT90), .B1(G104), .B2(G2105), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  NOR3_X1   g355(.A1(KEYINPUT90), .A2(G104), .A3(G2105), .ZN(new_n781));
  OAI221_X1 g356(.A(G2104), .B1(G116), .B2(new_n466), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(G128), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(new_n482), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G140), .B2(new_n468), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n778), .B1(new_n785), .B2(new_n683), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G2067), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G2084), .B2(new_n749), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n771), .A2(new_n776), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n683), .A2(G35), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT96), .Z(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G162), .B2(new_n683), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT29), .Z(new_n793));
  INV_X1    g368(.A(G2090), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT97), .Z(new_n796));
  NAND2_X1  g371(.A1(new_n683), .A2(G32), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n470), .A2(G105), .ZN(new_n798));
  NAND3_X1  g373(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT93), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT26), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n468), .A2(G141), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n611), .A2(G129), .ZN(new_n803));
  AND4_X1   g378(.A1(new_n798), .A2(new_n801), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT94), .Z(new_n805));
  OAI21_X1  g380(.A(new_n797), .B1(new_n805), .B2(new_n683), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT27), .B(G1996), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n737), .A2(new_n738), .B1(new_n794), .B2(new_n793), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n796), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n789), .A2(new_n810), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n722), .A2(new_n811), .ZN(G311));
  NAND2_X1  g387(.A1(new_n722), .A2(new_n811), .ZN(G150));
  NAND2_X1  g388(.A1(new_n604), .A2(G559), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT38), .ZN(new_n815));
  INV_X1    g390(.A(G55), .ZN(new_n816));
  INV_X1    g391(.A(G93), .ZN(new_n817));
  OAI22_X1  g392(.A1(new_n816), .A2(new_n505), .B1(new_n507), .B2(new_n817), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n819), .A2(new_n511), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n768), .A2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n821), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n547), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n815), .B(new_n825), .Z(new_n826));
  OR2_X1    g401(.A1(new_n826), .A2(KEYINPUT39), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(KEYINPUT39), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n827), .A2(new_n548), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n821), .A2(new_n548), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT37), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(G145));
  XOR2_X1   g407(.A(new_n805), .B(new_n785), .Z(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n835));
  INV_X1    g410(.A(G118), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n835), .A2(KEYINPUT101), .B1(new_n836), .B2(G2105), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(KEYINPUT101), .B2(new_n835), .ZN(new_n838));
  INV_X1    g413(.A(G130), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n838), .B1(new_n839), .B2(new_n482), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(new_n468), .B2(G142), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n694), .A2(new_n625), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n694), .A2(new_n625), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n842), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n845), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n847), .A2(new_n841), .A3(new_n843), .ZN(new_n848));
  INV_X1    g423(.A(new_n735), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n846), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n849), .B1(new_n846), .B2(new_n848), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT99), .ZN(new_n853));
  AOI221_X4 g428(.A(new_n853), .B1(new_n473), .B2(new_n496), .C1(new_n494), .C2(KEYINPUT4), .ZN(new_n854));
  AOI21_X1  g429(.A(KEYINPUT99), .B1(new_n495), .B2(new_n497), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n491), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(KEYINPUT100), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT100), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n858), .B(new_n491), .C1(new_n854), .C2(new_n855), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NOR3_X1   g435(.A1(new_n851), .A2(new_n852), .A3(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n860), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n846), .A2(new_n848), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(new_n735), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n862), .B1(new_n864), .B2(new_n850), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n834), .B1(new_n861), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT102), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n860), .B1(new_n851), .B2(new_n852), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n864), .A2(new_n862), .A3(new_n850), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n868), .A2(new_n833), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n866), .A2(new_n867), .A3(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n622), .B(new_n478), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(G162), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(G37), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n866), .A2(new_n867), .A3(new_n873), .A4(new_n870), .ZN(new_n876));
  XNOR2_X1  g451(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n877));
  AND3_X1   g452(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n877), .B1(new_n875), .B2(new_n876), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(G395));
  XNOR2_X1  g455(.A(G303), .B(KEYINPUT105), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(G305), .ZN(new_n882));
  XOR2_X1   g457(.A(G288), .B(G290), .Z(new_n883));
  INV_X1    g458(.A(KEYINPUT106), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n883), .A2(new_n884), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n882), .A2(new_n887), .A3(new_n885), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  OR3_X1    g464(.A1(new_n889), .A2(KEYINPUT107), .A3(KEYINPUT42), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT41), .ZN(new_n891));
  NOR2_X1   g466(.A1(G299), .A2(new_n604), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n892), .A2(KEYINPUT104), .ZN(new_n893));
  NAND2_X1  g468(.A1(G299), .A2(new_n604), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n563), .A2(KEYINPUT104), .A3(new_n567), .A4(new_n596), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n891), .B1(new_n893), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n892), .A2(KEYINPUT104), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n899), .A2(new_n896), .A3(KEYINPUT41), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n825), .B(new_n608), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n899), .A2(new_n896), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n903), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT42), .B1(new_n889), .B2(KEYINPUT107), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n890), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n905), .B1(new_n890), .B2(new_n906), .ZN(new_n908));
  OAI21_X1  g483(.A(G868), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(G868), .B2(new_n821), .ZN(G295));
  OAI21_X1  g485(.A(new_n909), .B1(G868), .B2(new_n821), .ZN(G331));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n912));
  INV_X1    g487(.A(new_n824), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n547), .A2(new_n823), .ZN(new_n914));
  OAI21_X1  g489(.A(G171), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n822), .A2(G301), .A3(new_n824), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(G286), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n915), .A2(G168), .A3(new_n916), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n918), .B(new_n919), .C1(new_n898), .C2(new_n900), .ZN(new_n920));
  INV_X1    g495(.A(new_n919), .ZN(new_n921));
  AOI21_X1  g496(.A(G168), .B1(new_n915), .B2(new_n916), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n904), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n920), .A2(new_n923), .A3(KEYINPUT108), .ZN(new_n924));
  AOI21_X1  g499(.A(G37), .B1(new_n924), .B2(new_n889), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n886), .A2(new_n888), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n926), .A2(new_n920), .A3(KEYINPUT108), .A4(new_n923), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n912), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT109), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT44), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n924), .A2(new_n889), .ZN(new_n931));
  INV_X1    g506(.A(G37), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n932), .A3(new_n927), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n925), .A2(new_n912), .A3(new_n927), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n930), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n934), .A2(new_n929), .A3(KEYINPUT44), .A4(new_n935), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(G397));
  XNOR2_X1  g514(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n940));
  INV_X1    g515(.A(G1384), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n940), .B1(new_n860), .B2(new_n941), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n469), .A2(new_n477), .A3(G40), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(KEYINPUT111), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n785), .B(G2067), .ZN(new_n946));
  INV_X1    g521(.A(G1996), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n946), .B1(new_n805), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n944), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n950), .A2(new_n947), .A3(new_n805), .ZN(new_n951));
  INV_X1    g526(.A(new_n945), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n694), .B(new_n697), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n949), .B(new_n951), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(G290), .B(G1986), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n954), .B1(new_n950), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT49), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n583), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(G1981), .B1(new_n582), .B2(KEYINPUT114), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT49), .B1(new_n580), .B2(new_n582), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n943), .A2(new_n941), .A3(new_n856), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n580), .A2(new_n582), .A3(KEYINPUT49), .ZN(new_n964));
  INV_X1    g539(.A(new_n582), .ZN(new_n965));
  AOI22_X1  g540(.A1(new_n543), .A2(G86), .B1(new_n545), .B2(G48), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n957), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n959), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n962), .A2(new_n963), .A3(new_n968), .A4(G8), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n574), .A2(G1976), .A3(new_n576), .ZN(new_n970));
  INV_X1    g545(.A(G1976), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT52), .B1(G288), .B2(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n963), .A2(new_n970), .A3(new_n972), .A4(G8), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n963), .A2(new_n970), .A3(G8), .ZN(new_n975));
  OR2_X1    g550(.A1(new_n975), .A2(KEYINPUT113), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n977), .B1(new_n975), .B2(KEYINPUT113), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n974), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(G303), .A2(G8), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n980), .B(KEYINPUT55), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT50), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n856), .A2(new_n983), .A3(new_n941), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n943), .ZN(new_n985));
  AOI22_X1  g560(.A1(new_n494), .A2(KEYINPUT4), .B1(new_n473), .B2(new_n496), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n941), .B1(new_n986), .B2(new_n490), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n987), .A2(KEYINPUT112), .A3(KEYINPUT50), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT112), .B1(new_n987), .B2(KEYINPUT50), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n985), .A2(new_n990), .A3(G2090), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n992), .A2(G1384), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n857), .A2(new_n859), .A3(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n469), .A2(new_n477), .A3(G40), .ZN(new_n995));
  INV_X1    g570(.A(new_n940), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n995), .B1(new_n987), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(G1971), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n982), .B(G8), .C1(new_n991), .C2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G8), .ZN(new_n1000));
  INV_X1    g575(.A(new_n998), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n943), .B1(KEYINPUT50), .B2(new_n987), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n983), .B1(new_n856), .B2(new_n941), .ZN(new_n1003));
  OR3_X1    g578(.A1(new_n1002), .A2(new_n1003), .A3(G2090), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1000), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n979), .B(new_n999), .C1(new_n1005), .C2(new_n982), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT120), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(new_n985), .B2(new_n990), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n987), .A2(KEYINPUT50), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT112), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n987), .A2(KEYINPUT112), .A3(KEYINPUT50), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1013), .A2(KEYINPUT120), .A3(new_n943), .A4(new_n984), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1008), .A2(new_n764), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n856), .A2(new_n941), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n995), .B1(new_n1016), .B2(new_n992), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n499), .A2(KEYINPUT116), .A3(new_n941), .A4(new_n940), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n941), .B(new_n940), .C1(new_n986), .C2(new_n490), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT116), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1017), .A2(KEYINPUT53), .A3(new_n723), .A4(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n994), .A2(new_n997), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1024), .B1(new_n1025), .B2(G2078), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1015), .A2(new_n1023), .A3(new_n1026), .A4(G301), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n1027), .A2(KEYINPUT54), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n994), .A2(KEYINPUT53), .A3(new_n723), .A4(new_n943), .ZN(new_n1029));
  OR2_X1    g604(.A1(new_n942), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1030), .A2(new_n1015), .A3(new_n1026), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(G171), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1006), .B1(new_n1028), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT126), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n498), .A2(new_n853), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n986), .A2(KEYINPUT99), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n490), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n992), .B1(new_n1037), .B2(G1384), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1038), .A2(new_n943), .A3(new_n1022), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n742), .ZN(new_n1040));
  INV_X1    g615(.A(G2084), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1013), .A2(new_n1041), .A3(new_n943), .A4(new_n984), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1000), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT125), .B1(G286), .B2(G8), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(G286), .A2(KEYINPUT125), .A3(G8), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1034), .B1(new_n1043), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1046), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(new_n1044), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n985), .A2(new_n990), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1051), .A2(new_n1041), .B1(new_n1039), .B2(new_n742), .ZN(new_n1052));
  OAI211_X1 g627(.A(KEYINPUT126), .B(new_n1050), .C1(new_n1052), .C2(new_n1000), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1048), .A2(new_n1053), .A3(KEYINPUT51), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1034), .B(new_n1055), .C1(new_n1043), .C2(new_n1047), .ZN(new_n1056));
  AOI21_X1  g631(.A(G1966), .B1(new_n1017), .B2(new_n1022), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1042), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1047), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1054), .A2(new_n1056), .A3(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1015), .A2(new_n1026), .A3(new_n1023), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(G171), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1030), .A2(G301), .A3(new_n1015), .A4(new_n1026), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1033), .A2(new_n1060), .A3(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT56), .B(G2072), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n994), .A2(new_n997), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT119), .ZN(new_n1070));
  INV_X1    g645(.A(G1956), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT119), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n994), .A2(new_n1073), .A3(new_n997), .A4(new_n1068), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1070), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT118), .ZN(new_n1076));
  NAND3_X1  g651(.A1(G299), .A2(new_n1076), .A3(KEYINPUT57), .ZN(new_n1077));
  OR2_X1    g652(.A1(new_n1076), .A2(KEYINPUT57), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1076), .A2(KEYINPUT57), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n563), .A2(new_n567), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1075), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1081), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1070), .A2(new_n1083), .A3(new_n1072), .A4(new_n1074), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1082), .A2(KEYINPUT61), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT124), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT124), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1082), .A2(new_n1087), .A3(KEYINPUT61), .A4(new_n1084), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1008), .A2(new_n753), .A3(new_n1014), .ZN(new_n1090));
  INV_X1    g665(.A(new_n963), .ZN(new_n1091));
  INV_X1    g666(.A(G2067), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1095), .A2(KEYINPUT60), .A3(new_n604), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT60), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n596), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1096), .B(new_n1098), .C1(KEYINPUT60), .C2(new_n1095), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT123), .B(KEYINPUT61), .Z(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1102), .B(G1341), .ZN(new_n1103));
  OAI22_X1  g678(.A1(new_n1025), .A2(G1996), .B1(new_n1091), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n547), .B1(KEYINPUT122), .B2(KEYINPUT59), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(KEYINPUT122), .B2(KEYINPUT59), .ZN(new_n1107));
  NOR2_X1   g682(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1104), .A2(new_n1108), .A3(new_n1105), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1100), .A2(new_n1101), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1089), .A2(new_n1099), .A3(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1082), .B1(new_n1095), .B2(new_n596), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n1084), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1067), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1048), .A2(new_n1053), .A3(KEYINPUT51), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1116));
  OAI21_X1  g691(.A(KEYINPUT62), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1054), .A2(new_n1118), .A3(new_n1056), .A4(new_n1059), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1006), .A2(new_n1062), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1117), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n979), .ZN(new_n1122));
  NOR2_X1   g697(.A1(G305), .A2(G1981), .ZN(new_n1123));
  NOR2_X1   g698(.A1(G288), .A2(G1976), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1123), .B1(new_n969), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT115), .ZN(new_n1126));
  OAI211_X1 g701(.A(G8), .B(new_n963), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1128));
  OAI22_X1  g703(.A1(new_n1122), .A2(new_n999), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT63), .ZN(new_n1130));
  OAI211_X1 g705(.A(G8), .B(G168), .C1(new_n1058), .C2(new_n1057), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1131), .A2(KEYINPUT117), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT117), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1133), .B1(new_n1043), .B2(G168), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1130), .B1(new_n1135), .B2(new_n1006), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n979), .A2(new_n999), .ZN(new_n1137));
  OAI21_X1  g712(.A(G8), .B1(new_n991), .B2(new_n998), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1130), .B1(new_n1138), .B2(new_n981), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1137), .B(new_n1139), .C1(new_n1132), .C2(new_n1134), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1129), .B1(new_n1136), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1121), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n956), .B1(new_n1114), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n950), .A2(new_n947), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1144), .B(KEYINPUT46), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n805), .A2(new_n946), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n945), .A2(new_n1146), .ZN(new_n1147));
  XOR2_X1   g722(.A(KEYINPUT127), .B(KEYINPUT47), .Z(new_n1148));
  AND3_X1   g723(.A1(new_n1145), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1148), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1150));
  NOR3_X1   g725(.A1(new_n944), .A2(G1986), .A3(G290), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT48), .ZN(new_n1152));
  OAI22_X1  g727(.A1(new_n1149), .A2(new_n1150), .B1(new_n954), .B2(new_n1152), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n949), .A2(new_n695), .A3(new_n697), .A4(new_n951), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n785), .A2(new_n1092), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n952), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1143), .A2(new_n1157), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g733(.A1(new_n875), .A2(new_n876), .ZN(new_n1160));
  INV_X1    g734(.A(G319), .ZN(new_n1161));
  NOR4_X1   g735(.A1(G229), .A2(new_n1161), .A3(G401), .A4(G227), .ZN(new_n1162));
  NAND3_X1  g736(.A1(new_n1160), .A2(new_n936), .A3(new_n1162), .ZN(G225));
  INV_X1    g737(.A(G225), .ZN(G308));
endmodule


