//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 1 0 1 0 1 1 1 0 1 0 1 1 1 0 1 0 0 0 1 1 0 0 1 1 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n636, new_n637, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n795, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  INV_X1    g001(.A(G211gat), .ZN(new_n203));
  OR2_X1    g002(.A1(KEYINPUT72), .A2(G218gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(KEYINPUT72), .A2(G218gat), .ZN(new_n205));
  AOI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n202), .B1(new_n206), .B2(KEYINPUT22), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(KEYINPUT73), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n207), .B(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G226gat), .ZN(new_n213));
  INV_X1    g012(.A(G233gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217));
  INV_X1    g016(.A(G169gat), .ZN(new_n218));
  INV_X1    g017(.A(G176gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n220), .B(KEYINPUT26), .ZN(new_n221));
  NAND2_X1  g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT67), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT67), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n224), .A2(G169gat), .A3(G176gat), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(KEYINPUT27), .B(G183gat), .ZN(new_n227));
  INV_X1    g026(.A(G190gat), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT28), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AND3_X1   g028(.A1(new_n227), .A2(KEYINPUT28), .A3(new_n228), .ZN(new_n230));
  OAI221_X1 g029(.A(new_n217), .B1(new_n221), .B2(new_n226), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n232));
  AOI22_X1  g031(.A1(new_n223), .A2(new_n225), .B1(new_n220), .B2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n228), .A2(G183gat), .ZN(new_n234));
  INV_X1    g033(.A(G183gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n235), .A2(G190gat), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT24), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n217), .A2(KEYINPUT24), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n232), .A2(G169gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n219), .A2(KEYINPUT66), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G176gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n239), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n233), .A2(new_n237), .A3(new_n238), .A4(new_n243), .ZN(new_n244));
  XOR2_X1   g043(.A(KEYINPUT65), .B(KEYINPUT25), .Z(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT25), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n248), .B1(new_n239), .B2(new_n219), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n233), .A2(new_n237), .A3(new_n238), .A4(new_n249), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n246), .A2(new_n247), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n247), .B1(new_n246), .B2(new_n250), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n231), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT74), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n246), .A2(new_n250), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT68), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n246), .A2(new_n247), .A3(new_n250), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n259), .A2(KEYINPUT74), .A3(new_n231), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n216), .B1(new_n255), .B2(new_n260), .ZN(new_n261));
  AND2_X1   g060(.A1(new_n256), .A2(new_n231), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n215), .A2(KEYINPUT29), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n212), .B1(new_n261), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n262), .A2(new_n215), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n255), .A2(new_n260), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n211), .B(new_n267), .C1(new_n268), .C2(new_n264), .ZN(new_n269));
  XNOR2_X1  g068(.A(G8gat), .B(G36gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(G64gat), .B(G92gat), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n270), .B(new_n271), .Z(new_n272));
  NAND4_X1  g071(.A1(new_n266), .A2(new_n269), .A3(KEYINPUT30), .A4(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT75), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n276));
  INV_X1    g075(.A(G134gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(G127gat), .ZN(new_n278));
  INV_X1    g077(.A(G127gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(G134gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT1), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(G113gat), .ZN(new_n283));
  INV_X1    g082(.A(G120gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G113gat), .A2(G120gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n276), .B1(new_n282), .B2(new_n287), .ZN(new_n288));
  AND2_X1   g087(.A1(G113gat), .A2(G120gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(G113gat), .A2(G120gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G127gat), .B(G134gat), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n291), .A2(new_n292), .A3(KEYINPUT70), .A4(new_n281), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n288), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT69), .B1(new_n289), .B2(new_n290), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT69), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n285), .A2(new_n296), .A3(new_n286), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n295), .A2(new_n297), .A3(new_n281), .ZN(new_n298));
  INV_X1    g097(.A(new_n292), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n253), .A2(new_n302), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n301), .B(new_n231), .C1(new_n251), .C2(new_n252), .ZN(new_n304));
  INV_X1    g103(.A(G227gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n305), .A2(new_n214), .ZN(new_n306));
  XOR2_X1   g105(.A(new_n306), .B(KEYINPUT64), .Z(new_n307));
  NAND3_X1  g106(.A1(new_n303), .A2(new_n304), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT32), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT33), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  XOR2_X1   g110(.A(G15gat), .B(G43gat), .Z(new_n312));
  XNOR2_X1  g111(.A(G71gat), .B(G99gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n312), .B(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n309), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n314), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n308), .B(KEYINPUT32), .C1(new_n310), .C2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n301), .B1(new_n259), .B2(new_n231), .ZN(new_n319));
  INV_X1    g118(.A(new_n304), .ZN(new_n320));
  OAI22_X1  g119(.A1(new_n319), .A2(new_n320), .B1(new_n305), .B2(new_n214), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n303), .A2(new_n304), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n307), .A2(KEYINPUT34), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n321), .A2(KEYINPUT34), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n318), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT79), .ZN(new_n327));
  INV_X1    g126(.A(G228gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n328), .A2(new_n214), .ZN(new_n329));
  INV_X1    g128(.A(new_n207), .ZN(new_n330));
  AND2_X1   g129(.A1(new_n208), .A2(KEYINPUT78), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n208), .A2(KEYINPUT78), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT29), .B1(new_n207), .B2(new_n331), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT3), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AND2_X1   g137(.A1(G155gat), .A2(G162gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(G155gat), .A2(G162gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G141gat), .B(G148gat), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT2), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n343), .B1(G155gat), .B2(G162gat), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n341), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(G141gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(G148gat), .ZN(new_n347));
  INV_X1    g146(.A(G148gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G141gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G155gat), .B(G162gat), .ZN(new_n351));
  INV_X1    g150(.A(G155gat), .ZN(new_n352));
  INV_X1    g151(.A(G162gat), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT2), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n350), .A2(new_n351), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n345), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n338), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n345), .A2(new_n355), .A3(new_n337), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT29), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n211), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n329), .B1(new_n357), .B2(new_n361), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n210), .B(new_n202), .C1(KEYINPUT22), .C2(new_n206), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n207), .A2(new_n209), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT29), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n356), .B1(new_n365), .B2(KEYINPUT3), .ZN(new_n366));
  INV_X1    g165(.A(new_n329), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n367), .B1(new_n211), .B2(new_n360), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(G22gat), .B1(new_n362), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT3), .B1(new_n334), .B2(new_n335), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n345), .A2(new_n355), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n361), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n373), .A2(new_n367), .B1(new_n366), .B2(new_n368), .ZN(new_n374));
  INV_X1    g173(.A(G22gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT77), .B(KEYINPUT31), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(G50gat), .ZN(new_n378));
  XOR2_X1   g177(.A(G78gat), .B(G106gat), .Z(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  AND4_X1   g179(.A1(new_n327), .A2(new_n370), .A3(new_n376), .A4(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT79), .B1(new_n374), .B2(new_n375), .ZN(new_n382));
  AOI22_X1  g181(.A1(new_n382), .A2(new_n380), .B1(new_n370), .B2(new_n376), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n315), .A2(new_n324), .A3(new_n317), .ZN(new_n385));
  AND3_X1   g184(.A1(new_n326), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n272), .B1(new_n266), .B2(new_n269), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT30), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n266), .A2(new_n269), .A3(new_n272), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n372), .A2(new_n294), .A3(new_n300), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT4), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n356), .A2(KEYINPUT3), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n301), .A2(new_n358), .A3(new_n394), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n372), .A2(new_n294), .A3(new_n300), .A4(KEYINPUT4), .ZN(new_n396));
  NAND2_X1  g195(.A1(G225gat), .A2(G233gat), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n393), .A2(new_n395), .A3(new_n396), .A4(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n397), .ZN(new_n399));
  INV_X1    g198(.A(new_n391), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n372), .B1(new_n300), .B2(new_n294), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n398), .A2(KEYINPUT5), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n358), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n337), .B1(new_n345), .B2(new_n355), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n399), .B1(new_n406), .B2(new_n301), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT5), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n407), .A2(new_n408), .A3(new_n393), .A4(new_n396), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  XOR2_X1   g209(.A(G1gat), .B(G29gat), .Z(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(KEYINPUT0), .ZN(new_n412));
  XNOR2_X1  g211(.A(G57gat), .B(G85gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT6), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n403), .A2(new_n414), .A3(new_n409), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n410), .A2(KEYINPUT6), .A3(new_n415), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT35), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AND4_X1   g220(.A1(new_n275), .A2(new_n386), .A3(new_n390), .A4(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n384), .A2(new_n385), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT71), .B1(new_n318), .B2(new_n325), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n324), .B1(new_n315), .B2(new_n317), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT71), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n424), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT76), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n419), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n416), .A2(KEYINPUT76), .A3(new_n418), .A4(new_n417), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(new_n432), .A3(new_n420), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n273), .A2(new_n274), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n273), .A2(new_n274), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n390), .B(new_n433), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  OAI211_X1 g235(.A(KEYINPUT81), .B(KEYINPUT35), .C1(new_n429), .C2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT71), .ZN(new_n439));
  AOI211_X1 g238(.A(new_n439), .B(new_n324), .C1(new_n315), .C2(new_n317), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n440), .A2(new_n425), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n389), .A2(new_n388), .ZN(new_n442));
  INV_X1    g241(.A(new_n387), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n433), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n441), .A2(new_n444), .A3(new_n275), .A4(new_n424), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT81), .B1(new_n445), .B2(KEYINPUT35), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n423), .B1(new_n438), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n441), .A2(KEYINPUT36), .A3(new_n385), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n326), .A2(new_n385), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT36), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n384), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n275), .A2(new_n390), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT80), .ZN(new_n456));
  OR2_X1    g255(.A1(new_n400), .A2(new_n401), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT39), .B1(new_n457), .B2(new_n399), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n393), .A2(new_n395), .A3(new_n396), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n458), .B1(new_n399), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n399), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n414), .B1(new_n461), .B2(KEYINPUT39), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n456), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT40), .ZN(new_n464));
  OR2_X1    g263(.A1(new_n463), .A2(KEYINPUT40), .ZN(new_n465));
  AND4_X1   g264(.A1(new_n416), .A2(new_n455), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n272), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n266), .A2(new_n269), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n467), .B1(new_n468), .B2(KEYINPUT37), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n469), .B1(KEYINPUT37), .B2(new_n468), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT38), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n389), .A2(new_n419), .A3(new_n420), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n267), .B1(new_n268), .B2(new_n264), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT37), .B1(new_n474), .B2(new_n211), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n261), .A2(new_n265), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n476), .A2(new_n212), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n471), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n473), .B1(new_n478), .B2(new_n469), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n384), .B1(new_n472), .B2(new_n479), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n452), .B(new_n454), .C1(new_n466), .C2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n447), .A2(new_n481), .ZN(new_n482));
  XOR2_X1   g281(.A(KEYINPUT85), .B(G29gat), .Z(new_n483));
  INV_X1    g282(.A(G36gat), .ZN(new_n484));
  OR3_X1    g283(.A1(new_n483), .A2(KEYINPUT86), .A3(new_n484), .ZN(new_n485));
  XOR2_X1   g284(.A(G43gat), .B(G50gat), .Z(new_n486));
  INV_X1    g285(.A(KEYINPUT15), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT87), .ZN(new_n489));
  OR3_X1    g288(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT86), .B1(new_n483), .B2(new_n484), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n485), .A2(new_n488), .A3(new_n492), .A4(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n486), .A2(new_n487), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n496), .B(KEYINPUT17), .ZN(new_n497));
  XNOR2_X1  g296(.A(G15gat), .B(G22gat), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT16), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n498), .B1(new_n499), .B2(G1gat), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT88), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n500), .B(new_n501), .C1(G1gat), .C2(new_n498), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n502), .B(G8gat), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n497), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(G229gat), .A2(G233gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n496), .A2(new_n503), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT18), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n505), .A2(KEYINPUT18), .A3(new_n506), .A4(new_n507), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT89), .B1(new_n496), .B2(new_n503), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(new_n507), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n506), .B(KEYINPUT13), .Z(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n510), .A2(new_n511), .A3(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G169gat), .B(G197gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n517), .B(KEYINPUT83), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(G113gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(new_n346), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n519), .B(new_n521), .ZN(new_n522));
  XOR2_X1   g321(.A(KEYINPUT84), .B(KEYINPUT12), .Z(new_n523));
  XOR2_X1   g322(.A(new_n522), .B(new_n523), .Z(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n516), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n510), .A2(new_n524), .A3(new_n511), .A4(new_n515), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n528), .A2(KEYINPUT90), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT90), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n530), .B1(new_n526), .B2(new_n527), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G232gat), .A2(G233gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT41), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(new_n536), .B(KEYINPUT96), .Z(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(G134gat), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n534), .A2(new_n535), .ZN(new_n540));
  NAND2_X1  g339(.A1(G99gat), .A2(G106gat), .ZN(new_n541));
  INV_X1    g340(.A(G85gat), .ZN(new_n542));
  INV_X1    g341(.A(G92gat), .ZN(new_n543));
  AOI22_X1  g342(.A1(KEYINPUT8), .A2(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(KEYINPUT97), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n545));
  NAND3_X1  g344(.A1(KEYINPUT97), .A2(G85gat), .A3(G92gat), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT7), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n544), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(G99gat), .B(G106gat), .Z(new_n550));
  XOR2_X1   g349(.A(new_n549), .B(new_n550), .Z(new_n551));
  AOI21_X1  g350(.A(new_n540), .B1(new_n496), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT99), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n551), .B(KEYINPUT98), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n497), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT100), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n553), .A2(KEYINPUT100), .A3(new_n555), .ZN(new_n559));
  XNOR2_X1  g358(.A(G190gat), .B(G218gat), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n560), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n556), .A2(new_n557), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n561), .A2(new_n353), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n353), .B1(new_n561), .B2(new_n563), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n539), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n566), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n568), .A2(new_n538), .A3(new_n564), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(G71gat), .A2(G78gat), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n571), .B(KEYINPUT91), .Z(new_n572));
  XOR2_X1   g371(.A(G57gat), .B(G64gat), .Z(new_n573));
  NAND2_X1  g372(.A1(G71gat), .A2(G78gat), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT9), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n572), .A2(new_n577), .A3(new_n574), .ZN(new_n578));
  INV_X1    g377(.A(new_n571), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(new_n574), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT92), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT92), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n579), .A2(new_n582), .A3(new_n574), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n581), .A2(new_n576), .A3(new_n573), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n578), .A2(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(KEYINPUT93), .B(KEYINPUT21), .Z(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT94), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT95), .ZN(new_n589));
  XNOR2_X1  g388(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XOR2_X1   g390(.A(G183gat), .B(G211gat), .Z(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT21), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n504), .B1(new_n594), .B2(new_n585), .ZN(new_n595));
  XNOR2_X1  g394(.A(G127gat), .B(G155gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(G231gat), .A2(G233gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n595), .B(new_n598), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n593), .A2(new_n599), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n570), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(G230gat), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n605), .A2(new_n214), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n551), .B(new_n585), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT10), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n551), .A2(KEYINPUT10), .A3(new_n578), .A4(new_n584), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n606), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NOR3_X1   g410(.A1(new_n607), .A2(new_n605), .A3(new_n214), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G120gat), .B(G148gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(G176gat), .B(G204gat), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n614), .B(new_n615), .Z(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n613), .A2(new_n617), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n482), .A2(new_n533), .A3(new_n604), .A4(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n622), .A2(new_n433), .ZN(new_n623));
  XNOR2_X1  g422(.A(KEYINPUT101), .B(G1gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(G1324gat));
  INV_X1    g424(.A(new_n455), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(KEYINPUT16), .B(G8gat), .Z(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(G8gat), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n629), .B1(new_n630), .B2(new_n627), .ZN(new_n631));
  MUX2_X1   g430(.A(new_n629), .B(new_n631), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g431(.A(G15gat), .B1(new_n622), .B2(new_n452), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n449), .A2(G15gat), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n633), .B1(new_n622), .B2(new_n634), .ZN(G1326gat));
  NOR2_X1   g434(.A1(new_n622), .A2(new_n384), .ZN(new_n636));
  XOR2_X1   g435(.A(KEYINPUT43), .B(G22gat), .Z(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(G1327gat));
  NAND2_X1  g437(.A1(new_n603), .A2(new_n621), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n567), .A2(new_n569), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n482), .A2(new_n641), .A3(new_n533), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n433), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n643), .A2(new_n644), .A3(new_n483), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT45), .ZN(new_n646));
  OAI21_X1  g445(.A(KEYINPUT35), .B1(new_n429), .B2(new_n436), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT81), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n437), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT102), .B1(new_n650), .B2(new_n423), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT102), .ZN(new_n652));
  AOI211_X1 g451(.A(new_n652), .B(new_n422), .C1(new_n649), .C2(new_n437), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n481), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n640), .A2(KEYINPUT44), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT44), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n657), .B1(new_n482), .B2(new_n570), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n528), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n639), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(new_n433), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n646), .B1(new_n664), .B2(new_n483), .ZN(G1328gat));
  NOR3_X1   g464(.A1(new_n642), .A2(G36gat), .A3(new_n626), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT103), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT46), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(G36gat), .B1(new_n663), .B2(new_n626), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n668), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n671), .A2(KEYINPUT104), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n673), .B1(new_n667), .B2(new_n668), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n669), .B(new_n670), .C1(new_n672), .C2(new_n674), .ZN(G1329gat));
  INV_X1    g474(.A(G43gat), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n452), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n655), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n447), .A2(new_n652), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n650), .A2(KEYINPUT102), .A3(new_n423), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n678), .B1(new_n681), .B2(new_n481), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n662), .B(new_n677), .C1(new_n682), .C2(new_n658), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n676), .B1(new_n642), .B2(new_n449), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(KEYINPUT106), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n683), .A2(new_n684), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT47), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT106), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n683), .A2(new_n690), .A3(new_n684), .A4(new_n685), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n687), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(KEYINPUT107), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT107), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n687), .A2(new_n689), .A3(new_n694), .A4(new_n691), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(G1330gat));
  NOR3_X1   g495(.A1(new_n642), .A2(G50gat), .A3(new_n384), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n660), .A2(new_n453), .A3(new_n662), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n697), .B1(new_n698), .B2(G50gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g499(.A(new_n621), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n604), .A2(new_n661), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n702), .B1(new_n681), .B2(new_n481), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(new_n644), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g504(.A(new_n626), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT108), .Z(new_n708));
  NOR2_X1   g507(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1333gat));
  INV_X1    g509(.A(new_n452), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n703), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n449), .A2(G71gat), .ZN(new_n713));
  AOI22_X1  g512(.A1(new_n712), .A2(G71gat), .B1(new_n703), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g514(.A1(new_n703), .A2(new_n453), .ZN(new_n716));
  XOR2_X1   g515(.A(KEYINPUT109), .B(G78gat), .Z(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(G1335gat));
  NAND2_X1  g517(.A1(new_n603), .A2(new_n661), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n719), .A2(new_n621), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n721), .B1(new_n656), .B2(new_n659), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n722), .A2(new_n644), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n719), .A2(new_n640), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n654), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT51), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n654), .A2(KEYINPUT51), .A3(new_n724), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n701), .A2(new_n542), .A3(new_n644), .ZN(new_n731));
  OAI22_X1  g530(.A1(new_n723), .A2(new_n542), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT110), .ZN(G1336gat));
  NAND3_X1  g532(.A1(new_n455), .A2(new_n543), .A3(new_n701), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n734), .B(KEYINPUT111), .Z(new_n735));
  NAND3_X1  g534(.A1(new_n725), .A2(KEYINPUT112), .A3(new_n726), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n735), .B(new_n736), .C1(new_n729), .C2(KEYINPUT112), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n455), .B(new_n720), .C1(new_n682), .C2(new_n658), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(G92gat), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT52), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT113), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n660), .A2(KEYINPUT113), .A3(new_n455), .A4(new_n720), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n743), .A2(G92gat), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT52), .B1(new_n729), .B2(new_n735), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n745), .A2(KEYINPUT114), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT114), .B1(new_n745), .B2(new_n746), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n741), .B1(new_n747), .B2(new_n748), .ZN(G1337gat));
  AND2_X1   g548(.A1(new_n722), .A2(new_n711), .ZN(new_n750));
  INV_X1    g549(.A(G99gat), .ZN(new_n751));
  OR3_X1    g550(.A1(new_n621), .A2(new_n449), .A3(G99gat), .ZN(new_n752));
  OAI22_X1  g551(.A1(new_n750), .A2(new_n751), .B1(new_n730), .B2(new_n752), .ZN(G1338gat));
  NAND2_X1  g552(.A1(new_n722), .A2(new_n453), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G106gat), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT53), .ZN(new_n756));
  OR3_X1    g555(.A1(new_n621), .A2(G106gat), .A3(new_n384), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n755), .B(new_n756), .C1(new_n730), .C2(new_n757), .ZN(new_n758));
  XOR2_X1   g557(.A(new_n757), .B(KEYINPUT115), .Z(new_n759));
  OAI211_X1 g558(.A(new_n736), .B(new_n759), .C1(new_n729), .C2(KEYINPUT112), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n760), .A2(new_n755), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n758), .B1(new_n761), .B2(new_n756), .ZN(G1339gat));
  INV_X1    g561(.A(KEYINPUT54), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n611), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n609), .A2(new_n610), .A3(new_n606), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n616), .B1(new_n611), .B2(new_n763), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n618), .B1(new_n769), .B2(KEYINPUT55), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(KEYINPUT55), .B2(new_n769), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n513), .A2(new_n514), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n506), .B1(new_n505), .B2(new_n507), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n522), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n527), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n776), .A2(new_n567), .A3(new_n569), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n528), .B(new_n770), .C1(KEYINPUT55), .C2(new_n769), .ZN(new_n778));
  OR2_X1    g577(.A1(new_n775), .A2(new_n621), .ZN(new_n779));
  AOI22_X1  g578(.A1(new_n567), .A2(new_n569), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n603), .B1(new_n777), .B2(new_n780), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n640), .A2(new_n661), .A3(new_n602), .A4(new_n621), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n783), .A2(new_n644), .A3(new_n626), .A4(new_n386), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n784), .A2(new_n283), .A3(new_n532), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n433), .B1(new_n781), .B2(new_n782), .ZN(new_n786));
  INV_X1    g585(.A(new_n429), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n455), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n528), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n785), .B1(new_n790), .B2(new_n283), .ZN(G1340gat));
  NOR3_X1   g590(.A1(new_n784), .A2(new_n284), .A3(new_n621), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n701), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n792), .B1(new_n793), .B2(new_n284), .ZN(G1341gat));
  NAND3_X1  g593(.A1(new_n789), .A2(new_n279), .A3(new_n602), .ZN(new_n795));
  OAI21_X1  g594(.A(G127gat), .B1(new_n784), .B2(new_n603), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(G1342gat));
  NAND2_X1  g596(.A1(new_n570), .A2(new_n626), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(KEYINPUT116), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n788), .A2(G134gat), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n801), .A2(KEYINPUT56), .ZN(new_n802));
  OAI21_X1  g601(.A(G134gat), .B1(new_n784), .B2(new_n640), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n801), .A2(KEYINPUT56), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(G1343gat));
  NAND2_X1  g604(.A1(new_n626), .A2(new_n644), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n711), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n384), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  XNOR2_X1  g609(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n768), .A2(KEYINPUT118), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT118), .B1(new_n768), .B2(new_n811), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n770), .B(KEYINPUT119), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n529), .B2(new_n531), .ZN(new_n815));
  OR2_X1    g614(.A1(new_n812), .A2(new_n813), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT119), .B1(new_n816), .B2(new_n770), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n779), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n640), .ZN(new_n819));
  INV_X1    g618(.A(new_n777), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n603), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n810), .B1(new_n822), .B2(new_n782), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT57), .B1(new_n783), .B2(new_n453), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n807), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n528), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n452), .A2(new_n453), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(KEYINPUT120), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n786), .A2(new_n829), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n830), .A2(new_n626), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n532), .A2(G141gat), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(KEYINPUT121), .ZN(new_n833));
  AOI22_X1  g632(.A1(new_n827), .A2(G141gat), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT58), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n346), .B1(new_n826), .B2(new_n533), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n831), .A2(new_n833), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n835), .ZN(new_n838));
  OAI22_X1  g637(.A1(new_n834), .A2(new_n835), .B1(new_n836), .B2(new_n838), .ZN(G1344gat));
  NAND3_X1  g638(.A1(new_n831), .A2(new_n348), .A3(new_n701), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT59), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n604), .A2(KEYINPUT122), .A3(new_n532), .A4(new_n621), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT122), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n640), .A2(new_n602), .A3(new_n621), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n843), .B1(new_n844), .B2(new_n533), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n777), .B1(new_n818), .B2(new_n640), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n842), .B(new_n845), .C1(new_n602), .C2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n453), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n808), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n783), .A2(new_n809), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(new_n701), .A3(new_n807), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n841), .B1(new_n852), .B2(G148gat), .ZN(new_n853));
  AOI211_X1 g652(.A(KEYINPUT59), .B(new_n348), .C1(new_n826), .C2(new_n701), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n840), .B1(new_n853), .B2(new_n854), .ZN(G1345gat));
  OAI21_X1  g654(.A(G155gat), .B1(new_n825), .B2(new_n603), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n831), .A2(new_n352), .A3(new_n602), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(G1346gat));
  OAI21_X1  g657(.A(G162gat), .B1(new_n825), .B2(new_n640), .ZN(new_n859));
  INV_X1    g658(.A(new_n799), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n830), .A2(new_n353), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(G1347gat));
  AOI21_X1  g661(.A(new_n644), .B1(new_n781), .B2(new_n782), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n863), .A2(new_n787), .A3(new_n455), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n864), .A2(G169gat), .A3(new_n661), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n865), .B(KEYINPUT123), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n626), .A2(new_n644), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n783), .A2(new_n386), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(KEYINPUT124), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT124), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n783), .A2(new_n870), .A3(new_n386), .A4(new_n867), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n218), .B1(new_n872), .B2(new_n533), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n866), .A2(new_n873), .ZN(G1348gat));
  AOI21_X1  g673(.A(new_n621), .B1(new_n240), .B2(new_n242), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n864), .A2(new_n621), .ZN(new_n876));
  AOI22_X1  g675(.A1(new_n872), .A2(new_n875), .B1(new_n876), .B2(new_n219), .ZN(G1349gat));
  NAND2_X1  g676(.A1(new_n602), .A2(new_n227), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n864), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n869), .A2(new_n602), .A3(new_n871), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n879), .B1(new_n880), .B2(G183gat), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n881), .B(KEYINPUT60), .Z(G1350gat));
  OR3_X1    g681(.A1(new_n864), .A2(G190gat), .A3(new_n640), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n869), .A2(new_n570), .A3(new_n871), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT125), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n885), .A3(G190gat), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n885), .B1(new_n884), .B2(G190gat), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n887), .A2(new_n888), .A3(KEYINPUT61), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n884), .A2(G190gat), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT125), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n890), .B1(new_n892), .B2(new_n886), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n883), .B1(new_n889), .B2(new_n893), .ZN(G1351gat));
  NAND2_X1  g693(.A1(new_n867), .A2(new_n452), .ZN(new_n895));
  INV_X1    g694(.A(G197gat), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n895), .A2(new_n532), .A3(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT126), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n898), .B1(new_n849), .B2(new_n850), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT57), .B1(new_n847), .B2(new_n453), .ZN(new_n900));
  INV_X1    g699(.A(new_n850), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n900), .A2(KEYINPUT126), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n897), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  AND4_X1   g702(.A1(new_n453), .A2(new_n863), .A3(new_n455), .A4(new_n452), .ZN(new_n904));
  AOI21_X1  g703(.A(G197gat), .B1(new_n904), .B2(new_n528), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n903), .A2(KEYINPUT127), .A3(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT127), .ZN(new_n908));
  INV_X1    g707(.A(new_n897), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n849), .A2(new_n898), .A3(new_n850), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT126), .B1(new_n900), .B2(new_n901), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n908), .B1(new_n912), .B2(new_n905), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n907), .A2(new_n913), .ZN(G1352gat));
  INV_X1    g713(.A(G204gat), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n904), .A2(new_n915), .A3(new_n701), .ZN(new_n916));
  XOR2_X1   g715(.A(new_n916), .B(KEYINPUT62), .Z(new_n917));
  AOI211_X1 g716(.A(new_n621), .B(new_n895), .C1(new_n910), .C2(new_n911), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n918), .B2(new_n915), .ZN(G1353gat));
  NAND3_X1  g718(.A1(new_n904), .A2(new_n203), .A3(new_n602), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n895), .A2(new_n603), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n851), .A2(new_n921), .ZN(new_n922));
  AND3_X1   g721(.A1(new_n922), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT63), .B1(new_n922), .B2(G211gat), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n920), .B1(new_n923), .B2(new_n924), .ZN(G1354gat));
  AOI21_X1  g724(.A(G218gat), .B1(new_n904), .B2(new_n570), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n895), .B1(new_n910), .B2(new_n911), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n640), .B1(new_n204), .B2(new_n205), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(G1355gat));
endmodule


